
module eth_clockgen_test_1 ( Clk, Reset, Divider, MdcEn, MdcEn_n, Mdc, 
        eth_top_test_point_11887_in, test_si, test_se );
  input [7:0] Divider;
  input Clk, Reset, eth_top_test_point_11887_in, test_si, test_se;
  output MdcEn, MdcEn_n, Mdc;
  wire   N15, N16, N17, N18, N19, N20, N21, n13, n23, n1, n56, n57, n58, n59,
         n60, n61, n43, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42;
  wire   [7:1] TempDivider;
  assign TempDivider[7] = Divider[7];
  assign TempDivider[6] = Divider[6];
  assign TempDivider[5] = Divider[5];
  assign TempDivider[4] = Divider[4];
  assign TempDivider[3] = Divider[3];
  assign TempDivider[2] = Divider[2];

  SDFFASX1 \Counter_reg[0]  ( .D(N15), .SI(test_si), .SE(test_se), .CLK(Clk), 
        .SETB(n42), .Q(n61), .QN(n41) );
  SDFFARX1 \Counter_reg[1]  ( .D(N16), .SI(n61), .SE(test_se), .CLK(Clk), 
        .RSTB(n42), .Q(n60), .QN(n40) );
  SDFFARX1 \Counter_reg[2]  ( .D(N17), .SI(n60), .SE(test_se), .CLK(Clk), 
        .RSTB(n42), .Q(n59), .QN(n39) );
  SDFFARX1 \Counter_reg[3]  ( .D(N18), .SI(n59), .SE(test_se), .CLK(Clk), 
        .RSTB(n42), .Q(n58), .QN(n38) );
  SDFFARX1 \Counter_reg[4]  ( .D(N19), .SI(n58), .SE(test_se), .CLK(Clk), 
        .RSTB(n42), .Q(n57) );
  SDFFARX1 \Counter_reg[5]  ( .D(N20), .SI(n57), .SE(test_se), .CLK(Clk), 
        .RSTB(n42), .Q(n56), .QN(n37) );
  SDFFARX1 \Counter_reg[6]  ( .D(N21), .SI(n56), .SE(test_se), .CLK(Clk), 
        .RSTB(n42), .Q(n1), .QN(n43) );
  SDFFARX1 Mdc_reg ( .D(n13), .SI(n1), .SE(test_se), .CLK(Clk), .RSTB(n42), 
        .Q(Mdc), .QN(n23) );
  INVX0 U3 ( .INP(eth_top_test_point_11887_in), .ZN(n42) );
  AO21X1 U4 ( .IN1(n2), .IN2(Mdc), .IN3(MdcEn), .Q(n13) );
  NAND2X0 U5 ( .IN1(n3), .IN2(n4), .QN(N21) );
  OR3X1 U6 ( .IN1(n2), .IN2(n5), .IN3(n6), .Q(n4) );
  INVX0 U7 ( .INP(TempDivider[7]), .ZN(n6) );
  AO21X1 U8 ( .IN1(n37), .IN2(n7), .IN3(n43), .Q(n3) );
  MUX21X1 U9 ( .IN1(n8), .IN2(n9), .S(n2), .Q(N20) );
  XNOR2X1 U10 ( .IN1(n37), .IN2(n7), .Q(n9) );
  AO21X1 U11 ( .IN1(TempDivider[6]), .IN2(n10), .IN3(n5), .Q(n8) );
  NOR2X0 U12 ( .IN1(n10), .IN2(TempDivider[6]), .QN(n5) );
  INVX0 U13 ( .INP(n11), .ZN(n10) );
  MUX21X1 U14 ( .IN1(n12), .IN2(n14), .S(n2), .Q(N19) );
  AO21X1 U15 ( .IN1(n15), .IN2(n57), .IN3(n7), .Q(n14) );
  AO21X1 U16 ( .IN1(TempDivider[5]), .IN2(n16), .IN3(n11), .Q(n12) );
  NOR2X0 U17 ( .IN1(n16), .IN2(TempDivider[5]), .QN(n11) );
  INVX0 U18 ( .INP(n17), .ZN(n16) );
  MUX21X1 U19 ( .IN1(n18), .IN2(n19), .S(n2), .Q(N18) );
  OAI21X1 U20 ( .IN1(n20), .IN2(n38), .IN3(n15), .QN(n19) );
  AO21X1 U21 ( .IN1(TempDivider[4]), .IN2(n21), .IN3(n17), .Q(n18) );
  NOR2X0 U22 ( .IN1(n21), .IN2(TempDivider[4]), .QN(n17) );
  INVX0 U23 ( .INP(n22), .ZN(n21) );
  MUX21X1 U24 ( .IN1(n24), .IN2(n25), .S(n2), .Q(N17) );
  OAI21X1 U25 ( .IN1(n26), .IN2(n39), .IN3(n27), .QN(n25) );
  AO21X1 U26 ( .IN1(TempDivider[3]), .IN2(n28), .IN3(n22), .Q(n24) );
  NOR2X0 U27 ( .IN1(n28), .IN2(TempDivider[3]), .QN(n22) );
  INVX0 U28 ( .INP(n29), .ZN(n28) );
  MUX21X1 U29 ( .IN1(n30), .IN2(n31), .S(n2), .Q(N16) );
  OAI21X1 U30 ( .IN1(n41), .IN2(n40), .IN3(n32), .QN(n31) );
  AO21X1 U31 ( .IN1(TempDivider[2]), .IN2(n33), .IN3(n29), .Q(n30) );
  NOR2X0 U32 ( .IN1(n33), .IN2(TempDivider[2]), .QN(n29) );
  INVX0 U33 ( .INP(n34), .ZN(n33) );
  MUX21X1 U34 ( .IN1(n34), .IN2(n41), .S(n2), .Q(N15) );
  NOR2X0 U35 ( .IN1(Divider[1]), .IN2(n35), .QN(n34) );
  NOR4X0 U36 ( .IN1(n36), .IN2(TempDivider[2]), .IN3(TempDivider[4]), .IN4(
        TempDivider[3]), .QN(n35) );
  OR3X1 U37 ( .IN1(TempDivider[6]), .IN2(TempDivider[7]), .IN3(TempDivider[5]), 
        .Q(n36) );
  NOR2X0 U38 ( .IN1(n23), .IN2(n2), .QN(MdcEn_n) );
  NOR2X0 U39 ( .IN1(Mdc), .IN2(n2), .QN(MdcEn) );
  NAND3X0 U40 ( .IN1(n43), .IN2(n7), .IN3(n37), .QN(n2) );
  NOR2X0 U41 ( .IN1(n57), .IN2(n15), .QN(n7) );
  NAND2X0 U42 ( .IN1(n38), .IN2(n20), .QN(n15) );
  INVX0 U43 ( .INP(n27), .ZN(n20) );
  NAND2X0 U44 ( .IN1(n39), .IN2(n26), .QN(n27) );
  INVX0 U45 ( .INP(n32), .ZN(n26) );
  NAND2X0 U46 ( .IN1(n40), .IN2(n41), .QN(n32) );
endmodule


module eth_shiftreg_test_1 ( Clk, Reset, MdcEn_n, Mdi, Fiad, Rgad, CtrlData, 
        WriteOp, ByteSelect, LatchByte, ShiftedBit, Prsd, LinkFail, 
        eth_top_test_point_11887_in, test_si, test_se );
  input [4:0] Fiad;
  input [4:0] Rgad;
  input [15:0] CtrlData;
  input [3:0] ByteSelect;
  input [1:0] LatchByte;
  output [15:0] Prsd;
  input Clk, Reset, MdcEn_n, Mdi, WriteOp, eth_top_test_point_11887_in,
         test_si, test_se;
  output ShiftedBit, LinkFail;
  wire   n62, n64, n66, n68, n70, n72, n74, n77, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n40, n41, n42,
         n43, n75, n78, n96, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n44;

  SDFFARX1 \ShiftReg_reg[0]  ( .D(n77), .SI(Prsd[15]), .SE(test_se), .CLK(Clk), 
        .RSTB(n44), .Q(n96) );
  SDFFARX1 \ShiftReg_reg[1]  ( .D(n74), .SI(n96), .SE(test_se), .CLK(Clk), 
        .RSTB(n44), .Q(n75), .QN(n39) );
  SDFFARX1 \ShiftReg_reg[2]  ( .D(n72), .SI(n75), .SE(test_se), .CLK(Clk), 
        .RSTB(n44), .Q(n43) );
  SDFFARX1 \ShiftReg_reg[3]  ( .D(n70), .SI(n43), .SE(test_se), .CLK(Clk), 
        .RSTB(n44), .Q(n42) );
  SDFFARX1 \ShiftReg_reg[4]  ( .D(n68), .SI(n42), .SE(test_se), .CLK(Clk), 
        .RSTB(n44), .Q(n41) );
  SDFFARX1 \ShiftReg_reg[5]  ( .D(n66), .SI(n41), .SE(test_se), .CLK(Clk), 
        .RSTB(n44), .Q(n78) );
  SDFFARX1 \ShiftReg_reg[6]  ( .D(n64), .SI(n78), .SE(test_se), .CLK(Clk), 
        .RSTB(n44), .Q(n40) );
  SDFFARX1 \ShiftReg_reg[7]  ( .D(n62), .SI(n40), .SE(test_se), .CLK(Clk), 
        .RSTB(n44), .Q(ShiftedBit) );
  SDFFARX1 \Prsd_reg[15]  ( .D(n95), .SI(Prsd[14]), .SE(test_se), .CLK(Clk), 
        .RSTB(n44), .Q(Prsd[15]) );
  SDFFARX1 \Prsd_reg[14]  ( .D(n94), .SI(Prsd[13]), .SE(test_se), .CLK(Clk), 
        .RSTB(n44), .Q(Prsd[14]) );
  SDFFARX1 \Prsd_reg[13]  ( .D(n93), .SI(Prsd[12]), .SE(test_se), .CLK(Clk), 
        .RSTB(n44), .Q(Prsd[13]) );
  SDFFARX1 \Prsd_reg[12]  ( .D(n92), .SI(Prsd[11]), .SE(test_se), .CLK(Clk), 
        .RSTB(n44), .Q(Prsd[12]) );
  SDFFARX1 \Prsd_reg[11]  ( .D(n91), .SI(Prsd[10]), .SE(test_se), .CLK(Clk), 
        .RSTB(n44), .Q(Prsd[11]) );
  SDFFARX1 \Prsd_reg[10]  ( .D(n90), .SI(Prsd[9]), .SE(test_se), .CLK(Clk), 
        .RSTB(n44), .Q(Prsd[10]) );
  SDFFARX1 \Prsd_reg[9]  ( .D(n89), .SI(Prsd[8]), .SE(test_se), .CLK(Clk), 
        .RSTB(n44), .Q(Prsd[9]) );
  SDFFARX1 \Prsd_reg[8]  ( .D(n88), .SI(Prsd[7]), .SE(test_se), .CLK(Clk), 
        .RSTB(n44), .Q(Prsd[8]) );
  SDFFARX1 \Prsd_reg[7]  ( .D(n87), .SI(Prsd[6]), .SE(test_se), .CLK(Clk), 
        .RSTB(n44), .Q(Prsd[7]) );
  SDFFARX1 \Prsd_reg[6]  ( .D(n86), .SI(Prsd[5]), .SE(test_se), .CLK(Clk), 
        .RSTB(n44), .Q(Prsd[6]) );
  SDFFARX1 \Prsd_reg[5]  ( .D(n85), .SI(Prsd[4]), .SE(test_se), .CLK(Clk), 
        .RSTB(n44), .Q(Prsd[5]) );
  SDFFARX1 \Prsd_reg[4]  ( .D(n84), .SI(Prsd[3]), .SE(test_se), .CLK(Clk), 
        .RSTB(n44), .Q(Prsd[4]) );
  SDFFARX1 \Prsd_reg[3]  ( .D(n83), .SI(Prsd[2]), .SE(test_se), .CLK(Clk), 
        .RSTB(n44), .Q(Prsd[3]) );
  SDFFARX1 \Prsd_reg[2]  ( .D(n82), .SI(Prsd[1]), .SE(test_se), .CLK(Clk), 
        .RSTB(n44), .Q(Prsd[2]) );
  SDFFARX1 \Prsd_reg[1]  ( .D(n81), .SI(Prsd[0]), .SE(test_se), .CLK(Clk), 
        .RSTB(n44), .Q(Prsd[1]) );
  SDFFARX1 \Prsd_reg[0]  ( .D(n80), .SI(LinkFail), .SE(test_se), .CLK(Clk), 
        .RSTB(n44), .Q(Prsd[0]) );
  SDFFARX1 LinkFail_reg ( .D(n79), .SI(test_si), .SE(test_se), .CLK(Clk), 
        .RSTB(n44), .Q(LinkFail) );
  INVX0 U3 ( .INP(eth_top_test_point_11887_in), .ZN(n44) );
  MUX21X1 U4 ( .IN1(Prsd[15]), .IN2(n40), .S(n1), .Q(n95) );
  MUX21X1 U5 ( .IN1(Prsd[14]), .IN2(n78), .S(n1), .Q(n94) );
  MUX21X1 U6 ( .IN1(Prsd[13]), .IN2(n41), .S(n1), .Q(n93) );
  MUX21X1 U7 ( .IN1(Prsd[12]), .IN2(n42), .S(n1), .Q(n92) );
  MUX21X1 U8 ( .IN1(Prsd[11]), .IN2(n43), .S(n1), .Q(n91) );
  MUX21X1 U9 ( .IN1(Prsd[10]), .IN2(n75), .S(n1), .Q(n90) );
  MUX21X1 U10 ( .IN1(Prsd[9]), .IN2(n96), .S(n1), .Q(n89) );
  MUX21X1 U11 ( .IN1(Prsd[8]), .IN2(Mdi), .S(n1), .Q(n88) );
  AND3X1 U12 ( .IN1(n2), .IN2(n3), .IN3(LatchByte[1]), .Q(n1) );
  INVX0 U13 ( .INP(LatchByte[0]), .ZN(n3) );
  MUX21X1 U14 ( .IN1(Prsd[7]), .IN2(n40), .S(n4), .Q(n87) );
  MUX21X1 U15 ( .IN1(Prsd[6]), .IN2(n78), .S(n4), .Q(n86) );
  MUX21X1 U16 ( .IN1(Prsd[5]), .IN2(n41), .S(n4), .Q(n85) );
  MUX21X1 U17 ( .IN1(Prsd[4]), .IN2(n42), .S(n4), .Q(n84) );
  MUX21X1 U18 ( .IN1(Prsd[3]), .IN2(n43), .S(n4), .Q(n83) );
  MUX21X1 U19 ( .IN1(Prsd[2]), .IN2(n75), .S(n4), .Q(n82) );
  MUX21X1 U20 ( .IN1(Prsd[1]), .IN2(n96), .S(n4), .Q(n81) );
  MUX21X1 U21 ( .IN1(Prsd[0]), .IN2(Mdi), .S(n4), .Q(n80) );
  MUX21X1 U22 ( .IN1(LinkFail), .IN2(n39), .S(n5), .Q(n79) );
  NOR4X0 U23 ( .IN1(n6), .IN2(Rgad[2]), .IN3(Rgad[4]), .IN4(Rgad[3]), .QN(n5)
         );
  NAND3X0 U24 ( .IN1(n4), .IN2(n7), .IN3(Rgad[0]), .QN(n6) );
  INVX0 U25 ( .INP(Rgad[1]), .ZN(n7) );
  AND2X1 U26 ( .IN1(LatchByte[0]), .IN2(n2), .Q(n4) );
  AO21X1 U27 ( .IN1(Mdi), .IN2(n2), .IN3(n8), .Q(n77) );
  MUX21X1 U28 ( .IN1(n96), .IN2(n9), .S(MdcEn_n), .Q(n8) );
  AO222X1 U29 ( .IN1(CtrlData[8]), .IN2(ByteSelect[2]), .IN3(Fiad[1]), .IN4(
        ByteSelect[0]), .IN5(CtrlData[0]), .IN6(ByteSelect[3]), .Q(n9) );
  MUX21X1 U30 ( .IN1(n75), .IN2(n10), .S(MdcEn_n), .Q(n74) );
  OR4X1 U31 ( .IN1(n11), .IN2(n12), .IN3(ByteSelect[1]), .IN4(n13), .Q(n10) );
  AND2X1 U32 ( .IN1(CtrlData[9]), .IN2(ByteSelect[2]), .Q(n13) );
  MUX21X1 U33 ( .IN1(n14), .IN2(Fiad[2]), .S(ByteSelect[0]), .Q(n12) );
  AND2X1 U34 ( .IN1(n15), .IN2(n96), .Q(n14) );
  AND2X1 U35 ( .IN1(CtrlData[1]), .IN2(ByteSelect[3]), .Q(n11) );
  AO21X1 U36 ( .IN1(n2), .IN2(n75), .IN3(n16), .Q(n72) );
  MUX21X1 U37 ( .IN1(n43), .IN2(n17), .S(MdcEn_n), .Q(n16) );
  AO221X1 U38 ( .IN1(CtrlData[10]), .IN2(ByteSelect[2]), .IN3(CtrlData[2]), 
        .IN4(ByteSelect[3]), .IN5(n18), .Q(n17) );
  AO22X1 U39 ( .IN1(ByteSelect[1]), .IN2(Rgad[0]), .IN3(Fiad[3]), .IN4(
        ByteSelect[0]), .Q(n18) );
  AO21X1 U40 ( .IN1(n2), .IN2(n43), .IN3(n19), .Q(n70) );
  MUX21X1 U41 ( .IN1(n42), .IN2(n20), .S(MdcEn_n), .Q(n19) );
  AO221X1 U42 ( .IN1(CtrlData[11]), .IN2(ByteSelect[2]), .IN3(CtrlData[3]), 
        .IN4(ByteSelect[3]), .IN5(n21), .Q(n20) );
  AO22X1 U43 ( .IN1(Rgad[1]), .IN2(ByteSelect[1]), .IN3(Fiad[4]), .IN4(
        ByteSelect[0]), .Q(n21) );
  AO21X1 U44 ( .IN1(n2), .IN2(n42), .IN3(n22), .Q(n68) );
  MUX21X1 U45 ( .IN1(n41), .IN2(n23), .S(MdcEn_n), .Q(n22) );
  AO221X1 U46 ( .IN1(CtrlData[12]), .IN2(ByteSelect[2]), .IN3(CtrlData[4]), 
        .IN4(ByteSelect[3]), .IN5(n24), .Q(n23) );
  AO22X1 U47 ( .IN1(Rgad[2]), .IN2(ByteSelect[1]), .IN3(WriteOp), .IN4(
        ByteSelect[0]), .Q(n24) );
  AO21X1 U48 ( .IN1(n2), .IN2(n41), .IN3(n25), .Q(n66) );
  MUX21X1 U49 ( .IN1(n78), .IN2(n26), .S(MdcEn_n), .Q(n25) );
  AO221X1 U50 ( .IN1(ByteSelect[0]), .IN2(n27), .IN3(Rgad[3]), .IN4(
        ByteSelect[1]), .IN5(n28), .Q(n26) );
  AO22X1 U51 ( .IN1(CtrlData[5]), .IN2(ByteSelect[3]), .IN3(CtrlData[13]), 
        .IN4(ByteSelect[2]), .Q(n28) );
  INVX0 U52 ( .INP(WriteOp), .ZN(n27) );
  MUX21X1 U53 ( .IN1(n40), .IN2(n29), .S(MdcEn_n), .Q(n64) );
  NAND4X0 U54 ( .IN1(n30), .IN2(n31), .IN3(n32), .IN4(n33), .QN(n29) );
  NAND2X0 U55 ( .IN1(CtrlData[14]), .IN2(ByteSelect[2]), .QN(n32) );
  NAND2X0 U56 ( .IN1(CtrlData[6]), .IN2(ByteSelect[3]), .QN(n31) );
  MUX21X1 U57 ( .IN1(n34), .IN2(n35), .S(ByteSelect[1]), .Q(n30) );
  INVX0 U58 ( .INP(Rgad[4]), .ZN(n35) );
  NAND2X0 U59 ( .IN1(n78), .IN2(n15), .QN(n34) );
  AO21X1 U60 ( .IN1(n2), .IN2(n40), .IN3(n36), .Q(n62) );
  MUX21X1 U61 ( .IN1(ShiftedBit), .IN2(n37), .S(MdcEn_n), .Q(n36) );
  AO222X1 U62 ( .IN1(CtrlData[15]), .IN2(ByteSelect[2]), .IN3(Fiad[0]), .IN4(
        ByteSelect[1]), .IN5(CtrlData[7]), .IN6(ByteSelect[3]), .Q(n37) );
  AND4X1 U63 ( .IN1(MdcEn_n), .IN2(n15), .IN3(n33), .IN4(n38), .Q(n2) );
  INVX0 U64 ( .INP(ByteSelect[1]), .ZN(n38) );
  INVX0 U65 ( .INP(ByteSelect[0]), .ZN(n33) );
  NOR2X0 U66 ( .IN1(ByteSelect[2]), .IN2(ByteSelect[3]), .QN(n15) );
endmodule


module eth_outputcontrol_test_1 ( Clk, Reset, InProgress, ShiftedBit, 
        BitCounter, WriteOp, NoPre, MdcEn_n, Mdo, MdoEn, 
        eth_top_test_point_11887_in, test_si, test_se );
  input [6:0] BitCounter;
  input Clk, Reset, InProgress, ShiftedBit, WriteOp, NoPre, MdcEn_n,
         eth_top_test_point_11887_in, test_si, test_se;
  output Mdo, MdoEn;
  wire   n25, n27, n29, n31, n33, n36, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15;

  SDFFARX1 MdoEn_2d_reg ( .D(n36), .SI(test_si), .SE(test_se), .CLK(Clk), 
        .RSTB(n15), .Q(n1) );
  SDFFARX1 MdoEn_d_reg ( .D(n33), .SI(n1), .SE(test_se), .CLK(Clk), .RSTB(n15), 
        .Q(n3) );
  SDFFARX1 MdoEn_reg ( .D(n31), .SI(n3), .SE(test_se), .CLK(Clk), .RSTB(n15), 
        .Q(MdoEn) );
  SDFFARX1 Mdo_2d_reg ( .D(n29), .SI(MdoEn), .SE(test_se), .CLK(Clk), .RSTB(
        n15), .Q(n2) );
  SDFFARX1 Mdo_d_reg ( .D(n27), .SI(n2), .SE(test_se), .CLK(Clk), .RSTB(n15), 
        .Q(n4) );
  SDFFARX1 Mdo_reg ( .D(n25), .SI(n4), .SE(test_se), .CLK(Clk), .RSTB(n15), 
        .Q(Mdo) );
  INVX0 U3 ( .INP(eth_top_test_point_11887_in), .ZN(n15) );
  MUX21X1 U4 ( .IN1(n1), .IN2(n5), .S(MdcEn_n), .Q(n36) );
  OA21X1 U5 ( .IN1(n6), .IN2(WriteOp), .IN3(InProgress), .Q(n5) );
  NOR2X0 U6 ( .IN1(BitCounter[6]), .IN2(n7), .QN(n6) );
  OA21X1 U7 ( .IN1(BitCounter[4]), .IN2(n8), .IN3(BitCounter[5]), .Q(n7) );
  AND3X1 U8 ( .IN1(BitCounter[2]), .IN2(BitCounter[1]), .IN3(BitCounter[3]), 
        .Q(n8) );
  MUX21X1 U9 ( .IN1(n3), .IN2(n1), .S(MdcEn_n), .Q(n33) );
  MUX21X1 U10 ( .IN1(MdoEn), .IN2(n3), .S(MdcEn_n), .Q(n31) );
  MUX21X1 U11 ( .IN1(n2), .IN2(n9), .S(MdcEn_n), .Q(n29) );
  NOR3X0 U12 ( .IN1(BitCounter[5]), .IN2(BitCounter[6]), .IN3(n10), .QN(n9) );
  AND3X1 U13 ( .IN1(n11), .IN2(NoPre), .IN3(n12), .Q(n10) );
  NOR4X0 U14 ( .IN1(BitCounter[4]), .IN2(BitCounter[3]), .IN3(BitCounter[2]), 
        .IN4(BitCounter[1]), .QN(n12) );
  NOR2X0 U15 ( .IN1(BitCounter[0]), .IN2(n13), .QN(n11) );
  INVX0 U16 ( .INP(InProgress), .ZN(n13) );
  MUX21X1 U17 ( .IN1(n4), .IN2(n14), .S(MdcEn_n), .Q(n27) );
  OR2X1 U18 ( .IN1(ShiftedBit), .IN2(n2), .Q(n14) );
  MUX21X1 U19 ( .IN1(Mdo), .IN2(n4), .S(MdcEn_n), .Q(n25) );
endmodule


module eth_miim_DW01_inc_0 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  XOR2X1 U2 ( .IN1(carry[6]), .IN2(A[6]), .Q(SUM[6]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module eth_miim_test_1 ( Clk, Reset, Divider, NoPre, CtrlData, Rgad, Fiad, 
        WCtrlData, RStat, ScanStat, Mdi, Mdo, MdoEn, Mdc, Busy, Prsd, LinkFail, 
        Nvalid, WCtrlDataStart, RStatStart, UpdateMIIRX_DATAReg, 
        eth_top_test_point_11887_in, test_si, test_so, test_se );
  input [7:0] Divider;
  input [15:0] CtrlData;
  input [4:0] Rgad;
  input [4:0] Fiad;
  output [15:0] Prsd;
  input Clk, Reset, NoPre, WCtrlData, RStat, ScanStat, Mdi,
         eth_top_test_point_11887_in, test_si, test_se;
  output Mdo, MdoEn, Mdc, Busy, LinkFail, Nvalid, WCtrlDataStart, RStatStart,
         UpdateMIIRX_DATAReg, test_so;
  wire   EndBusy_d, N9, WCtrlData_q1, RStat_q1, ScanStat_q1, MdcEn, RStat_q2,
         WCtrlData_q2, InProgress, WriteOp, N39, N40, N41, N42, N43, N44, N45,
         MdcEn_n, ShiftedBit, n49, n50, n51, n52, n53, n55, n58, n60, n64, n65,
         n66, n67, n68, n69, n70, n73, n75, n77, n79, n81, n83, n85, n87, n89,
         n91, n95, n100, n102, n105, n110, n112, n114, n117, n125, n133, n135,
         n136, n137, n138, n139, n140, n5, n6, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n54, n56, n94, n98, n101, n1, n2, n3, n4, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n57, n59, n61;
  wire   [1:0] LatchByte;
  wire   [6:0] BitCounter;
  wire   [3:0] ByteSelect;
  assign test_so = ShiftedBit;

  SDFFARX1 ScanStat_q1_reg ( .D(ScanStat), .SI(n50), .SE(test_se), .CLK(n1), 
        .RSTB(n61), .Q(ScanStat_q1) );
  SDFFARX1 ScanStat_q2_reg ( .D(ScanStat_q1), .SI(ScanStat_q1), .SE(test_se), 
        .CLK(n1), .RSTB(n61), .Q(n46), .QN(n6) );
  SDFFARX1 SyncStatMdcEn_reg ( .D(n125), .SI(n46), .SE(test_se), .CLK(n1), 
        .RSTB(n61), .Q(n45), .QN(n59) );
  SDFFARX1 RStat_q1_reg ( .D(RStat), .SI(RStatStart), .SE(test_se), .CLK(n1), 
        .RSTB(n61), .Q(RStat_q1) );
  SDFFARX1 RStat_q2_reg ( .D(RStat_q1), .SI(RStat_q1), .SE(test_se), .CLK(n1), 
        .RSTB(n61), .Q(RStat_q2), .QN(n49) );
  SDFFARX1 RStat_q3_reg ( .D(RStat_q2), .SI(RStat_q2), .SE(test_se), .CLK(n1), 
        .RSTB(n61), .Q(n50) );
  SDFFARX1 WCtrlData_q1_reg ( .D(WCtrlData), .SI(WCtrlDataStart), .SE(test_se), 
        .CLK(n1), .RSTB(n61), .Q(WCtrlData_q1) );
  SDFFARX1 WCtrlData_q2_reg ( .D(WCtrlData_q1), .SI(WCtrlData_q1), .SE(test_se), .CLK(n1), .RSTB(n61), .Q(WCtrlData_q2), .QN(n51) );
  SDFFARX1 WCtrlData_q3_reg ( .D(WCtrlData_q2), .SI(WCtrlData_q2), .SE(test_se), .CLK(n1), .RSTB(n61), .Q(n52) );
  SDFFARX1 \BitCounter_reg[0]  ( .D(n117), .SI(test_si), .SE(test_se), .CLK(n1), .RSTB(n61), .Q(BitCounter[0]), .QN(n70) );
  SDFFARX1 InProgress_reg ( .D(n140), .SI(n47), .SE(test_se), .CLK(n1), .RSTB(
        n61), .Q(InProgress), .QN(n69) );
  SDFFARX1 InProgress_q1_reg ( .D(n114), .SI(n56), .SE(test_se), .CLK(n1), 
        .RSTB(n61), .Q(n44) );
  SDFFARX1 InProgress_q2_reg ( .D(n112), .SI(n44), .SE(test_se), .CLK(n1), 
        .RSTB(n61), .Q(n43) );
  SDFFARX1 InProgress_q3_reg ( .D(n110), .SI(n43), .SE(test_se), .CLK(n1), 
        .RSTB(n61), .Q(n47), .QN(n57) );
  SDFFARX1 EndBusy_d_reg ( .D(n133), .SI(BitCounter[6]), .SE(test_se), .CLK(n1), .RSTB(n61), .Q(EndBusy_d) );
  SDFFARX1 EndBusy_reg ( .D(EndBusy_d), .SI(EndBusy_d), .SE(test_se), .CLK(n1), 
        .RSTB(n61), .Q(n56), .QN(n37) );
  SDFFARX1 WCtrlDataStart_reg ( .D(n137), .SI(n42), .SE(test_se), .CLK(n1), 
        .RSTB(n61), .Q(WCtrlDataStart), .QN(n60) );
  SDFFARX1 WCtrlDataStart_q_reg ( .D(n105), .SI(n48), .SE(test_se), .CLK(n1), 
        .RSTB(n61), .Q(n42) );
  SDFFARX1 UpdateMIIRX_DATAReg_reg ( .D(N9), .SI(n45), .SE(test_se), .CLK(n1), 
        .RSTB(n61), .Q(UpdateMIIRX_DATAReg) );
  SDFFARX1 WCtrlDataStart_q1_reg ( .D(n102), .SI(UpdateMIIRX_DATAReg), .SE(
        test_se), .CLK(n1), .RSTB(n61), .Q(n41), .QN(n36) );
  SDFFARX1 WCtrlDataStart_q2_reg ( .D(n100), .SI(n41), .SE(test_se), .CLK(n1), 
        .RSTB(n61), .Q(n48), .QN(n98) );
  SDFFARX1 RStatStart_reg ( .D(n138), .SI(n54), .SE(test_se), .CLK(n1), .RSTB(
        n61), .Q(RStatStart), .QN(n58) );
  SDFFARX1 RStatStart_q1_reg ( .D(n101), .SI(Nvalid), .SE(test_se), .CLK(n1), 
        .RSTB(n61), .Q(n40), .QN(n5) );
  SDFFARX1 RStatStart_q2_reg ( .D(n95), .SI(n40), .SE(test_se), .CLK(n1), 
        .RSTB(n61), .Q(n54), .QN(n94) );
  SDFFARX1 Nvalid_reg ( .D(n139), .SI(LatchByte[1]), .SE(test_se), .CLK(n1), 
        .RSTB(n61), .Q(Nvalid), .QN(n53) );
  SDFFARX1 WriteOp_reg ( .D(n136), .SI(n52), .SE(test_se), .CLK(n1), .RSTB(n61), .Q(WriteOp), .QN(n55) );
  SDFFARX1 \BitCounter_reg[5]  ( .D(n91), .SI(BitCounter[4]), .SE(test_se), 
        .CLK(n1), .RSTB(n61), .Q(BitCounter[5]), .QN(n68) );
  SDFFARX1 \BitCounter_reg[1]  ( .D(n89), .SI(BitCounter[0]), .SE(test_se), 
        .CLK(n1), .RSTB(n61), .Q(BitCounter[1]), .QN(n67) );
  SDFFARX1 \BitCounter_reg[2]  ( .D(n87), .SI(BitCounter[1]), .SE(test_se), 
        .CLK(n1), .RSTB(n61), .Q(BitCounter[2]), .QN(n66) );
  SDFFARX1 \BitCounter_reg[3]  ( .D(n85), .SI(BitCounter[2]), .SE(test_se), 
        .CLK(n1), .RSTB(n61), .Q(BitCounter[3]), .QN(n135) );
  SDFFARX1 \BitCounter_reg[4]  ( .D(n83), .SI(BitCounter[3]), .SE(test_se), 
        .CLK(n1), .RSTB(n61), .Q(BitCounter[4]), .QN(n64) );
  SDFFARX1 \BitCounter_reg[6]  ( .D(n81), .SI(BitCounter[5]), .SE(test_se), 
        .CLK(n1), .RSTB(n61), .Q(BitCounter[6]), .QN(n65) );
  SDFFARX1 LatchByte1_d_reg ( .D(n79), .SI(n38), .SE(test_se), .CLK(n1), 
        .RSTB(n61), .Q(n39) );
  SDFFARX1 \LatchByte_reg[1]  ( .D(n77), .SI(LatchByte[0]), .SE(test_se), 
        .CLK(n1), .RSTB(n61), .Q(LatchByte[1]) );
  SDFFARX1 LatchByte0_d_reg ( .D(n75), .SI(InProgress), .SE(test_se), .CLK(n1), 
        .RSTB(n61), .Q(n38) );
  SDFFARX1 \LatchByte_reg[0]  ( .D(n73), .SI(n39), .SE(test_se), .CLK(n1), 
        .RSTB(n61), .Q(LatchByte[0]) );
  eth_clockgen_test_1 clkgen ( .Clk(n1), .Reset(Reset), .Divider(Divider), 
        .MdcEn(MdcEn), .MdcEn_n(MdcEn_n), .Mdc(Mdc), 
        .eth_top_test_point_11887_in(eth_top_test_point_11887_in), .test_si(
        WriteOp), .test_se(test_se) );
  eth_shiftreg_test_1 shftrg ( .Clk(n1), .Reset(Reset), .MdcEn_n(MdcEn_n), 
        .Mdi(Mdi), .Fiad(Fiad), .Rgad(Rgad), .CtrlData(CtrlData), .WriteOp(
        WriteOp), .ByteSelect(ByteSelect), .LatchByte(LatchByte), .ShiftedBit(
        ShiftedBit), .Prsd(Prsd), .LinkFail(LinkFail), 
        .eth_top_test_point_11887_in(eth_top_test_point_11887_in), .test_si(
        Mdo), .test_se(test_se) );
  eth_outputcontrol_test_1 outctrl ( .Clk(n1), .Reset(Reset), .InProgress(
        InProgress), .ShiftedBit(ShiftedBit), .BitCounter(BitCounter), 
        .WriteOp(WriteOp), .NoPre(NoPre), .MdcEn_n(MdcEn_n), .Mdo(Mdo), 
        .MdoEn(MdoEn), .eth_top_test_point_11887_in(
        eth_top_test_point_11887_in), .test_si(Mdc), .test_se(test_se) );
  eth_miim_DW01_inc_0 add_412 ( .A(BitCounter), .SUM({N45, N44, N43, N42, N41, 
        N40, N39}) );
  INVX1 U3 ( .INP(eth_top_test_point_11887_in), .ZN(n61) );
  DELLN1X2 U4 ( .INP(Clk), .Z(n1) );
  INVX0 U5 ( .INP(n2), .ZN(n95) );
  MUX21X1 U6 ( .IN1(n5), .IN2(n94), .S(n3), .Q(n2) );
  OAI22X1 U7 ( .IN1(n68), .IN2(MdcEn), .IN3(n4), .IN4(n7), .QN(n91) );
  NOR2X0 U8 ( .IN1(n8), .IN2(N44), .QN(n4) );
  AO22X1 U9 ( .IN1(n3), .IN2(BitCounter[1]), .IN3(N40), .IN4(n9), .Q(n89) );
  AO22X1 U10 ( .IN1(n3), .IN2(BitCounter[2]), .IN3(N41), .IN4(n9), .Q(n87) );
  AO22X1 U11 ( .IN1(n3), .IN2(BitCounter[3]), .IN3(N42), .IN4(n9), .Q(n85) );
  AO22X1 U12 ( .IN1(n3), .IN2(BitCounter[4]), .IN3(N43), .IN4(n9), .Q(n83) );
  AO22X1 U13 ( .IN1(n3), .IN2(BitCounter[6]), .IN3(N45), .IN4(n9), .Q(n81) );
  NOR2X0 U14 ( .IN1(n7), .IN2(n8), .QN(n9) );
  AO22X1 U15 ( .IN1(n3), .IN2(n39), .IN3(n10), .IN4(n135), .Q(n79) );
  MUX21X1 U16 ( .IN1(n39), .IN2(LatchByte[1]), .S(n3), .Q(n77) );
  AO22X1 U17 ( .IN1(n3), .IN2(n38), .IN3(n10), .IN4(BitCounter[3]), .Q(n75) );
  AND3X1 U18 ( .IN1(n11), .IN2(n12), .IN3(n55), .Q(n10) );
  MUX21X1 U19 ( .IN1(n38), .IN2(LatchByte[0]), .S(n3), .Q(n73) );
  AO22X1 U20 ( .IN1(MdcEn), .IN2(n13), .IN3(n14), .IN4(InProgress), .Q(n140)
         );
  OR2X1 U21 ( .IN1(n15), .IN2(n3), .Q(n14) );
  NOR2X0 U22 ( .IN1(n133), .IN2(n16), .QN(n139) );
  OA21X1 U23 ( .IN1(n6), .IN2(n45), .IN3(n53), .Q(n16) );
  NOR2X0 U24 ( .IN1(n17), .IN2(n56), .QN(n138) );
  OA21X1 U25 ( .IN1(n49), .IN2(n50), .IN3(n58), .Q(n17) );
  NOR2X0 U26 ( .IN1(n18), .IN2(n56), .QN(n137) );
  OA21X1 U27 ( .IN1(n51), .IN2(n52), .IN3(n60), .Q(n18) );
  MUX21X1 U28 ( .IN1(WriteOp), .IN2(n19), .S(n20), .Q(n136) );
  NOR2X0 U29 ( .IN1(n21), .IN2(n3), .QN(n20) );
  OA21X1 U30 ( .IN1(n22), .IN2(InProgress), .IN3(n15), .Q(n21) );
  NAND3X0 U31 ( .IN1(n11), .IN2(BitCounter[3]), .IN3(n22), .QN(n15) );
  AND4X1 U32 ( .IN1(BitCounter[4]), .IN2(BitCounter[2]), .IN3(n65), .IN4(n23), 
        .Q(n11) );
  NOR3X0 U33 ( .IN1(n67), .IN2(n70), .IN3(n68), .QN(n23) );
  INVX0 U34 ( .INP(n13), .ZN(n22) );
  AO221X1 U35 ( .IN1(n94), .IN2(n40), .IN3(n98), .IN4(n41), .IN5(n24), .Q(n13)
         );
  NOR4X0 U36 ( .IN1(n59), .IN2(InProgress), .IN3(n44), .IN4(n43), .QN(n24) );
  NOR2X0 U37 ( .IN1(n36), .IN2(n48), .QN(n19) );
  NOR2X0 U38 ( .IN1(n43), .IN2(n57), .QN(n133) );
  INVX0 U39 ( .INP(n25), .ZN(n125) );
  MUX21X1 U40 ( .IN1(n6), .IN2(n59), .S(n3), .Q(n25) );
  OAI22X1 U41 ( .IN1(n70), .IN2(MdcEn), .IN3(n26), .IN4(n7), .QN(n117) );
  INVX0 U42 ( .INP(n12), .ZN(n7) );
  NOR2X0 U43 ( .IN1(n8), .IN2(N39), .QN(n26) );
  INVX0 U44 ( .INP(n27), .ZN(n8) );
  AO21X1 U45 ( .IN1(n3), .IN2(n44), .IN3(n12), .Q(n114) );
  NOR2X0 U46 ( .IN1(n3), .IN2(n69), .QN(n12) );
  MUX21X1 U47 ( .IN1(n44), .IN2(n43), .S(n3), .Q(n112) );
  MUX21X1 U48 ( .IN1(n43), .IN2(n47), .S(n3), .Q(n110) );
  MUX21X1 U49 ( .IN1(WCtrlDataStart), .IN2(n42), .S(n56), .Q(n105) );
  MUX21X1 U50 ( .IN1(WCtrlDataStart), .IN2(n41), .S(n3), .Q(n102) );
  MUX21X1 U51 ( .IN1(RStatStart), .IN2(n40), .S(n3), .Q(n101) );
  MUX21X1 U52 ( .IN1(n41), .IN2(n48), .S(n3), .Q(n100) );
  INVX0 U53 ( .INP(MdcEn), .ZN(n3) );
  NOR2X0 U54 ( .IN1(n37), .IN2(n42), .QN(N9) );
  NOR2X0 U55 ( .IN1(n135), .IN2(n28), .QN(ByteSelect[3]) );
  NOR2X0 U56 ( .IN1(BitCounter[3]), .IN2(n28), .QN(ByteSelect[2]) );
  NAND3X0 U57 ( .IN1(WriteOp), .IN2(BitCounter[4]), .IN3(n29), .QN(n28) );
  AND3X1 U58 ( .IN1(n64), .IN2(BitCounter[3]), .IN3(n29), .Q(ByteSelect[1]) );
  OAI21X1 U59 ( .IN1(n69), .IN2(n27), .IN3(n30), .QN(ByteSelect[0]) );
  NAND4X0 U60 ( .IN1(n29), .IN2(n64), .IN3(n135), .IN4(n31), .QN(n30) );
  NOR3X0 U61 ( .IN1(n68), .IN2(n69), .IN3(n32), .QN(n29) );
  NAND4X0 U62 ( .IN1(n68), .IN2(n64), .IN3(n33), .IN4(n135), .QN(n27) );
  NOR2X0 U63 ( .IN1(n32), .IN2(n31), .QN(n33) );
  INVX0 U64 ( .INP(NoPre), .ZN(n31) );
  NAND4X0 U65 ( .IN1(n70), .IN2(n67), .IN3(n66), .IN4(n65), .QN(n32) );
  NAND4X0 U66 ( .IN1(n53), .IN2(n59), .IN3(n34), .IN4(n35), .QN(Busy) );
  NOR4X0 U67 ( .IN1(RStatStart), .IN2(n56), .IN3(WCtrlDataStart), .IN4(n47), 
        .QN(n35) );
  NOR3X0 U68 ( .IN1(InProgress), .IN2(WCtrlData), .IN3(RStat), .QN(n34) );
endmodule


module eth_register_8_00_test_0 ( DataIn, DataOut, Write, Clk, Reset, 
        SyncReset, eth_top_test_point_11887_in, test_si, test_se );
  input [7:0] DataIn;
  output [7:0] DataOut;
  input Write, Clk, Reset, SyncReset, eth_top_test_point_11887_in, test_si,
         test_se;
  wire   n13, n14, n15, n16, n17, n18, n19, n20, n1, n2, n3, n4;

  SDFFARX1 \DataOut_reg[7]  ( .D(n20), .SI(DataOut[6]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[7]) );
  SDFFARX1 \DataOut_reg[6]  ( .D(n19), .SI(DataOut[5]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[6]) );
  SDFFARX1 \DataOut_reg[5]  ( .D(n18), .SI(DataOut[4]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[5]) );
  SDFFARX1 \DataOut_reg[4]  ( .D(n17), .SI(DataOut[3]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[4]) );
  SDFFARX1 \DataOut_reg[3]  ( .D(n16), .SI(DataOut[2]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[3]) );
  SDFFARX1 \DataOut_reg[2]  ( .D(n15), .SI(DataOut[1]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[2]) );
  SDFFARX1 \DataOut_reg[1]  ( .D(n14), .SI(DataOut[0]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[1]) );
  SDFFARX1 \DataOut_reg[0]  ( .D(n13), .SI(test_si), .SE(test_se), .CLK(Clk), 
        .RSTB(n4), .Q(DataOut[0]) );
  INVX0 U2 ( .INP(eth_top_test_point_11887_in), .ZN(n4) );
  AO22X1 U3 ( .IN1(DataIn[7]), .IN2(n1), .IN3(n2), .IN4(DataOut[7]), .Q(n20)
         );
  AO22X1 U4 ( .IN1(DataIn[6]), .IN2(n1), .IN3(n2), .IN4(DataOut[6]), .Q(n19)
         );
  AO22X1 U5 ( .IN1(DataIn[5]), .IN2(n1), .IN3(n2), .IN4(DataOut[5]), .Q(n18)
         );
  AO22X1 U6 ( .IN1(DataIn[4]), .IN2(n1), .IN3(n2), .IN4(DataOut[4]), .Q(n17)
         );
  AO22X1 U7 ( .IN1(DataIn[3]), .IN2(n1), .IN3(n2), .IN4(DataOut[3]), .Q(n16)
         );
  AO22X1 U8 ( .IN1(DataIn[2]), .IN2(n1), .IN3(n2), .IN4(DataOut[2]), .Q(n15)
         );
  AO22X1 U9 ( .IN1(DataIn[1]), .IN2(n1), .IN3(n2), .IN4(DataOut[1]), .Q(n14)
         );
  AO22X1 U10 ( .IN1(DataIn[0]), .IN2(n1), .IN3(n2), .IN4(DataOut[0]), .Q(n13)
         );
  NOR2X0 U11 ( .IN1(n1), .IN2(SyncReset), .QN(n2) );
  NOR2X0 U12 ( .IN1(n3), .IN2(SyncReset), .QN(n1) );
  INVX0 U13 ( .INP(Write), .ZN(n3) );
endmodule


module eth_register_8_a0_test_1 ( DataIn, DataOut, Write, Clk, Reset, 
        SyncReset, eth_top_test_point_11887_in, test_si, test_se );
  input [7:0] DataIn;
  output [7:0] DataOut;
  input Write, Clk, Reset, SyncReset, eth_top_test_point_11887_in, test_si,
         test_se;
  wire   n13, n14, n15, n16, n17, n18, n19, n20, n1, n2, n3, n4;

  SDFFASX1 \DataOut_reg[7]  ( .D(n20), .SI(DataOut[6]), .SE(test_se), .CLK(Clk), .SETB(n4), .Q(DataOut[7]) );
  SDFFARX1 \DataOut_reg[6]  ( .D(n19), .SI(DataOut[5]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[6]) );
  SDFFASX1 \DataOut_reg[5]  ( .D(n18), .SI(DataOut[4]), .SE(test_se), .CLK(Clk), .SETB(n4), .Q(DataOut[5]) );
  SDFFARX1 \DataOut_reg[4]  ( .D(n17), .SI(DataOut[3]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[4]) );
  SDFFARX1 \DataOut_reg[3]  ( .D(n16), .SI(DataOut[2]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[3]) );
  SDFFARX1 \DataOut_reg[2]  ( .D(n15), .SI(DataOut[1]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[2]) );
  SDFFARX1 \DataOut_reg[1]  ( .D(n14), .SI(DataOut[0]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[1]) );
  SDFFARX1 \DataOut_reg[0]  ( .D(n13), .SI(test_si), .SE(test_se), .CLK(Clk), 
        .RSTB(n4), .Q(DataOut[0]) );
  INVX0 U3 ( .INP(eth_top_test_point_11887_in), .ZN(n4) );
  AO221X1 U4 ( .IN1(n1), .IN2(DataOut[7]), .IN3(DataIn[7]), .IN4(n2), .IN5(
        SyncReset), .Q(n20) );
  AO22X1 U5 ( .IN1(DataIn[6]), .IN2(n2), .IN3(n1), .IN4(DataOut[6]), .Q(n19)
         );
  AO221X1 U6 ( .IN1(n1), .IN2(DataOut[5]), .IN3(DataIn[5]), .IN4(n2), .IN5(
        SyncReset), .Q(n18) );
  AO22X1 U7 ( .IN1(DataIn[4]), .IN2(n2), .IN3(n1), .IN4(DataOut[4]), .Q(n17)
         );
  AO22X1 U8 ( .IN1(DataIn[3]), .IN2(n2), .IN3(n1), .IN4(DataOut[3]), .Q(n16)
         );
  AO22X1 U9 ( .IN1(DataIn[2]), .IN2(n2), .IN3(n1), .IN4(DataOut[2]), .Q(n15)
         );
  AO22X1 U10 ( .IN1(DataIn[1]), .IN2(n2), .IN3(n1), .IN4(DataOut[1]), .Q(n14)
         );
  AO22X1 U11 ( .IN1(DataIn[0]), .IN2(n2), .IN3(n1), .IN4(DataOut[0]), .Q(n13)
         );
  NOR2X0 U12 ( .IN1(n2), .IN2(SyncReset), .QN(n1) );
  NOR2X0 U13 ( .IN1(n3), .IN2(SyncReset), .QN(n2) );
  INVX0 U14 ( .INP(Write), .ZN(n3) );
endmodule


module eth_register_1_0_test_0 ( DataIn, DataOut, Write, Clk, Reset, SyncReset, 
        eth_top_test_point_11887_in, test_si, test_se );
  input [0:0] DataIn;
  output [0:0] DataOut;
  input Write, Clk, Reset, SyncReset, eth_top_test_point_11887_in, test_si,
         test_se;
  wire   n5, n1, n2, n3;

  SDFFARX1 \DataOut_reg[0]  ( .D(n5), .SI(test_si), .SE(test_se), .CLK(Clk), 
        .RSTB(n3), .Q(DataOut[0]) );
  INVX0 U2 ( .INP(eth_top_test_point_11887_in), .ZN(n3) );
  NOR2X0 U3 ( .IN1(SyncReset), .IN2(n1), .QN(n5) );
  INVX0 U4 ( .INP(n2), .ZN(n1) );
  MUX21X1 U5 ( .IN1(DataOut[0]), .IN2(DataIn[0]), .S(Write), .Q(n2) );
endmodule


module eth_register_7_00_test_1 ( DataIn, DataOut, Write, Clk, Reset, 
        SyncReset, eth_top_test_point_11887_in, test_si, test_se );
  input [6:0] DataIn;
  output [6:0] DataOut;
  input Write, Clk, Reset, SyncReset, eth_top_test_point_11887_in, test_si,
         test_se;
  wire   n12, n13, n14, n15, n16, n17, n18, n1, n2, n3, n4;

  SDFFARX1 \DataOut_reg[6]  ( .D(n18), .SI(DataOut[5]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[6]) );
  SDFFARX1 \DataOut_reg[5]  ( .D(n17), .SI(DataOut[4]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[5]) );
  SDFFARX1 \DataOut_reg[4]  ( .D(n16), .SI(DataOut[3]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[4]) );
  SDFFARX1 \DataOut_reg[3]  ( .D(n15), .SI(DataOut[2]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[3]) );
  SDFFARX1 \DataOut_reg[2]  ( .D(n14), .SI(DataOut[1]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[2]) );
  SDFFARX1 \DataOut_reg[1]  ( .D(n13), .SI(DataOut[0]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[1]) );
  SDFFARX1 \DataOut_reg[0]  ( .D(n12), .SI(test_si), .SE(test_se), .CLK(Clk), 
        .RSTB(n4), .Q(DataOut[0]) );
  INVX0 U2 ( .INP(eth_top_test_point_11887_in), .ZN(n4) );
  AO22X1 U3 ( .IN1(DataIn[6]), .IN2(n1), .IN3(n2), .IN4(DataOut[6]), .Q(n18)
         );
  AO22X1 U4 ( .IN1(DataIn[5]), .IN2(n1), .IN3(n2), .IN4(DataOut[5]), .Q(n17)
         );
  AO22X1 U5 ( .IN1(DataIn[4]), .IN2(n1), .IN3(n2), .IN4(DataOut[4]), .Q(n16)
         );
  AO22X1 U6 ( .IN1(DataIn[3]), .IN2(n1), .IN3(n2), .IN4(DataOut[3]), .Q(n15)
         );
  AO22X1 U7 ( .IN1(DataIn[2]), .IN2(n1), .IN3(n2), .IN4(DataOut[2]), .Q(n14)
         );
  AO22X1 U8 ( .IN1(DataIn[1]), .IN2(n1), .IN3(n2), .IN4(DataOut[1]), .Q(n13)
         );
  AO22X1 U9 ( .IN1(DataIn[0]), .IN2(n1), .IN3(n2), .IN4(DataOut[0]), .Q(n12)
         );
  NOR2X0 U10 ( .IN1(n1), .IN2(SyncReset), .QN(n2) );
  NOR2X0 U11 ( .IN1(n3), .IN2(SyncReset), .QN(n1) );
  INVX0 U12 ( .INP(Write), .ZN(n3) );
endmodule


module eth_register_7_12_test_0 ( DataIn, DataOut, Write, Clk, Reset, 
        SyncReset, eth_top_test_point_11887_in, test_si, test_se );
  input [6:0] DataIn;
  output [6:0] DataOut;
  input Write, Clk, Reset, SyncReset, eth_top_test_point_11887_in, test_si,
         test_se;
  wire   n12, n13, n14, n15, n16, n17, n18, n1, n2, n3, n4;

  SDFFARX1 \DataOut_reg[6]  ( .D(n18), .SI(DataOut[5]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[6]) );
  SDFFARX1 \DataOut_reg[5]  ( .D(n17), .SI(DataOut[4]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[5]) );
  SDFFASX1 \DataOut_reg[4]  ( .D(n16), .SI(DataOut[3]), .SE(test_se), .CLK(Clk), .SETB(n4), .Q(DataOut[4]) );
  SDFFARX1 \DataOut_reg[3]  ( .D(n15), .SI(DataOut[2]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[3]) );
  SDFFARX1 \DataOut_reg[2]  ( .D(n14), .SI(DataOut[1]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[2]) );
  SDFFASX1 \DataOut_reg[1]  ( .D(n13), .SI(DataOut[0]), .SE(test_se), .CLK(Clk), .SETB(n4), .Q(DataOut[1]) );
  SDFFARX1 \DataOut_reg[0]  ( .D(n12), .SI(test_si), .SE(test_se), .CLK(Clk), 
        .RSTB(n4), .Q(DataOut[0]) );
  INVX0 U3 ( .INP(eth_top_test_point_11887_in), .ZN(n4) );
  AO22X1 U4 ( .IN1(DataIn[6]), .IN2(n1), .IN3(n2), .IN4(DataOut[6]), .Q(n18)
         );
  AO22X1 U5 ( .IN1(DataIn[5]), .IN2(n1), .IN3(n2), .IN4(DataOut[5]), .Q(n17)
         );
  AO221X1 U6 ( .IN1(n2), .IN2(DataOut[4]), .IN3(DataIn[4]), .IN4(n1), .IN5(
        SyncReset), .Q(n16) );
  AO22X1 U7 ( .IN1(DataIn[3]), .IN2(n1), .IN3(n2), .IN4(DataOut[3]), .Q(n15)
         );
  AO22X1 U8 ( .IN1(DataIn[2]), .IN2(n1), .IN3(n2), .IN4(DataOut[2]), .Q(n14)
         );
  AO221X1 U9 ( .IN1(n2), .IN2(DataOut[1]), .IN3(DataIn[1]), .IN4(n1), .IN5(
        SyncReset), .Q(n13) );
  AO22X1 U10 ( .IN1(DataIn[0]), .IN2(n1), .IN3(n2), .IN4(DataOut[0]), .Q(n12)
         );
  NOR2X0 U11 ( .IN1(n1), .IN2(SyncReset), .QN(n2) );
  NOR2X0 U12 ( .IN1(n3), .IN2(SyncReset), .QN(n1) );
  INVX0 U13 ( .INP(Write), .ZN(n3) );
endmodule


module eth_register_7_0c_test_1 ( DataIn, DataOut, Write, Clk, Reset, 
        SyncReset, eth_top_test_point_11887_in, test_si, test_se );
  input [6:0] DataIn;
  output [6:0] DataOut;
  input Write, Clk, Reset, SyncReset, eth_top_test_point_11887_in, test_si,
         test_se;
  wire   n12, n13, n14, n15, n16, n17, n18, n1, n2, n3, n4;

  SDFFARX1 \DataOut_reg[6]  ( .D(n18), .SI(DataOut[5]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[6]) );
  SDFFARX1 \DataOut_reg[5]  ( .D(n17), .SI(DataOut[4]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[5]) );
  SDFFARX1 \DataOut_reg[4]  ( .D(n16), .SI(DataOut[3]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[4]) );
  SDFFASX1 \DataOut_reg[3]  ( .D(n15), .SI(DataOut[2]), .SE(test_se), .CLK(Clk), .SETB(n4), .Q(DataOut[3]) );
  SDFFASX1 \DataOut_reg[2]  ( .D(n14), .SI(DataOut[1]), .SE(test_se), .CLK(Clk), .SETB(n4), .Q(DataOut[2]) );
  SDFFARX1 \DataOut_reg[1]  ( .D(n13), .SI(DataOut[0]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[1]) );
  SDFFARX1 \DataOut_reg[0]  ( .D(n12), .SI(test_si), .SE(test_se), .CLK(Clk), 
        .RSTB(n4), .Q(DataOut[0]) );
  INVX0 U3 ( .INP(eth_top_test_point_11887_in), .ZN(n4) );
  AO22X1 U4 ( .IN1(DataIn[6]), .IN2(n1), .IN3(n2), .IN4(DataOut[6]), .Q(n18)
         );
  AO22X1 U5 ( .IN1(DataIn[5]), .IN2(n1), .IN3(n2), .IN4(DataOut[5]), .Q(n17)
         );
  AO22X1 U6 ( .IN1(DataIn[4]), .IN2(n1), .IN3(n2), .IN4(DataOut[4]), .Q(n16)
         );
  AO221X1 U7 ( .IN1(n2), .IN2(DataOut[3]), .IN3(DataIn[3]), .IN4(n1), .IN5(
        SyncReset), .Q(n15) );
  AO221X1 U8 ( .IN1(n2), .IN2(DataOut[2]), .IN3(DataIn[2]), .IN4(n1), .IN5(
        SyncReset), .Q(n14) );
  AO22X1 U9 ( .IN1(DataIn[1]), .IN2(n1), .IN3(n2), .IN4(DataOut[1]), .Q(n13)
         );
  AO22X1 U10 ( .IN1(DataIn[0]), .IN2(n1), .IN3(n2), .IN4(DataOut[0]), .Q(n12)
         );
  NOR2X0 U11 ( .IN1(n1), .IN2(SyncReset), .QN(n2) );
  NOR2X0 U12 ( .IN1(n3), .IN2(SyncReset), .QN(n1) );
  INVX0 U13 ( .INP(Write), .ZN(n3) );
endmodule


module eth_register_7_12_test_1 ( DataIn, DataOut, Write, Clk, Reset, 
        SyncReset, eth_top_test_point_11887_in, test_si, test_se );
  input [6:0] DataIn;
  output [6:0] DataOut;
  input Write, Clk, Reset, SyncReset, eth_top_test_point_11887_in, test_si,
         test_se;
  wire   n19, n20, n21, n22, n23, n24, n25, n1, n2, n3, n4;

  SDFFARX1 \DataOut_reg[6]  ( .D(n19), .SI(DataOut[5]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[6]) );
  SDFFARX1 \DataOut_reg[5]  ( .D(n20), .SI(DataOut[4]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[5]) );
  SDFFASX1 \DataOut_reg[4]  ( .D(n21), .SI(DataOut[3]), .SE(test_se), .CLK(Clk), .SETB(n4), .Q(DataOut[4]) );
  SDFFARX1 \DataOut_reg[3]  ( .D(n22), .SI(DataOut[2]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[3]) );
  SDFFARX1 \DataOut_reg[2]  ( .D(n23), .SI(DataOut[1]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[2]) );
  SDFFASX1 \DataOut_reg[1]  ( .D(n24), .SI(DataOut[0]), .SE(test_se), .CLK(Clk), .SETB(n4), .Q(DataOut[1]) );
  SDFFARX1 \DataOut_reg[0]  ( .D(n25), .SI(test_si), .SE(test_se), .CLK(Clk), 
        .RSTB(n4), .Q(DataOut[0]) );
  INVX0 U3 ( .INP(eth_top_test_point_11887_in), .ZN(n4) );
  AO22X1 U4 ( .IN1(DataIn[0]), .IN2(n1), .IN3(n2), .IN4(DataOut[0]), .Q(n25)
         );
  AO221X1 U5 ( .IN1(n2), .IN2(DataOut[1]), .IN3(DataIn[1]), .IN4(n1), .IN5(
        SyncReset), .Q(n24) );
  AO22X1 U6 ( .IN1(DataIn[2]), .IN2(n1), .IN3(n2), .IN4(DataOut[2]), .Q(n23)
         );
  AO22X1 U7 ( .IN1(DataIn[3]), .IN2(n1), .IN3(n2), .IN4(DataOut[3]), .Q(n22)
         );
  AO221X1 U8 ( .IN1(n2), .IN2(DataOut[4]), .IN3(DataIn[4]), .IN4(n1), .IN5(
        SyncReset), .Q(n21) );
  AO22X1 U9 ( .IN1(DataIn[5]), .IN2(n1), .IN3(n2), .IN4(DataOut[5]), .Q(n20)
         );
  AO22X1 U10 ( .IN1(DataIn[6]), .IN2(n1), .IN3(n2), .IN4(DataOut[6]), .Q(n19)
         );
  NOR2X0 U11 ( .IN1(n1), .IN2(SyncReset), .QN(n2) );
  NOR2X0 U12 ( .IN1(n3), .IN2(SyncReset), .QN(n1) );
  INVX0 U13 ( .INP(Write), .ZN(n3) );
endmodule


module eth_register_8_00_test_20 ( DataIn, DataOut, Write, Clk, Reset, 
        SyncReset, eth_top_test_point_11887_in, test_si, test_se );
  input [7:0] DataIn;
  output [7:0] DataOut;
  input Write, Clk, Reset, SyncReset, eth_top_test_point_11887_in, test_si,
         test_se;
  wire   n21, n22, n23, n24, n25, n26, n27, n28, n1, n2, n3, n4;

  SDFFARX1 \DataOut_reg[7]  ( .D(n21), .SI(DataOut[6]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[7]) );
  SDFFARX1 \DataOut_reg[6]  ( .D(n22), .SI(DataOut[5]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[6]) );
  SDFFARX1 \DataOut_reg[5]  ( .D(n23), .SI(DataOut[4]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[5]) );
  SDFFARX1 \DataOut_reg[4]  ( .D(n24), .SI(DataOut[3]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[4]) );
  SDFFARX1 \DataOut_reg[3]  ( .D(n25), .SI(DataOut[2]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[3]) );
  SDFFARX1 \DataOut_reg[2]  ( .D(n26), .SI(DataOut[1]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[2]) );
  SDFFARX1 \DataOut_reg[1]  ( .D(n27), .SI(DataOut[0]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[1]) );
  SDFFARX1 \DataOut_reg[0]  ( .D(n28), .SI(test_si), .SE(test_se), .CLK(Clk), 
        .RSTB(n4), .Q(DataOut[0]) );
  INVX0 U2 ( .INP(eth_top_test_point_11887_in), .ZN(n4) );
  AO22X1 U3 ( .IN1(DataIn[0]), .IN2(n1), .IN3(n2), .IN4(DataOut[0]), .Q(n28)
         );
  AO22X1 U4 ( .IN1(DataIn[1]), .IN2(n1), .IN3(n2), .IN4(DataOut[1]), .Q(n27)
         );
  AO22X1 U5 ( .IN1(DataIn[2]), .IN2(n1), .IN3(n2), .IN4(DataOut[2]), .Q(n26)
         );
  AO22X1 U6 ( .IN1(DataIn[3]), .IN2(n1), .IN3(n2), .IN4(DataOut[3]), .Q(n25)
         );
  AO22X1 U7 ( .IN1(DataIn[4]), .IN2(n1), .IN3(n2), .IN4(DataOut[4]), .Q(n24)
         );
  AO22X1 U8 ( .IN1(DataIn[5]), .IN2(n1), .IN3(n2), .IN4(DataOut[5]), .Q(n23)
         );
  AO22X1 U9 ( .IN1(DataIn[6]), .IN2(n1), .IN3(n2), .IN4(DataOut[6]), .Q(n22)
         );
  AO22X1 U10 ( .IN1(DataIn[7]), .IN2(n1), .IN3(n2), .IN4(DataOut[7]), .Q(n21)
         );
  NOR2X0 U11 ( .IN1(n1), .IN2(SyncReset), .QN(n2) );
  NOR2X0 U12 ( .IN1(n3), .IN2(SyncReset), .QN(n1) );
  INVX0 U13 ( .INP(Write), .ZN(n3) );
endmodule


module eth_register_8_06_test_1 ( DataIn, DataOut, Write, Clk, Reset, 
        SyncReset, eth_top_test_point_11887_in, test_si, test_se );
  input [7:0] DataIn;
  output [7:0] DataOut;
  input Write, Clk, Reset, SyncReset, eth_top_test_point_11887_in, test_si,
         test_se;
  wire   n13, n14, n15, n16, n17, n18, n19, n20, n1, n2, n3, n4;

  SDFFARX1 \DataOut_reg[7]  ( .D(n20), .SI(DataOut[6]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[7]) );
  SDFFARX1 \DataOut_reg[6]  ( .D(n19), .SI(DataOut[5]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[6]) );
  SDFFARX1 \DataOut_reg[5]  ( .D(n18), .SI(DataOut[4]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[5]) );
  SDFFARX1 \DataOut_reg[4]  ( .D(n17), .SI(DataOut[3]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[4]) );
  SDFFARX1 \DataOut_reg[3]  ( .D(n16), .SI(DataOut[2]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[3]) );
  SDFFASX1 \DataOut_reg[2]  ( .D(n15), .SI(DataOut[1]), .SE(test_se), .CLK(Clk), .SETB(n4), .Q(DataOut[2]) );
  SDFFASX1 \DataOut_reg[1]  ( .D(n14), .SI(DataOut[0]), .SE(test_se), .CLK(Clk), .SETB(n4), .Q(DataOut[1]) );
  SDFFARX1 \DataOut_reg[0]  ( .D(n13), .SI(test_si), .SE(test_se), .CLK(Clk), 
        .RSTB(n4), .Q(DataOut[0]) );
  INVX0 U3 ( .INP(eth_top_test_point_11887_in), .ZN(n4) );
  AO22X1 U4 ( .IN1(DataIn[7]), .IN2(n1), .IN3(n2), .IN4(DataOut[7]), .Q(n20)
         );
  AO22X1 U5 ( .IN1(DataIn[6]), .IN2(n1), .IN3(n2), .IN4(DataOut[6]), .Q(n19)
         );
  AO22X1 U6 ( .IN1(DataIn[5]), .IN2(n1), .IN3(n2), .IN4(DataOut[5]), .Q(n18)
         );
  AO22X1 U7 ( .IN1(DataIn[4]), .IN2(n1), .IN3(n2), .IN4(DataOut[4]), .Q(n17)
         );
  AO22X1 U8 ( .IN1(DataIn[3]), .IN2(n1), .IN3(n2), .IN4(DataOut[3]), .Q(n16)
         );
  AO221X1 U9 ( .IN1(n2), .IN2(DataOut[2]), .IN3(DataIn[2]), .IN4(n1), .IN5(
        SyncReset), .Q(n15) );
  AO221X1 U10 ( .IN1(n2), .IN2(DataOut[1]), .IN3(DataIn[1]), .IN4(n1), .IN5(
        SyncReset), .Q(n14) );
  AO22X1 U11 ( .IN1(DataIn[0]), .IN2(n1), .IN3(n2), .IN4(DataOut[0]), .Q(n13)
         );
  NOR2X0 U12 ( .IN1(n1), .IN2(SyncReset), .QN(n2) );
  NOR2X0 U13 ( .IN1(n3), .IN2(SyncReset), .QN(n1) );
  INVX0 U14 ( .INP(Write), .ZN(n3) );
endmodule


module eth_register_8_40_test_0 ( DataIn, DataOut, Write, Clk, Reset, 
        SyncReset, eth_top_test_point_11887_in, test_si, test_se );
  input [7:0] DataIn;
  output [7:0] DataOut;
  input Write, Clk, Reset, SyncReset, eth_top_test_point_11887_in, test_si,
         test_se;
  wire   n13, n14, n15, n16, n17, n18, n19, n20, n1, n2, n3, n4;

  SDFFARX1 \DataOut_reg[7]  ( .D(n20), .SI(DataOut[6]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[7]) );
  SDFFASX1 \DataOut_reg[6]  ( .D(n19), .SI(DataOut[5]), .SE(test_se), .CLK(Clk), .SETB(n4), .Q(DataOut[6]) );
  SDFFARX1 \DataOut_reg[5]  ( .D(n18), .SI(DataOut[4]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[5]) );
  SDFFARX1 \DataOut_reg[4]  ( .D(n17), .SI(DataOut[3]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[4]) );
  SDFFARX1 \DataOut_reg[3]  ( .D(n16), .SI(DataOut[2]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[3]) );
  SDFFARX1 \DataOut_reg[2]  ( .D(n15), .SI(DataOut[1]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[2]) );
  SDFFARX1 \DataOut_reg[1]  ( .D(n14), .SI(DataOut[0]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[1]) );
  SDFFARX1 \DataOut_reg[0]  ( .D(n13), .SI(test_si), .SE(test_se), .CLK(Clk), 
        .RSTB(n4), .Q(DataOut[0]) );
  INVX0 U3 ( .INP(eth_top_test_point_11887_in), .ZN(n4) );
  AO22X1 U4 ( .IN1(DataIn[7]), .IN2(n1), .IN3(n2), .IN4(DataOut[7]), .Q(n20)
         );
  AO221X1 U5 ( .IN1(n2), .IN2(DataOut[6]), .IN3(DataIn[6]), .IN4(n1), .IN5(
        SyncReset), .Q(n19) );
  AO22X1 U6 ( .IN1(DataIn[5]), .IN2(n1), .IN3(n2), .IN4(DataOut[5]), .Q(n18)
         );
  AO22X1 U7 ( .IN1(DataIn[4]), .IN2(n1), .IN3(n2), .IN4(DataOut[4]), .Q(n17)
         );
  AO22X1 U8 ( .IN1(DataIn[3]), .IN2(n1), .IN3(n2), .IN4(DataOut[3]), .Q(n16)
         );
  AO22X1 U9 ( .IN1(DataIn[2]), .IN2(n1), .IN3(n2), .IN4(DataOut[2]), .Q(n15)
         );
  AO22X1 U10 ( .IN1(DataIn[1]), .IN2(n1), .IN3(n2), .IN4(DataOut[1]), .Q(n14)
         );
  AO22X1 U11 ( .IN1(DataIn[0]), .IN2(n1), .IN3(n2), .IN4(DataOut[0]), .Q(n13)
         );
  NOR2X0 U12 ( .IN1(n1), .IN2(SyncReset), .QN(n2) );
  NOR2X0 U13 ( .IN1(n3), .IN2(SyncReset), .QN(n1) );
  INVX0 U14 ( .INP(Write), .ZN(n3) );
endmodule


module eth_register_8_00_test_19 ( DataIn, DataOut, Write, Clk, Reset, 
        SyncReset, eth_top_test_point_11887_in, test_si, test_se );
  input [7:0] DataIn;
  output [7:0] DataOut;
  input Write, Clk, Reset, SyncReset, eth_top_test_point_11887_in, test_si,
         test_se;
  wire   n21, n22, n23, n24, n25, n26, n27, n28, n1, n2, n3, n4;

  SDFFARX1 \DataOut_reg[7]  ( .D(n21), .SI(DataOut[6]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[7]) );
  SDFFARX1 \DataOut_reg[6]  ( .D(n22), .SI(DataOut[5]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[6]) );
  SDFFARX1 \DataOut_reg[5]  ( .D(n23), .SI(DataOut[4]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[5]) );
  SDFFARX1 \DataOut_reg[4]  ( .D(n24), .SI(DataOut[3]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[4]) );
  SDFFARX1 \DataOut_reg[3]  ( .D(n25), .SI(DataOut[2]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[3]) );
  SDFFARX1 \DataOut_reg[2]  ( .D(n26), .SI(DataOut[1]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[2]) );
  SDFFARX1 \DataOut_reg[1]  ( .D(n27), .SI(DataOut[0]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[1]) );
  SDFFARX1 \DataOut_reg[0]  ( .D(n28), .SI(test_si), .SE(test_se), .CLK(Clk), 
        .RSTB(n4), .Q(DataOut[0]) );
  INVX0 U2 ( .INP(eth_top_test_point_11887_in), .ZN(n4) );
  AO22X1 U3 ( .IN1(DataIn[0]), .IN2(n1), .IN3(n2), .IN4(DataOut[0]), .Q(n28)
         );
  AO22X1 U4 ( .IN1(DataIn[1]), .IN2(n1), .IN3(n2), .IN4(DataOut[1]), .Q(n27)
         );
  AO22X1 U5 ( .IN1(DataIn[2]), .IN2(n1), .IN3(n2), .IN4(DataOut[2]), .Q(n26)
         );
  AO22X1 U6 ( .IN1(DataIn[3]), .IN2(n1), .IN3(n2), .IN4(DataOut[3]), .Q(n25)
         );
  AO22X1 U7 ( .IN1(DataIn[4]), .IN2(n1), .IN3(n2), .IN4(DataOut[4]), .Q(n24)
         );
  AO22X1 U8 ( .IN1(DataIn[5]), .IN2(n1), .IN3(n2), .IN4(DataOut[5]), .Q(n23)
         );
  AO22X1 U9 ( .IN1(DataIn[6]), .IN2(n1), .IN3(n2), .IN4(DataOut[6]), .Q(n22)
         );
  AO22X1 U10 ( .IN1(DataIn[7]), .IN2(n1), .IN3(n2), .IN4(DataOut[7]), .Q(n21)
         );
  NOR2X0 U11 ( .IN1(n1), .IN2(SyncReset), .QN(n2) );
  NOR2X0 U12 ( .IN1(n3), .IN2(SyncReset), .QN(n1) );
  INVX0 U13 ( .INP(Write), .ZN(n3) );
endmodule


module eth_register_6_3f_test_1 ( DataIn, DataOut, Write, Clk, Reset, 
        SyncReset, eth_top_test_point_11887_in, test_si, test_se );
  input [5:0] DataIn;
  output [5:0] DataOut;
  input Write, Clk, Reset, SyncReset, eth_top_test_point_11887_in, test_si,
         test_se;
  wire   n9, n10, n11, n12, n13, n14, n1, n2, n3, n4, n5, n6, n7;

  SDFFASX1 \DataOut_reg[5]  ( .D(n14), .SI(DataOut[4]), .SE(test_se), .CLK(Clk), .SETB(n7), .Q(DataOut[5]) );
  SDFFASX1 \DataOut_reg[4]  ( .D(n13), .SI(DataOut[3]), .SE(test_se), .CLK(Clk), .SETB(n7), .Q(DataOut[4]) );
  SDFFASX1 \DataOut_reg[3]  ( .D(n12), .SI(DataOut[2]), .SE(test_se), .CLK(Clk), .SETB(n7), .Q(DataOut[3]) );
  SDFFASX1 \DataOut_reg[2]  ( .D(n11), .SI(DataOut[1]), .SE(test_se), .CLK(Clk), .SETB(n7), .Q(DataOut[2]) );
  SDFFASX1 \DataOut_reg[1]  ( .D(n10), .SI(DataOut[0]), .SE(test_se), .CLK(Clk), .SETB(n7), .Q(DataOut[1]) );
  SDFFASX1 \DataOut_reg[0]  ( .D(n9), .SI(test_si), .SE(test_se), .CLK(Clk), 
        .SETB(n7), .Q(DataOut[0]) );
  INVX0 U3 ( .INP(eth_top_test_point_11887_in), .ZN(n7) );
  OR2X1 U4 ( .IN1(SyncReset), .IN2(n1), .Q(n9) );
  MUX21X1 U5 ( .IN1(DataOut[0]), .IN2(DataIn[0]), .S(Write), .Q(n1) );
  OR2X1 U6 ( .IN1(SyncReset), .IN2(n2), .Q(n14) );
  MUX21X1 U7 ( .IN1(DataOut[5]), .IN2(DataIn[5]), .S(Write), .Q(n2) );
  OR2X1 U8 ( .IN1(SyncReset), .IN2(n3), .Q(n13) );
  MUX21X1 U9 ( .IN1(DataOut[4]), .IN2(DataIn[4]), .S(Write), .Q(n3) );
  OR2X1 U10 ( .IN1(SyncReset), .IN2(n4), .Q(n12) );
  MUX21X1 U11 ( .IN1(DataOut[3]), .IN2(DataIn[3]), .S(Write), .Q(n4) );
  OR2X1 U12 ( .IN1(SyncReset), .IN2(n5), .Q(n11) );
  MUX21X1 U13 ( .IN1(DataOut[2]), .IN2(DataIn[2]), .S(Write), .Q(n5) );
  OR2X1 U14 ( .IN1(SyncReset), .IN2(n6), .Q(n10) );
  MUX21X1 U15 ( .IN1(DataOut[1]), .IN2(DataIn[1]), .S(Write), .Q(n6) );
endmodule


module eth_register_4_f_test_1 ( DataIn, DataOut, Write, Clk, Reset, SyncReset, 
        eth_top_test_point_11887_in, test_si, test_se );
  input [3:0] DataIn;
  output [3:0] DataOut;
  input Write, Clk, Reset, SyncReset, eth_top_test_point_11887_in, test_si,
         test_se;
  wire   n7, n8, n9, n10, n1, n2, n3, n4, n5;

  SDFFASX1 \DataOut_reg[3]  ( .D(n10), .SI(DataOut[2]), .SE(test_se), .CLK(Clk), .SETB(n5), .Q(DataOut[3]) );
  SDFFASX1 \DataOut_reg[2]  ( .D(n9), .SI(DataOut[1]), .SE(test_se), .CLK(Clk), 
        .SETB(n5), .Q(DataOut[2]) );
  SDFFASX1 \DataOut_reg[1]  ( .D(n8), .SI(DataOut[0]), .SE(test_se), .CLK(Clk), 
        .SETB(n5), .Q(DataOut[1]) );
  SDFFASX1 \DataOut_reg[0]  ( .D(n7), .SI(test_si), .SE(test_se), .CLK(Clk), 
        .SETB(n5), .Q(DataOut[0]) );
  INVX0 U3 ( .INP(eth_top_test_point_11887_in), .ZN(n5) );
  OR2X1 U4 ( .IN1(SyncReset), .IN2(n1), .Q(n9) );
  MUX21X1 U5 ( .IN1(DataOut[2]), .IN2(DataIn[2]), .S(Write), .Q(n1) );
  OR2X1 U6 ( .IN1(SyncReset), .IN2(n2), .Q(n8) );
  MUX21X1 U7 ( .IN1(DataOut[1]), .IN2(DataIn[1]), .S(Write), .Q(n2) );
  OR2X1 U8 ( .IN1(SyncReset), .IN2(n3), .Q(n7) );
  MUX21X1 U9 ( .IN1(DataOut[0]), .IN2(DataIn[0]), .S(Write), .Q(n3) );
  OR2X1 U10 ( .IN1(SyncReset), .IN2(n4), .Q(n10) );
  MUX21X1 U11 ( .IN1(DataOut[3]), .IN2(DataIn[3]), .S(Write), .Q(n4) );
endmodule


module eth_register_8_40_test_1 ( DataIn, DataOut, Write, Clk, Reset, 
        SyncReset, eth_top_test_point_11887_in, test_si, test_se );
  input [7:0] DataIn;
  output [7:0] DataOut;
  input Write, Clk, Reset, SyncReset, eth_top_test_point_11887_in, test_si,
         test_se;
  wire   n21, n22, n23, n24, n25, n26, n27, n28, n1, n2, n3, n4;

  SDFFARX1 \DataOut_reg[7]  ( .D(n21), .SI(DataOut[6]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[7]) );
  SDFFASX1 \DataOut_reg[6]  ( .D(n22), .SI(DataOut[5]), .SE(test_se), .CLK(Clk), .SETB(n4), .Q(DataOut[6]) );
  SDFFARX1 \DataOut_reg[5]  ( .D(n23), .SI(DataOut[4]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[5]) );
  SDFFARX1 \DataOut_reg[4]  ( .D(n24), .SI(DataOut[3]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[4]) );
  SDFFARX1 \DataOut_reg[3]  ( .D(n25), .SI(DataOut[2]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[3]) );
  SDFFARX1 \DataOut_reg[2]  ( .D(n26), .SI(DataOut[1]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[2]) );
  SDFFARX1 \DataOut_reg[1]  ( .D(n27), .SI(DataOut[0]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[1]) );
  SDFFARX1 \DataOut_reg[0]  ( .D(n28), .SI(test_si), .SE(test_se), .CLK(Clk), 
        .RSTB(n4), .Q(DataOut[0]) );
  INVX0 U3 ( .INP(eth_top_test_point_11887_in), .ZN(n4) );
  AO22X1 U4 ( .IN1(DataIn[0]), .IN2(n1), .IN3(n2), .IN4(DataOut[0]), .Q(n28)
         );
  AO22X1 U5 ( .IN1(DataIn[1]), .IN2(n1), .IN3(n2), .IN4(DataOut[1]), .Q(n27)
         );
  AO22X1 U6 ( .IN1(DataIn[2]), .IN2(n1), .IN3(n2), .IN4(DataOut[2]), .Q(n26)
         );
  AO22X1 U7 ( .IN1(DataIn[3]), .IN2(n1), .IN3(n2), .IN4(DataOut[3]), .Q(n25)
         );
  AO22X1 U8 ( .IN1(DataIn[4]), .IN2(n1), .IN3(n2), .IN4(DataOut[4]), .Q(n24)
         );
  AO22X1 U9 ( .IN1(DataIn[5]), .IN2(n1), .IN3(n2), .IN4(DataOut[5]), .Q(n23)
         );
  AO221X1 U10 ( .IN1(n2), .IN2(DataOut[6]), .IN3(DataIn[6]), .IN4(n1), .IN5(
        SyncReset), .Q(n22) );
  AO22X1 U11 ( .IN1(DataIn[7]), .IN2(n1), .IN3(n2), .IN4(DataOut[7]), .Q(n21)
         );
  NOR2X0 U12 ( .IN1(n1), .IN2(SyncReset), .QN(n2) );
  NOR2X0 U13 ( .IN1(n3), .IN2(SyncReset), .QN(n1) );
  INVX0 U14 ( .INP(Write), .ZN(n3) );
endmodule


module eth_register_3_0_test_1 ( DataIn, DataOut, Write, Clk, Reset, SyncReset, 
        eth_top_test_point_11887_in, test_si, test_se );
  input [2:0] DataIn;
  output [2:0] DataOut;
  input Write, Clk, Reset, SyncReset, eth_top_test_point_11887_in, test_si,
         test_se;
  wire   n7, n8, n9, n1, n2, n3, n4;

  SDFFARX1 \DataOut_reg[2]  ( .D(n9), .SI(DataOut[1]), .SE(test_se), .CLK(Clk), 
        .RSTB(n4), .Q(DataOut[2]) );
  SDFFARX1 \DataOut_reg[1]  ( .D(n8), .SI(DataOut[0]), .SE(test_se), .CLK(Clk), 
        .RSTB(n4), .Q(DataOut[1]) );
  SDFFARX1 \DataOut_reg[0]  ( .D(n7), .SI(test_si), .SE(test_se), .CLK(Clk), 
        .RSTB(n4), .Q(DataOut[0]) );
  INVX0 U2 ( .INP(eth_top_test_point_11887_in), .ZN(n4) );
  AO22X1 U3 ( .IN1(DataIn[2]), .IN2(n1), .IN3(n2), .IN4(DataOut[2]), .Q(n9) );
  AO22X1 U4 ( .IN1(DataIn[1]), .IN2(n1), .IN3(n2), .IN4(DataOut[1]), .Q(n8) );
  AO22X1 U5 ( .IN1(DataIn[0]), .IN2(n1), .IN3(n2), .IN4(DataOut[0]), .Q(n7) );
  NOR2X0 U6 ( .IN1(SyncReset), .IN2(Write), .QN(n2) );
  NOR2X0 U7 ( .IN1(n3), .IN2(SyncReset), .QN(n1) );
  INVX0 U8 ( .INP(Write), .ZN(n3) );
endmodule


module eth_register_8_64_test_1 ( DataIn, DataOut, Write, Clk, Reset, 
        SyncReset, eth_top_test_point_11887_in, test_si, test_se );
  input [7:0] DataIn;
  output [7:0] DataOut;
  input Write, Clk, Reset, SyncReset, eth_top_test_point_11887_in, test_si,
         test_se;
  wire   n13, n14, n15, n16, n17, n18, n19, n20, n1, n2, n3, n4;

  SDFFARX1 \DataOut_reg[7]  ( .D(n20), .SI(DataOut[6]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[7]) );
  SDFFASX1 \DataOut_reg[6]  ( .D(n19), .SI(DataOut[5]), .SE(test_se), .CLK(Clk), .SETB(n4), .Q(DataOut[6]) );
  SDFFASX1 \DataOut_reg[5]  ( .D(n18), .SI(DataOut[4]), .SE(test_se), .CLK(Clk), .SETB(n4), .Q(DataOut[5]) );
  SDFFARX1 \DataOut_reg[4]  ( .D(n17), .SI(DataOut[3]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[4]) );
  SDFFARX1 \DataOut_reg[3]  ( .D(n16), .SI(DataOut[2]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[3]) );
  SDFFASX1 \DataOut_reg[2]  ( .D(n15), .SI(DataOut[1]), .SE(test_se), .CLK(Clk), .SETB(n4), .Q(DataOut[2]) );
  SDFFARX1 \DataOut_reg[1]  ( .D(n14), .SI(DataOut[0]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[1]) );
  SDFFARX1 \DataOut_reg[0]  ( .D(n13), .SI(test_si), .SE(test_se), .CLK(Clk), 
        .RSTB(n4), .Q(DataOut[0]) );
  INVX0 U3 ( .INP(eth_top_test_point_11887_in), .ZN(n4) );
  AO22X1 U4 ( .IN1(DataIn[7]), .IN2(n1), .IN3(n2), .IN4(DataOut[7]), .Q(n20)
         );
  AO221X1 U5 ( .IN1(n2), .IN2(DataOut[6]), .IN3(DataIn[6]), .IN4(n1), .IN5(
        SyncReset), .Q(n19) );
  AO221X1 U6 ( .IN1(n2), .IN2(DataOut[5]), .IN3(DataIn[5]), .IN4(n1), .IN5(
        SyncReset), .Q(n18) );
  AO22X1 U7 ( .IN1(DataIn[4]), .IN2(n1), .IN3(n2), .IN4(DataOut[4]), .Q(n17)
         );
  AO22X1 U8 ( .IN1(DataIn[3]), .IN2(n1), .IN3(n2), .IN4(DataOut[3]), .Q(n16)
         );
  AO221X1 U9 ( .IN1(n2), .IN2(DataOut[2]), .IN3(DataIn[2]), .IN4(n1), .IN5(
        SyncReset), .Q(n15) );
  AO22X1 U10 ( .IN1(DataIn[1]), .IN2(n1), .IN3(n2), .IN4(DataOut[1]), .Q(n14)
         );
  AO22X1 U11 ( .IN1(DataIn[0]), .IN2(n1), .IN3(n2), .IN4(DataOut[0]), .Q(n13)
         );
  NOR2X0 U12 ( .IN1(n1), .IN2(SyncReset), .QN(n2) );
  NOR2X0 U13 ( .IN1(n3), .IN2(SyncReset), .QN(n1) );
  INVX0 U14 ( .INP(Write), .ZN(n3) );
endmodule


module eth_register_1_0_test_2 ( DataIn, DataOut, Write, Clk, Reset, SyncReset, 
        eth_top_test_point_11887_in, test_si, test_se );
  input [0:0] DataIn;
  output [0:0] DataOut;
  input Write, Clk, Reset, SyncReset, eth_top_test_point_11887_in, test_si,
         test_se;
  wire   n6, n1, n2, n3;

  SDFFARX1 \DataOut_reg[0]  ( .D(n6), .SI(test_si), .SE(test_se), .CLK(Clk), 
        .RSTB(n3), .Q(DataOut[0]) );
  INVX0 U2 ( .INP(eth_top_test_point_11887_in), .ZN(n3) );
  NOR2X0 U3 ( .IN1(SyncReset), .IN2(n1), .QN(n6) );
  INVX0 U4 ( .INP(n2), .ZN(n1) );
  MUX21X1 U5 ( .IN1(DataOut[0]), .IN2(DataIn[0]), .S(Write), .Q(n2) );
endmodule


module eth_register_WIDTH1_RESET_VALUE0_test_0 ( DataIn, DataOut, Write, Clk, 
        Reset, SyncReset, eth_top_test_point_11887_in, test_si, test_se );
  input [0:0] DataIn;
  output [0:0] DataOut;
  input Write, Clk, Reset, SyncReset, eth_top_test_point_11887_in, test_si,
         test_se;
  wire   n5, n1, n2, n3;

  SDFFARX1 \DataOut_reg[0]  ( .D(n5), .SI(test_si), .SE(test_se), .CLK(Clk), 
        .RSTB(n3), .Q(DataOut[0]) );
  INVX0 U2 ( .INP(eth_top_test_point_11887_in), .ZN(n3) );
  NOR2X0 U3 ( .IN1(SyncReset), .IN2(n1), .QN(n5) );
  INVX0 U4 ( .INP(n2), .ZN(n1) );
  MUX21X1 U5 ( .IN1(DataOut[0]), .IN2(DataIn[0]), .S(Write), .Q(n2) );
endmodule


module eth_register_WIDTH1_RESET_VALUE0_test_2 ( DataIn, DataOut, Write, Clk, 
        Reset, SyncReset, eth_top_test_point_11887_in, test_si, test_se );
  input [0:0] DataIn;
  output [0:0] DataOut;
  input Write, Clk, Reset, SyncReset, eth_top_test_point_11887_in, test_si,
         test_se;
  wire   n6, n1, n2, n3;

  SDFFARX1 \DataOut_reg[0]  ( .D(n6), .SI(test_si), .SE(test_se), .CLK(Clk), 
        .RSTB(n3), .Q(DataOut[0]) );
  INVX0 U2 ( .INP(eth_top_test_point_11887_in), .ZN(n3) );
  NOR2X0 U3 ( .IN1(SyncReset), .IN2(n1), .QN(n6) );
  INVX0 U4 ( .INP(n2), .ZN(n1) );
  MUX21X1 U5 ( .IN1(DataOut[0]), .IN2(DataIn[0]), .S(Write), .Q(n2) );
endmodule


module eth_register_WIDTH1_RESET_VALUE0_test_1 ( DataIn, DataOut, Write, Clk, 
        Reset, SyncReset, eth_top_test_point_11887_in, test_si, test_se );
  input [0:0] DataIn;
  output [0:0] DataOut;
  input Write, Clk, Reset, SyncReset, eth_top_test_point_11887_in, test_si,
         test_se;
  wire   n6, n1, n2, n3;

  SDFFARX1 \DataOut_reg[0]  ( .D(n6), .SI(test_si), .SE(test_se), .CLK(Clk), 
        .RSTB(n3), .Q(DataOut[0]) );
  INVX0 U2 ( .INP(eth_top_test_point_11887_in), .ZN(n3) );
  NOR2X0 U3 ( .IN1(SyncReset), .IN2(n1), .QN(n6) );
  INVX0 U4 ( .INP(n2), .ZN(n1) );
  MUX21X1 U5 ( .IN1(DataOut[0]), .IN2(DataIn[0]), .S(Write), .Q(n2) );
endmodule


module eth_register_5_00_test_0 ( DataIn, DataOut, Write, Clk, Reset, 
        SyncReset, eth_top_test_point_11887_in, test_si, test_se );
  input [4:0] DataIn;
  output [4:0] DataOut;
  input Write, Clk, Reset, SyncReset, eth_top_test_point_11887_in, test_si,
         test_se;
  wire   n10, n11, n12, n13, n14, n1, n2, n3, n4;

  SDFFARX1 \DataOut_reg[4]  ( .D(n14), .SI(DataOut[3]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[4]) );
  SDFFARX1 \DataOut_reg[3]  ( .D(n13), .SI(DataOut[2]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[3]) );
  SDFFARX1 \DataOut_reg[2]  ( .D(n12), .SI(DataOut[1]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[2]) );
  SDFFARX1 \DataOut_reg[1]  ( .D(n11), .SI(DataOut[0]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[1]) );
  SDFFARX1 \DataOut_reg[0]  ( .D(n10), .SI(test_si), .SE(test_se), .CLK(Clk), 
        .RSTB(n4), .Q(DataOut[0]) );
  INVX0 U2 ( .INP(eth_top_test_point_11887_in), .ZN(n4) );
  AO22X1 U3 ( .IN1(DataIn[4]), .IN2(n1), .IN3(n2), .IN4(DataOut[4]), .Q(n14)
         );
  AO22X1 U4 ( .IN1(DataIn[3]), .IN2(n1), .IN3(n2), .IN4(DataOut[3]), .Q(n13)
         );
  AO22X1 U5 ( .IN1(DataIn[2]), .IN2(n1), .IN3(n2), .IN4(DataOut[2]), .Q(n12)
         );
  AO22X1 U6 ( .IN1(DataIn[1]), .IN2(n1), .IN3(n2), .IN4(DataOut[1]), .Q(n11)
         );
  AO22X1 U7 ( .IN1(DataIn[0]), .IN2(n1), .IN3(n2), .IN4(DataOut[0]), .Q(n10)
         );
  NOR2X0 U8 ( .IN1(n1), .IN2(SyncReset), .QN(n2) );
  NOR2X0 U9 ( .IN1(n3), .IN2(SyncReset), .QN(n1) );
  INVX0 U10 ( .INP(Write), .ZN(n3) );
endmodule


module eth_register_5_00_test_1 ( DataIn, DataOut, Write, Clk, Reset, 
        SyncReset, eth_top_test_point_11887_in, test_si, test_se );
  input [4:0] DataIn;
  output [4:0] DataOut;
  input Write, Clk, Reset, SyncReset, eth_top_test_point_11887_in, test_si,
         test_se;
  wire   n15, n16, n17, n18, n19, n1, n2, n3, n4;

  SDFFARX1 \DataOut_reg[4]  ( .D(n15), .SI(DataOut[3]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[4]) );
  SDFFARX1 \DataOut_reg[3]  ( .D(n16), .SI(DataOut[2]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[3]) );
  SDFFARX1 \DataOut_reg[2]  ( .D(n17), .SI(DataOut[1]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[2]) );
  SDFFARX1 \DataOut_reg[1]  ( .D(n18), .SI(DataOut[0]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[1]) );
  SDFFARX1 \DataOut_reg[0]  ( .D(n19), .SI(test_si), .SE(test_se), .CLK(Clk), 
        .RSTB(n4), .Q(DataOut[0]) );
  INVX0 U2 ( .INP(eth_top_test_point_11887_in), .ZN(n4) );
  AO22X1 U3 ( .IN1(DataIn[0]), .IN2(n1), .IN3(n2), .IN4(DataOut[0]), .Q(n19)
         );
  AO22X1 U4 ( .IN1(DataIn[1]), .IN2(n1), .IN3(n2), .IN4(DataOut[1]), .Q(n18)
         );
  AO22X1 U5 ( .IN1(DataIn[2]), .IN2(n1), .IN3(n2), .IN4(DataOut[2]), .Q(n17)
         );
  AO22X1 U6 ( .IN1(DataIn[3]), .IN2(n1), .IN3(n2), .IN4(DataOut[3]), .Q(n16)
         );
  AO22X1 U7 ( .IN1(DataIn[4]), .IN2(n1), .IN3(n2), .IN4(DataOut[4]), .Q(n15)
         );
  NOR2X0 U8 ( .IN1(n1), .IN2(SyncReset), .QN(n2) );
  NOR2X0 U9 ( .IN1(n3), .IN2(SyncReset), .QN(n1) );
  INVX0 U10 ( .INP(Write), .ZN(n3) );
endmodule


module eth_register_8_00_test_18 ( DataIn, DataOut, Write, Clk, Reset, 
        SyncReset, eth_top_test_point_11887_in, test_si, test_se );
  input [7:0] DataIn;
  output [7:0] DataOut;
  input Write, Clk, Reset, SyncReset, eth_top_test_point_11887_in, test_si,
         test_se;
  wire   n21, n22, n23, n24, n25, n26, n27, n28, n1, n2, n3, n4;

  SDFFARX1 \DataOut_reg[7]  ( .D(n21), .SI(DataOut[6]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[7]) );
  SDFFARX1 \DataOut_reg[6]  ( .D(n22), .SI(DataOut[5]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[6]) );
  SDFFARX1 \DataOut_reg[5]  ( .D(n23), .SI(DataOut[4]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[5]) );
  SDFFARX1 \DataOut_reg[4]  ( .D(n24), .SI(DataOut[3]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[4]) );
  SDFFARX1 \DataOut_reg[3]  ( .D(n25), .SI(DataOut[2]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[3]) );
  SDFFARX1 \DataOut_reg[2]  ( .D(n26), .SI(DataOut[1]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[2]) );
  SDFFARX1 \DataOut_reg[1]  ( .D(n27), .SI(DataOut[0]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[1]) );
  SDFFARX1 \DataOut_reg[0]  ( .D(n28), .SI(test_si), .SE(test_se), .CLK(Clk), 
        .RSTB(n4), .Q(DataOut[0]) );
  INVX0 U2 ( .INP(eth_top_test_point_11887_in), .ZN(n4) );
  AO22X1 U3 ( .IN1(DataIn[0]), .IN2(n1), .IN3(n2), .IN4(DataOut[0]), .Q(n28)
         );
  AO22X1 U4 ( .IN1(DataIn[1]), .IN2(n1), .IN3(n2), .IN4(DataOut[1]), .Q(n27)
         );
  AO22X1 U5 ( .IN1(DataIn[2]), .IN2(n1), .IN3(n2), .IN4(DataOut[2]), .Q(n26)
         );
  AO22X1 U6 ( .IN1(DataIn[3]), .IN2(n1), .IN3(n2), .IN4(DataOut[3]), .Q(n25)
         );
  AO22X1 U7 ( .IN1(DataIn[4]), .IN2(n1), .IN3(n2), .IN4(DataOut[4]), .Q(n24)
         );
  AO22X1 U8 ( .IN1(DataIn[5]), .IN2(n1), .IN3(n2), .IN4(DataOut[5]), .Q(n23)
         );
  AO22X1 U9 ( .IN1(DataIn[6]), .IN2(n1), .IN3(n2), .IN4(DataOut[6]), .Q(n22)
         );
  AO22X1 U10 ( .IN1(DataIn[7]), .IN2(n1), .IN3(n2), .IN4(DataOut[7]), .Q(n21)
         );
  NOR2X0 U11 ( .IN1(n1), .IN2(SyncReset), .QN(n2) );
  NOR2X0 U12 ( .IN1(n3), .IN2(SyncReset), .QN(n1) );
  INVX0 U13 ( .INP(Write), .ZN(n3) );
endmodule


module eth_register_8_00_test_17 ( DataIn, DataOut, Write, Clk, Reset, 
        SyncReset, eth_top_test_point_11887_in, test_si, test_se );
  input [7:0] DataIn;
  output [7:0] DataOut;
  input Write, Clk, Reset, SyncReset, eth_top_test_point_11887_in, test_si,
         test_se;
  wire   n21, n22, n23, n24, n25, n26, n27, n28, n1, n2, n3, n4;

  SDFFARX1 \DataOut_reg[7]  ( .D(n21), .SI(DataOut[6]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[7]) );
  SDFFARX1 \DataOut_reg[6]  ( .D(n22), .SI(DataOut[5]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[6]) );
  SDFFARX1 \DataOut_reg[5]  ( .D(n23), .SI(DataOut[4]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[5]) );
  SDFFARX1 \DataOut_reg[4]  ( .D(n24), .SI(DataOut[3]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[4]) );
  SDFFARX1 \DataOut_reg[3]  ( .D(n25), .SI(DataOut[2]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[3]) );
  SDFFARX1 \DataOut_reg[2]  ( .D(n26), .SI(DataOut[1]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[2]) );
  SDFFARX1 \DataOut_reg[1]  ( .D(n27), .SI(DataOut[0]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[1]) );
  SDFFARX1 \DataOut_reg[0]  ( .D(n28), .SI(test_si), .SE(test_se), .CLK(Clk), 
        .RSTB(n4), .Q(DataOut[0]) );
  INVX0 U2 ( .INP(eth_top_test_point_11887_in), .ZN(n4) );
  AO22X1 U3 ( .IN1(DataIn[0]), .IN2(n1), .IN3(n2), .IN4(DataOut[0]), .Q(n28)
         );
  AO22X1 U4 ( .IN1(DataIn[1]), .IN2(n1), .IN3(n2), .IN4(DataOut[1]), .Q(n27)
         );
  AO22X1 U5 ( .IN1(DataIn[2]), .IN2(n1), .IN3(n2), .IN4(DataOut[2]), .Q(n26)
         );
  AO22X1 U6 ( .IN1(DataIn[3]), .IN2(n1), .IN3(n2), .IN4(DataOut[3]), .Q(n25)
         );
  AO22X1 U7 ( .IN1(DataIn[4]), .IN2(n1), .IN3(n2), .IN4(DataOut[4]), .Q(n24)
         );
  AO22X1 U8 ( .IN1(DataIn[5]), .IN2(n1), .IN3(n2), .IN4(DataOut[5]), .Q(n23)
         );
  AO22X1 U9 ( .IN1(DataIn[6]), .IN2(n1), .IN3(n2), .IN4(DataOut[6]), .Q(n22)
         );
  AO22X1 U10 ( .IN1(DataIn[7]), .IN2(n1), .IN3(n2), .IN4(DataOut[7]), .Q(n21)
         );
  NOR2X0 U11 ( .IN1(n1), .IN2(SyncReset), .QN(n2) );
  NOR2X0 U12 ( .IN1(n3), .IN2(SyncReset), .QN(n1) );
  INVX0 U13 ( .INP(Write), .ZN(n3) );
endmodule


module eth_register_16_0000_test_1 ( DataIn, DataOut, Write, Clk, Reset, 
        SyncReset, eth_top_test_point_11887_in, test_si, test_se );
  input [15:0] DataIn;
  output [15:0] DataOut;
  input Write, Clk, Reset, SyncReset, eth_top_test_point_11887_in, test_si,
         test_se;
  wire   n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n1, n2, n3, n4;

  SDFFARX1 \DataOut_reg[15]  ( .D(n36), .SI(DataOut[14]), .SE(test_se), .CLK(
        Clk), .RSTB(n4), .Q(DataOut[15]) );
  SDFFARX1 \DataOut_reg[14]  ( .D(n35), .SI(DataOut[13]), .SE(test_se), .CLK(
        Clk), .RSTB(n4), .Q(DataOut[14]) );
  SDFFARX1 \DataOut_reg[13]  ( .D(n34), .SI(DataOut[12]), .SE(test_se), .CLK(
        Clk), .RSTB(n4), .Q(DataOut[13]) );
  SDFFARX1 \DataOut_reg[12]  ( .D(n33), .SI(DataOut[11]), .SE(test_se), .CLK(
        Clk), .RSTB(n4), .Q(DataOut[12]) );
  SDFFARX1 \DataOut_reg[11]  ( .D(n32), .SI(DataOut[10]), .SE(test_se), .CLK(
        Clk), .RSTB(n4), .Q(DataOut[11]) );
  SDFFARX1 \DataOut_reg[10]  ( .D(n31), .SI(DataOut[9]), .SE(test_se), .CLK(
        Clk), .RSTB(n4), .Q(DataOut[10]) );
  SDFFARX1 \DataOut_reg[9]  ( .D(n30), .SI(DataOut[8]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[9]) );
  SDFFARX1 \DataOut_reg[8]  ( .D(n29), .SI(DataOut[7]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[8]) );
  SDFFARX1 \DataOut_reg[7]  ( .D(n28), .SI(DataOut[6]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[7]) );
  SDFFARX1 \DataOut_reg[6]  ( .D(n27), .SI(DataOut[5]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[6]) );
  SDFFARX1 \DataOut_reg[5]  ( .D(n26), .SI(DataOut[4]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[5]) );
  SDFFARX1 \DataOut_reg[4]  ( .D(n25), .SI(DataOut[3]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[4]) );
  SDFFARX1 \DataOut_reg[3]  ( .D(n24), .SI(DataOut[2]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[3]) );
  SDFFARX1 \DataOut_reg[2]  ( .D(n23), .SI(DataOut[1]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[2]) );
  SDFFARX1 \DataOut_reg[1]  ( .D(n22), .SI(DataOut[0]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[1]) );
  SDFFARX1 \DataOut_reg[0]  ( .D(n21), .SI(test_si), .SE(test_se), .CLK(Clk), 
        .RSTB(n4), .Q(DataOut[0]) );
  INVX0 U2 ( .INP(eth_top_test_point_11887_in), .ZN(n4) );
  AO22X1 U3 ( .IN1(DataIn[15]), .IN2(n1), .IN3(n2), .IN4(DataOut[15]), .Q(n36)
         );
  AO22X1 U4 ( .IN1(DataIn[14]), .IN2(n1), .IN3(n2), .IN4(DataOut[14]), .Q(n35)
         );
  AO22X1 U5 ( .IN1(DataIn[13]), .IN2(n1), .IN3(n2), .IN4(DataOut[13]), .Q(n34)
         );
  AO22X1 U6 ( .IN1(DataIn[12]), .IN2(n1), .IN3(n2), .IN4(DataOut[12]), .Q(n33)
         );
  AO22X1 U7 ( .IN1(DataIn[11]), .IN2(n1), .IN3(n2), .IN4(DataOut[11]), .Q(n32)
         );
  AO22X1 U8 ( .IN1(DataIn[10]), .IN2(n1), .IN3(n2), .IN4(DataOut[10]), .Q(n31)
         );
  AO22X1 U9 ( .IN1(DataIn[9]), .IN2(n1), .IN3(n2), .IN4(DataOut[9]), .Q(n30)
         );
  AO22X1 U10 ( .IN1(DataIn[8]), .IN2(n1), .IN3(n2), .IN4(DataOut[8]), .Q(n29)
         );
  AO22X1 U11 ( .IN1(DataIn[7]), .IN2(n1), .IN3(n2), .IN4(DataOut[7]), .Q(n28)
         );
  AO22X1 U12 ( .IN1(DataIn[6]), .IN2(n1), .IN3(n2), .IN4(DataOut[6]), .Q(n27)
         );
  AO22X1 U13 ( .IN1(DataIn[5]), .IN2(n1), .IN3(n2), .IN4(DataOut[5]), .Q(n26)
         );
  AO22X1 U14 ( .IN1(DataIn[4]), .IN2(n1), .IN3(n2), .IN4(DataOut[4]), .Q(n25)
         );
  AO22X1 U15 ( .IN1(DataIn[3]), .IN2(n1), .IN3(n2), .IN4(DataOut[3]), .Q(n24)
         );
  AO22X1 U16 ( .IN1(DataIn[2]), .IN2(n1), .IN3(n2), .IN4(DataOut[2]), .Q(n23)
         );
  AO22X1 U17 ( .IN1(DataIn[1]), .IN2(n1), .IN3(n2), .IN4(DataOut[1]), .Q(n22)
         );
  AO22X1 U18 ( .IN1(DataIn[0]), .IN2(n1), .IN3(n2), .IN4(DataOut[0]), .Q(n21)
         );
  NOR2X0 U19 ( .IN1(n1), .IN2(SyncReset), .QN(n2) );
  NOR2X0 U20 ( .IN1(n3), .IN2(SyncReset), .QN(n1) );
  INVX0 U21 ( .INP(Write), .ZN(n3) );
endmodule


module eth_register_8_00_test_16 ( DataIn, DataOut, Write, Clk, Reset, 
        SyncReset, eth_top_test_point_11887_in, test_si, test_se );
  input [7:0] DataIn;
  output [7:0] DataOut;
  input Write, Clk, Reset, SyncReset, eth_top_test_point_11887_in, test_si,
         test_se;
  wire   n21, n22, n23, n24, n25, n26, n27, n28, n1, n2, n3, n4;

  SDFFARX1 \DataOut_reg[7]  ( .D(n21), .SI(DataOut[6]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[7]) );
  SDFFARX1 \DataOut_reg[6]  ( .D(n22), .SI(DataOut[5]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[6]) );
  SDFFARX1 \DataOut_reg[5]  ( .D(n23), .SI(DataOut[4]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[5]) );
  SDFFARX1 \DataOut_reg[4]  ( .D(n24), .SI(DataOut[3]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[4]) );
  SDFFARX1 \DataOut_reg[3]  ( .D(n25), .SI(DataOut[2]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[3]) );
  SDFFARX1 \DataOut_reg[2]  ( .D(n26), .SI(DataOut[1]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[2]) );
  SDFFARX1 \DataOut_reg[1]  ( .D(n27), .SI(DataOut[0]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[1]) );
  SDFFARX1 \DataOut_reg[0]  ( .D(n28), .SI(test_si), .SE(test_se), .CLK(Clk), 
        .RSTB(n4), .Q(DataOut[0]) );
  INVX0 U2 ( .INP(eth_top_test_point_11887_in), .ZN(n4) );
  AO22X1 U3 ( .IN1(DataIn[0]), .IN2(n1), .IN3(n2), .IN4(DataOut[0]), .Q(n28)
         );
  AO22X1 U4 ( .IN1(DataIn[1]), .IN2(n1), .IN3(n2), .IN4(DataOut[1]), .Q(n27)
         );
  AO22X1 U5 ( .IN1(DataIn[2]), .IN2(n1), .IN3(n2), .IN4(DataOut[2]), .Q(n26)
         );
  AO22X1 U6 ( .IN1(DataIn[3]), .IN2(n1), .IN3(n2), .IN4(DataOut[3]), .Q(n25)
         );
  AO22X1 U7 ( .IN1(DataIn[4]), .IN2(n1), .IN3(n2), .IN4(DataOut[4]), .Q(n24)
         );
  AO22X1 U8 ( .IN1(DataIn[5]), .IN2(n1), .IN3(n2), .IN4(DataOut[5]), .Q(n23)
         );
  AO22X1 U9 ( .IN1(DataIn[6]), .IN2(n1), .IN3(n2), .IN4(DataOut[6]), .Q(n22)
         );
  AO22X1 U10 ( .IN1(DataIn[7]), .IN2(n1), .IN3(n2), .IN4(DataOut[7]), .Q(n21)
         );
  NOR2X0 U11 ( .IN1(n1), .IN2(SyncReset), .QN(n2) );
  NOR2X0 U12 ( .IN1(n3), .IN2(SyncReset), .QN(n1) );
  INVX0 U13 ( .INP(Write), .ZN(n3) );
endmodule


module eth_register_8_00_test_15 ( DataIn, DataOut, Write, Clk, Reset, 
        SyncReset, eth_top_test_point_11887_in, test_si, test_se );
  input [7:0] DataIn;
  output [7:0] DataOut;
  input Write, Clk, Reset, SyncReset, eth_top_test_point_11887_in, test_si,
         test_se;
  wire   n21, n22, n23, n24, n25, n26, n27, n28, n1, n2, n3, n4;

  SDFFARX1 \DataOut_reg[7]  ( .D(n21), .SI(DataOut[6]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[7]) );
  SDFFARX1 \DataOut_reg[6]  ( .D(n22), .SI(DataOut[5]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[6]) );
  SDFFARX1 \DataOut_reg[5]  ( .D(n23), .SI(DataOut[4]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[5]) );
  SDFFARX1 \DataOut_reg[4]  ( .D(n24), .SI(DataOut[3]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[4]) );
  SDFFARX1 \DataOut_reg[3]  ( .D(n25), .SI(DataOut[2]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[3]) );
  SDFFARX1 \DataOut_reg[2]  ( .D(n26), .SI(DataOut[1]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[2]) );
  SDFFARX1 \DataOut_reg[1]  ( .D(n27), .SI(DataOut[0]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[1]) );
  SDFFARX1 \DataOut_reg[0]  ( .D(n28), .SI(test_si), .SE(test_se), .CLK(Clk), 
        .RSTB(n4), .Q(DataOut[0]) );
  INVX0 U2 ( .INP(eth_top_test_point_11887_in), .ZN(n4) );
  AO22X1 U3 ( .IN1(DataIn[0]), .IN2(n1), .IN3(n2), .IN4(DataOut[0]), .Q(n28)
         );
  AO22X1 U4 ( .IN1(DataIn[1]), .IN2(n1), .IN3(n2), .IN4(DataOut[1]), .Q(n27)
         );
  AO22X1 U5 ( .IN1(DataIn[2]), .IN2(n1), .IN3(n2), .IN4(DataOut[2]), .Q(n26)
         );
  AO22X1 U6 ( .IN1(DataIn[3]), .IN2(n1), .IN3(n2), .IN4(DataOut[3]), .Q(n25)
         );
  AO22X1 U7 ( .IN1(DataIn[4]), .IN2(n1), .IN3(n2), .IN4(DataOut[4]), .Q(n24)
         );
  AO22X1 U8 ( .IN1(DataIn[5]), .IN2(n1), .IN3(n2), .IN4(DataOut[5]), .Q(n23)
         );
  AO22X1 U9 ( .IN1(DataIn[6]), .IN2(n1), .IN3(n2), .IN4(DataOut[6]), .Q(n22)
         );
  AO22X1 U10 ( .IN1(DataIn[7]), .IN2(n1), .IN3(n2), .IN4(DataOut[7]), .Q(n21)
         );
  NOR2X0 U11 ( .IN1(n1), .IN2(SyncReset), .QN(n2) );
  NOR2X0 U12 ( .IN1(n3), .IN2(SyncReset), .QN(n1) );
  INVX0 U13 ( .INP(Write), .ZN(n3) );
endmodule


module eth_register_8_00_test_14 ( DataIn, DataOut, Write, Clk, Reset, 
        SyncReset, eth_top_test_point_11887_in, test_si, test_se );
  input [7:0] DataIn;
  output [7:0] DataOut;
  input Write, Clk, Reset, SyncReset, eth_top_test_point_11887_in, test_si,
         test_se;
  wire   n21, n22, n23, n24, n25, n26, n27, n28, n1, n2, n3, n4;

  SDFFARX1 \DataOut_reg[7]  ( .D(n21), .SI(DataOut[6]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[7]) );
  SDFFARX1 \DataOut_reg[6]  ( .D(n22), .SI(DataOut[5]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[6]) );
  SDFFARX1 \DataOut_reg[5]  ( .D(n23), .SI(DataOut[4]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[5]) );
  SDFFARX1 \DataOut_reg[4]  ( .D(n24), .SI(DataOut[3]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[4]) );
  SDFFARX1 \DataOut_reg[3]  ( .D(n25), .SI(DataOut[2]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[3]) );
  SDFFARX1 \DataOut_reg[2]  ( .D(n26), .SI(DataOut[1]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[2]) );
  SDFFARX1 \DataOut_reg[1]  ( .D(n27), .SI(DataOut[0]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[1]) );
  SDFFARX1 \DataOut_reg[0]  ( .D(n28), .SI(test_si), .SE(test_se), .CLK(Clk), 
        .RSTB(n4), .Q(DataOut[0]) );
  INVX0 U2 ( .INP(eth_top_test_point_11887_in), .ZN(n4) );
  AO22X1 U3 ( .IN1(DataIn[0]), .IN2(n1), .IN3(n2), .IN4(DataOut[0]), .Q(n28)
         );
  AO22X1 U4 ( .IN1(DataIn[1]), .IN2(n1), .IN3(n2), .IN4(DataOut[1]), .Q(n27)
         );
  AO22X1 U5 ( .IN1(DataIn[2]), .IN2(n1), .IN3(n2), .IN4(DataOut[2]), .Q(n26)
         );
  AO22X1 U6 ( .IN1(DataIn[3]), .IN2(n1), .IN3(n2), .IN4(DataOut[3]), .Q(n25)
         );
  AO22X1 U7 ( .IN1(DataIn[4]), .IN2(n1), .IN3(n2), .IN4(DataOut[4]), .Q(n24)
         );
  AO22X1 U8 ( .IN1(DataIn[5]), .IN2(n1), .IN3(n2), .IN4(DataOut[5]), .Q(n23)
         );
  AO22X1 U9 ( .IN1(DataIn[6]), .IN2(n1), .IN3(n2), .IN4(DataOut[6]), .Q(n22)
         );
  AO22X1 U10 ( .IN1(DataIn[7]), .IN2(n1), .IN3(n2), .IN4(DataOut[7]), .Q(n21)
         );
  NOR2X0 U11 ( .IN1(n1), .IN2(SyncReset), .QN(n2) );
  NOR2X0 U12 ( .IN1(n3), .IN2(SyncReset), .QN(n1) );
  INVX0 U13 ( .INP(Write), .ZN(n3) );
endmodule


module eth_register_8_00_test_13 ( DataIn, DataOut, Write, Clk, Reset, 
        SyncReset, eth_top_test_point_11887_in, test_si, test_se );
  input [7:0] DataIn;
  output [7:0] DataOut;
  input Write, Clk, Reset, SyncReset, eth_top_test_point_11887_in, test_si,
         test_se;
  wire   n21, n22, n23, n24, n25, n26, n27, n28, n1, n2, n3, n4;

  SDFFARX1 \DataOut_reg[7]  ( .D(n21), .SI(DataOut[6]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[7]) );
  SDFFARX1 \DataOut_reg[6]  ( .D(n22), .SI(DataOut[5]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[6]) );
  SDFFARX1 \DataOut_reg[5]  ( .D(n23), .SI(DataOut[4]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[5]) );
  SDFFARX1 \DataOut_reg[4]  ( .D(n24), .SI(DataOut[3]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[4]) );
  SDFFARX1 \DataOut_reg[3]  ( .D(n25), .SI(DataOut[2]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[3]) );
  SDFFARX1 \DataOut_reg[2]  ( .D(n26), .SI(DataOut[1]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[2]) );
  SDFFARX1 \DataOut_reg[1]  ( .D(n27), .SI(DataOut[0]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[1]) );
  SDFFARX1 \DataOut_reg[0]  ( .D(n28), .SI(test_si), .SE(test_se), .CLK(Clk), 
        .RSTB(n4), .Q(DataOut[0]) );
  INVX0 U2 ( .INP(eth_top_test_point_11887_in), .ZN(n4) );
  AO22X1 U3 ( .IN1(DataIn[0]), .IN2(n1), .IN3(n2), .IN4(DataOut[0]), .Q(n28)
         );
  AO22X1 U4 ( .IN1(DataIn[1]), .IN2(n1), .IN3(n2), .IN4(DataOut[1]), .Q(n27)
         );
  AO22X1 U5 ( .IN1(DataIn[2]), .IN2(n1), .IN3(n2), .IN4(DataOut[2]), .Q(n26)
         );
  AO22X1 U6 ( .IN1(DataIn[3]), .IN2(n1), .IN3(n2), .IN4(DataOut[3]), .Q(n25)
         );
  AO22X1 U7 ( .IN1(DataIn[4]), .IN2(n1), .IN3(n2), .IN4(DataOut[4]), .Q(n24)
         );
  AO22X1 U8 ( .IN1(DataIn[5]), .IN2(n1), .IN3(n2), .IN4(DataOut[5]), .Q(n23)
         );
  AO22X1 U9 ( .IN1(DataIn[6]), .IN2(n1), .IN3(n2), .IN4(DataOut[6]), .Q(n22)
         );
  AO22X1 U10 ( .IN1(DataIn[7]), .IN2(n1), .IN3(n2), .IN4(DataOut[7]), .Q(n21)
         );
  NOR2X0 U11 ( .IN1(n1), .IN2(SyncReset), .QN(n2) );
  NOR2X0 U12 ( .IN1(n3), .IN2(SyncReset), .QN(n1) );
  INVX0 U13 ( .INP(Write), .ZN(n3) );
endmodule


module eth_register_8_00_test_12 ( DataIn, DataOut, Write, Clk, Reset, 
        SyncReset, eth_top_test_point_11887_in, test_si, test_se );
  input [7:0] DataIn;
  output [7:0] DataOut;
  input Write, Clk, Reset, SyncReset, eth_top_test_point_11887_in, test_si,
         test_se;
  wire   n21, n22, n23, n24, n25, n26, n27, n28, n1, n2, n3, n4;

  SDFFARX1 \DataOut_reg[7]  ( .D(n21), .SI(DataOut[6]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[7]) );
  SDFFARX1 \DataOut_reg[6]  ( .D(n22), .SI(DataOut[5]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[6]) );
  SDFFARX1 \DataOut_reg[5]  ( .D(n23), .SI(DataOut[4]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[5]) );
  SDFFARX1 \DataOut_reg[4]  ( .D(n24), .SI(DataOut[3]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[4]) );
  SDFFARX1 \DataOut_reg[3]  ( .D(n25), .SI(DataOut[2]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[3]) );
  SDFFARX1 \DataOut_reg[2]  ( .D(n26), .SI(DataOut[1]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[2]) );
  SDFFARX1 \DataOut_reg[1]  ( .D(n27), .SI(DataOut[0]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[1]) );
  SDFFARX1 \DataOut_reg[0]  ( .D(n28), .SI(test_si), .SE(test_se), .CLK(Clk), 
        .RSTB(n4), .Q(DataOut[0]) );
  INVX0 U2 ( .INP(eth_top_test_point_11887_in), .ZN(n4) );
  AO22X1 U3 ( .IN1(DataIn[0]), .IN2(n1), .IN3(n2), .IN4(DataOut[0]), .Q(n28)
         );
  AO22X1 U4 ( .IN1(DataIn[1]), .IN2(n1), .IN3(n2), .IN4(DataOut[1]), .Q(n27)
         );
  AO22X1 U5 ( .IN1(DataIn[2]), .IN2(n1), .IN3(n2), .IN4(DataOut[2]), .Q(n26)
         );
  AO22X1 U6 ( .IN1(DataIn[3]), .IN2(n1), .IN3(n2), .IN4(DataOut[3]), .Q(n25)
         );
  AO22X1 U7 ( .IN1(DataIn[4]), .IN2(n1), .IN3(n2), .IN4(DataOut[4]), .Q(n24)
         );
  AO22X1 U8 ( .IN1(DataIn[5]), .IN2(n1), .IN3(n2), .IN4(DataOut[5]), .Q(n23)
         );
  AO22X1 U9 ( .IN1(DataIn[6]), .IN2(n1), .IN3(n2), .IN4(DataOut[6]), .Q(n22)
         );
  AO22X1 U10 ( .IN1(DataIn[7]), .IN2(n1), .IN3(n2), .IN4(DataOut[7]), .Q(n21)
         );
  NOR2X0 U11 ( .IN1(n1), .IN2(SyncReset), .QN(n2) );
  NOR2X0 U12 ( .IN1(n3), .IN2(SyncReset), .QN(n1) );
  INVX0 U13 ( .INP(Write), .ZN(n3) );
endmodule


module eth_register_8_00_test_11 ( DataIn, DataOut, Write, Clk, Reset, 
        SyncReset, eth_top_test_point_11887_in, test_si, test_se );
  input [7:0] DataIn;
  output [7:0] DataOut;
  input Write, Clk, Reset, SyncReset, eth_top_test_point_11887_in, test_si,
         test_se;
  wire   n21, n22, n23, n24, n25, n26, n27, n28, n1, n2, n3, n4;

  SDFFARX1 \DataOut_reg[7]  ( .D(n21), .SI(DataOut[6]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[7]) );
  SDFFARX1 \DataOut_reg[6]  ( .D(n22), .SI(DataOut[5]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[6]) );
  SDFFARX1 \DataOut_reg[5]  ( .D(n23), .SI(DataOut[4]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[5]) );
  SDFFARX1 \DataOut_reg[4]  ( .D(n24), .SI(DataOut[3]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[4]) );
  SDFFARX1 \DataOut_reg[3]  ( .D(n25), .SI(DataOut[2]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[3]) );
  SDFFARX1 \DataOut_reg[2]  ( .D(n26), .SI(DataOut[1]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[2]) );
  SDFFARX1 \DataOut_reg[1]  ( .D(n27), .SI(DataOut[0]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[1]) );
  SDFFARX1 \DataOut_reg[0]  ( .D(n28), .SI(test_si), .SE(test_se), .CLK(Clk), 
        .RSTB(n4), .Q(DataOut[0]) );
  INVX0 U2 ( .INP(eth_top_test_point_11887_in), .ZN(n4) );
  AO22X1 U3 ( .IN1(DataIn[0]), .IN2(n1), .IN3(n2), .IN4(DataOut[0]), .Q(n28)
         );
  AO22X1 U4 ( .IN1(DataIn[1]), .IN2(n1), .IN3(n2), .IN4(DataOut[1]), .Q(n27)
         );
  AO22X1 U5 ( .IN1(DataIn[2]), .IN2(n1), .IN3(n2), .IN4(DataOut[2]), .Q(n26)
         );
  AO22X1 U6 ( .IN1(DataIn[3]), .IN2(n1), .IN3(n2), .IN4(DataOut[3]), .Q(n25)
         );
  AO22X1 U7 ( .IN1(DataIn[4]), .IN2(n1), .IN3(n2), .IN4(DataOut[4]), .Q(n24)
         );
  AO22X1 U8 ( .IN1(DataIn[5]), .IN2(n1), .IN3(n2), .IN4(DataOut[5]), .Q(n23)
         );
  AO22X1 U9 ( .IN1(DataIn[6]), .IN2(n1), .IN3(n2), .IN4(DataOut[6]), .Q(n22)
         );
  AO22X1 U10 ( .IN1(DataIn[7]), .IN2(n1), .IN3(n2), .IN4(DataOut[7]), .Q(n21)
         );
  NOR2X0 U11 ( .IN1(n1), .IN2(SyncReset), .QN(n2) );
  NOR2X0 U12 ( .IN1(n3), .IN2(SyncReset), .QN(n1) );
  INVX0 U13 ( .INP(Write), .ZN(n3) );
endmodule


module eth_register_8_00_test_10 ( DataIn, DataOut, Write, Clk, Reset, 
        SyncReset, eth_top_test_point_11887_in, test_si, test_se );
  input [7:0] DataIn;
  output [7:0] DataOut;
  input Write, Clk, Reset, SyncReset, eth_top_test_point_11887_in, test_si,
         test_se;
  wire   n21, n22, n23, n24, n25, n26, n27, n28, n1, n2, n3, n4;

  SDFFARX1 \DataOut_reg[7]  ( .D(n21), .SI(DataOut[6]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[7]) );
  SDFFARX1 \DataOut_reg[6]  ( .D(n22), .SI(DataOut[5]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[6]) );
  SDFFARX1 \DataOut_reg[5]  ( .D(n23), .SI(DataOut[4]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[5]) );
  SDFFARX1 \DataOut_reg[4]  ( .D(n24), .SI(DataOut[3]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[4]) );
  SDFFARX1 \DataOut_reg[3]  ( .D(n25), .SI(DataOut[2]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[3]) );
  SDFFARX1 \DataOut_reg[2]  ( .D(n26), .SI(DataOut[1]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[2]) );
  SDFFARX1 \DataOut_reg[1]  ( .D(n27), .SI(DataOut[0]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[1]) );
  SDFFARX1 \DataOut_reg[0]  ( .D(n28), .SI(test_si), .SE(test_se), .CLK(Clk), 
        .RSTB(n4), .Q(DataOut[0]) );
  INVX0 U2 ( .INP(eth_top_test_point_11887_in), .ZN(n4) );
  AO22X1 U3 ( .IN1(DataIn[0]), .IN2(n1), .IN3(n2), .IN4(DataOut[0]), .Q(n28)
         );
  AO22X1 U4 ( .IN1(DataIn[1]), .IN2(n1), .IN3(n2), .IN4(DataOut[1]), .Q(n27)
         );
  AO22X1 U5 ( .IN1(DataIn[2]), .IN2(n1), .IN3(n2), .IN4(DataOut[2]), .Q(n26)
         );
  AO22X1 U6 ( .IN1(DataIn[3]), .IN2(n1), .IN3(n2), .IN4(DataOut[3]), .Q(n25)
         );
  AO22X1 U7 ( .IN1(DataIn[4]), .IN2(n1), .IN3(n2), .IN4(DataOut[4]), .Q(n24)
         );
  AO22X1 U8 ( .IN1(DataIn[5]), .IN2(n1), .IN3(n2), .IN4(DataOut[5]), .Q(n23)
         );
  AO22X1 U9 ( .IN1(DataIn[6]), .IN2(n1), .IN3(n2), .IN4(DataOut[6]), .Q(n22)
         );
  AO22X1 U10 ( .IN1(DataIn[7]), .IN2(n1), .IN3(n2), .IN4(DataOut[7]), .Q(n21)
         );
  NOR2X0 U11 ( .IN1(n1), .IN2(SyncReset), .QN(n2) );
  NOR2X0 U12 ( .IN1(n3), .IN2(SyncReset), .QN(n1) );
  INVX0 U13 ( .INP(Write), .ZN(n3) );
endmodule


module eth_register_8_00_test_9 ( DataIn, DataOut, Write, Clk, Reset, 
        SyncReset, eth_top_test_point_11887_in, test_si, test_se );
  input [7:0] DataIn;
  output [7:0] DataOut;
  input Write, Clk, Reset, SyncReset, eth_top_test_point_11887_in, test_si,
         test_se;
  wire   n21, n22, n23, n24, n25, n26, n27, n28, n1, n2, n3, n4;

  SDFFARX1 \DataOut_reg[7]  ( .D(n21), .SI(DataOut[6]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[7]) );
  SDFFARX1 \DataOut_reg[6]  ( .D(n22), .SI(DataOut[5]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[6]) );
  SDFFARX1 \DataOut_reg[5]  ( .D(n23), .SI(DataOut[4]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[5]) );
  SDFFARX1 \DataOut_reg[4]  ( .D(n24), .SI(DataOut[3]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[4]) );
  SDFFARX1 \DataOut_reg[3]  ( .D(n25), .SI(DataOut[2]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[3]) );
  SDFFARX1 \DataOut_reg[2]  ( .D(n26), .SI(DataOut[1]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[2]) );
  SDFFARX1 \DataOut_reg[1]  ( .D(n27), .SI(DataOut[0]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[1]) );
  SDFFARX1 \DataOut_reg[0]  ( .D(n28), .SI(test_si), .SE(test_se), .CLK(Clk), 
        .RSTB(n4), .Q(DataOut[0]) );
  INVX0 U2 ( .INP(eth_top_test_point_11887_in), .ZN(n4) );
  AO22X1 U3 ( .IN1(DataIn[0]), .IN2(n1), .IN3(n2), .IN4(DataOut[0]), .Q(n28)
         );
  AO22X1 U4 ( .IN1(DataIn[1]), .IN2(n1), .IN3(n2), .IN4(DataOut[1]), .Q(n27)
         );
  AO22X1 U5 ( .IN1(DataIn[2]), .IN2(n1), .IN3(n2), .IN4(DataOut[2]), .Q(n26)
         );
  AO22X1 U6 ( .IN1(DataIn[3]), .IN2(n1), .IN3(n2), .IN4(DataOut[3]), .Q(n25)
         );
  AO22X1 U7 ( .IN1(DataIn[4]), .IN2(n1), .IN3(n2), .IN4(DataOut[4]), .Q(n24)
         );
  AO22X1 U8 ( .IN1(DataIn[5]), .IN2(n1), .IN3(n2), .IN4(DataOut[5]), .Q(n23)
         );
  AO22X1 U9 ( .IN1(DataIn[6]), .IN2(n1), .IN3(n2), .IN4(DataOut[6]), .Q(n22)
         );
  AO22X1 U10 ( .IN1(DataIn[7]), .IN2(n1), .IN3(n2), .IN4(DataOut[7]), .Q(n21)
         );
  NOR2X0 U11 ( .IN1(n1), .IN2(SyncReset), .QN(n2) );
  NOR2X0 U12 ( .IN1(n3), .IN2(SyncReset), .QN(n1) );
  INVX0 U13 ( .INP(Write), .ZN(n3) );
endmodule


module eth_register_8_00_test_8 ( DataIn, DataOut, Write, Clk, Reset, 
        SyncReset, eth_top_test_point_11887_in, test_si, test_se );
  input [7:0] DataIn;
  output [7:0] DataOut;
  input Write, Clk, Reset, SyncReset, eth_top_test_point_11887_in, test_si,
         test_se;
  wire   n21, n22, n23, n24, n25, n26, n27, n28, n1, n2, n3, n4;

  SDFFARX1 \DataOut_reg[7]  ( .D(n21), .SI(DataOut[6]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[7]) );
  SDFFARX1 \DataOut_reg[6]  ( .D(n22), .SI(DataOut[5]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[6]) );
  SDFFARX1 \DataOut_reg[5]  ( .D(n23), .SI(DataOut[4]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[5]) );
  SDFFARX1 \DataOut_reg[4]  ( .D(n24), .SI(DataOut[3]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[4]) );
  SDFFARX1 \DataOut_reg[3]  ( .D(n25), .SI(DataOut[2]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[3]) );
  SDFFARX1 \DataOut_reg[2]  ( .D(n26), .SI(DataOut[1]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[2]) );
  SDFFARX1 \DataOut_reg[1]  ( .D(n27), .SI(DataOut[0]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[1]) );
  SDFFARX1 \DataOut_reg[0]  ( .D(n28), .SI(test_si), .SE(test_se), .CLK(Clk), 
        .RSTB(n4), .Q(DataOut[0]) );
  INVX0 U2 ( .INP(eth_top_test_point_11887_in), .ZN(n4) );
  AO22X1 U3 ( .IN1(DataIn[0]), .IN2(n1), .IN3(n2), .IN4(DataOut[0]), .Q(n28)
         );
  AO22X1 U4 ( .IN1(DataIn[1]), .IN2(n1), .IN3(n2), .IN4(DataOut[1]), .Q(n27)
         );
  AO22X1 U5 ( .IN1(DataIn[2]), .IN2(n1), .IN3(n2), .IN4(DataOut[2]), .Q(n26)
         );
  AO22X1 U6 ( .IN1(DataIn[3]), .IN2(n1), .IN3(n2), .IN4(DataOut[3]), .Q(n25)
         );
  AO22X1 U7 ( .IN1(DataIn[4]), .IN2(n1), .IN3(n2), .IN4(DataOut[4]), .Q(n24)
         );
  AO22X1 U8 ( .IN1(DataIn[5]), .IN2(n1), .IN3(n2), .IN4(DataOut[5]), .Q(n23)
         );
  AO22X1 U9 ( .IN1(DataIn[6]), .IN2(n1), .IN3(n2), .IN4(DataOut[6]), .Q(n22)
         );
  AO22X1 U10 ( .IN1(DataIn[7]), .IN2(n1), .IN3(n2), .IN4(DataOut[7]), .Q(n21)
         );
  NOR2X0 U11 ( .IN1(n1), .IN2(SyncReset), .QN(n2) );
  NOR2X0 U12 ( .IN1(n3), .IN2(SyncReset), .QN(n1) );
  INVX0 U13 ( .INP(Write), .ZN(n3) );
endmodule


module eth_register_8_00_test_7 ( DataIn, DataOut, Write, Clk, Reset, 
        SyncReset, eth_top_test_point_11887_in, test_si, test_se );
  input [7:0] DataIn;
  output [7:0] DataOut;
  input Write, Clk, Reset, SyncReset, eth_top_test_point_11887_in, test_si,
         test_se;
  wire   n21, n22, n23, n24, n25, n26, n27, n28, n1, n2, n3, n4;

  SDFFARX1 \DataOut_reg[7]  ( .D(n21), .SI(DataOut[6]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[7]) );
  SDFFARX1 \DataOut_reg[6]  ( .D(n22), .SI(DataOut[5]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[6]) );
  SDFFARX1 \DataOut_reg[5]  ( .D(n23), .SI(DataOut[4]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[5]) );
  SDFFARX1 \DataOut_reg[4]  ( .D(n24), .SI(DataOut[3]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[4]) );
  SDFFARX1 \DataOut_reg[3]  ( .D(n25), .SI(DataOut[2]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[3]) );
  SDFFARX1 \DataOut_reg[2]  ( .D(n26), .SI(DataOut[1]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[2]) );
  SDFFARX1 \DataOut_reg[1]  ( .D(n27), .SI(DataOut[0]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[1]) );
  SDFFARX1 \DataOut_reg[0]  ( .D(n28), .SI(test_si), .SE(test_se), .CLK(Clk), 
        .RSTB(n4), .Q(DataOut[0]) );
  INVX0 U2 ( .INP(eth_top_test_point_11887_in), .ZN(n4) );
  AO22X1 U3 ( .IN1(DataIn[0]), .IN2(n1), .IN3(n2), .IN4(DataOut[0]), .Q(n28)
         );
  AO22X1 U4 ( .IN1(DataIn[1]), .IN2(n1), .IN3(n2), .IN4(DataOut[1]), .Q(n27)
         );
  AO22X1 U5 ( .IN1(DataIn[2]), .IN2(n1), .IN3(n2), .IN4(DataOut[2]), .Q(n26)
         );
  AO22X1 U6 ( .IN1(DataIn[3]), .IN2(n1), .IN3(n2), .IN4(DataOut[3]), .Q(n25)
         );
  AO22X1 U7 ( .IN1(DataIn[4]), .IN2(n1), .IN3(n2), .IN4(DataOut[4]), .Q(n24)
         );
  AO22X1 U8 ( .IN1(DataIn[5]), .IN2(n1), .IN3(n2), .IN4(DataOut[5]), .Q(n23)
         );
  AO22X1 U9 ( .IN1(DataIn[6]), .IN2(n1), .IN3(n2), .IN4(DataOut[6]), .Q(n22)
         );
  AO22X1 U10 ( .IN1(DataIn[7]), .IN2(n1), .IN3(n2), .IN4(DataOut[7]), .Q(n21)
         );
  NOR2X0 U11 ( .IN1(n1), .IN2(SyncReset), .QN(n2) );
  NOR2X0 U12 ( .IN1(n3), .IN2(SyncReset), .QN(n1) );
  INVX0 U13 ( .INP(Write), .ZN(n3) );
endmodule


module eth_register_8_00_test_6 ( DataIn, DataOut, Write, Clk, Reset, 
        SyncReset, eth_top_test_point_11887_in, test_si, test_se );
  input [7:0] DataIn;
  output [7:0] DataOut;
  input Write, Clk, Reset, SyncReset, eth_top_test_point_11887_in, test_si,
         test_se;
  wire   n21, n22, n23, n24, n25, n26, n27, n28, n1, n2, n3, n4;

  SDFFARX1 \DataOut_reg[7]  ( .D(n21), .SI(DataOut[6]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[7]) );
  SDFFARX1 \DataOut_reg[6]  ( .D(n22), .SI(DataOut[5]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[6]) );
  SDFFARX1 \DataOut_reg[5]  ( .D(n23), .SI(DataOut[4]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[5]) );
  SDFFARX1 \DataOut_reg[4]  ( .D(n24), .SI(DataOut[3]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[4]) );
  SDFFARX1 \DataOut_reg[3]  ( .D(n25), .SI(DataOut[2]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[3]) );
  SDFFARX1 \DataOut_reg[2]  ( .D(n26), .SI(DataOut[1]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[2]) );
  SDFFARX1 \DataOut_reg[1]  ( .D(n27), .SI(DataOut[0]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[1]) );
  SDFFARX1 \DataOut_reg[0]  ( .D(n28), .SI(test_si), .SE(test_se), .CLK(Clk), 
        .RSTB(n4), .Q(DataOut[0]) );
  INVX0 U2 ( .INP(eth_top_test_point_11887_in), .ZN(n4) );
  AO22X1 U3 ( .IN1(DataIn[0]), .IN2(n1), .IN3(n2), .IN4(DataOut[0]), .Q(n28)
         );
  AO22X1 U4 ( .IN1(DataIn[1]), .IN2(n1), .IN3(n2), .IN4(DataOut[1]), .Q(n27)
         );
  AO22X1 U5 ( .IN1(DataIn[2]), .IN2(n1), .IN3(n2), .IN4(DataOut[2]), .Q(n26)
         );
  AO22X1 U6 ( .IN1(DataIn[3]), .IN2(n1), .IN3(n2), .IN4(DataOut[3]), .Q(n25)
         );
  AO22X1 U7 ( .IN1(DataIn[4]), .IN2(n1), .IN3(n2), .IN4(DataOut[4]), .Q(n24)
         );
  AO22X1 U8 ( .IN1(DataIn[5]), .IN2(n1), .IN3(n2), .IN4(DataOut[5]), .Q(n23)
         );
  AO22X1 U9 ( .IN1(DataIn[6]), .IN2(n1), .IN3(n2), .IN4(DataOut[6]), .Q(n22)
         );
  AO22X1 U10 ( .IN1(DataIn[7]), .IN2(n1), .IN3(n2), .IN4(DataOut[7]), .Q(n21)
         );
  NOR2X0 U11 ( .IN1(n1), .IN2(SyncReset), .QN(n2) );
  NOR2X0 U12 ( .IN1(n3), .IN2(SyncReset), .QN(n1) );
  INVX0 U13 ( .INP(Write), .ZN(n3) );
endmodule


module eth_register_8_00_test_5 ( DataIn, DataOut, Write, Clk, Reset, 
        SyncReset, eth_top_test_point_11887_in, test_si, test_se );
  input [7:0] DataIn;
  output [7:0] DataOut;
  input Write, Clk, Reset, SyncReset, eth_top_test_point_11887_in, test_si,
         test_se;
  wire   n21, n22, n23, n24, n25, n26, n27, n28, n1, n2, n3, n4;

  SDFFARX1 \DataOut_reg[7]  ( .D(n21), .SI(DataOut[6]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[7]) );
  SDFFARX1 \DataOut_reg[6]  ( .D(n22), .SI(DataOut[5]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[6]) );
  SDFFARX1 \DataOut_reg[5]  ( .D(n23), .SI(DataOut[4]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[5]) );
  SDFFARX1 \DataOut_reg[4]  ( .D(n24), .SI(DataOut[3]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[4]) );
  SDFFARX1 \DataOut_reg[3]  ( .D(n25), .SI(DataOut[2]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[3]) );
  SDFFARX1 \DataOut_reg[2]  ( .D(n26), .SI(DataOut[1]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[2]) );
  SDFFARX1 \DataOut_reg[1]  ( .D(n27), .SI(DataOut[0]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[1]) );
  SDFFARX1 \DataOut_reg[0]  ( .D(n28), .SI(test_si), .SE(test_se), .CLK(Clk), 
        .RSTB(n4), .Q(DataOut[0]) );
  INVX0 U2 ( .INP(eth_top_test_point_11887_in), .ZN(n4) );
  AO22X1 U3 ( .IN1(DataIn[0]), .IN2(n1), .IN3(n2), .IN4(DataOut[0]), .Q(n28)
         );
  AO22X1 U4 ( .IN1(DataIn[1]), .IN2(n1), .IN3(n2), .IN4(DataOut[1]), .Q(n27)
         );
  AO22X1 U5 ( .IN1(DataIn[2]), .IN2(n1), .IN3(n2), .IN4(DataOut[2]), .Q(n26)
         );
  AO22X1 U6 ( .IN1(DataIn[3]), .IN2(n1), .IN3(n2), .IN4(DataOut[3]), .Q(n25)
         );
  AO22X1 U7 ( .IN1(DataIn[4]), .IN2(n1), .IN3(n2), .IN4(DataOut[4]), .Q(n24)
         );
  AO22X1 U8 ( .IN1(DataIn[5]), .IN2(n1), .IN3(n2), .IN4(DataOut[5]), .Q(n23)
         );
  AO22X1 U9 ( .IN1(DataIn[6]), .IN2(n1), .IN3(n2), .IN4(DataOut[6]), .Q(n22)
         );
  AO22X1 U10 ( .IN1(DataIn[7]), .IN2(n1), .IN3(n2), .IN4(DataOut[7]), .Q(n21)
         );
  NOR2X0 U11 ( .IN1(n1), .IN2(SyncReset), .QN(n2) );
  NOR2X0 U12 ( .IN1(n3), .IN2(SyncReset), .QN(n1) );
  INVX0 U13 ( .INP(Write), .ZN(n3) );
endmodule


module eth_register_8_00_test_4 ( DataIn, DataOut, Write, Clk, Reset, 
        SyncReset, eth_top_test_point_11887_in, test_si, test_se );
  input [7:0] DataIn;
  output [7:0] DataOut;
  input Write, Clk, Reset, SyncReset, eth_top_test_point_11887_in, test_si,
         test_se;
  wire   n21, n22, n23, n24, n25, n26, n27, n28, n1, n2, n3, n4;

  SDFFARX1 \DataOut_reg[7]  ( .D(n21), .SI(DataOut[6]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[7]) );
  SDFFARX1 \DataOut_reg[6]  ( .D(n22), .SI(DataOut[5]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[6]) );
  SDFFARX1 \DataOut_reg[5]  ( .D(n23), .SI(DataOut[4]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[5]) );
  SDFFARX1 \DataOut_reg[4]  ( .D(n24), .SI(DataOut[3]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[4]) );
  SDFFARX1 \DataOut_reg[3]  ( .D(n25), .SI(DataOut[2]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[3]) );
  SDFFARX1 \DataOut_reg[2]  ( .D(n26), .SI(DataOut[1]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[2]) );
  SDFFARX1 \DataOut_reg[1]  ( .D(n27), .SI(DataOut[0]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[1]) );
  SDFFARX1 \DataOut_reg[0]  ( .D(n28), .SI(test_si), .SE(test_se), .CLK(Clk), 
        .RSTB(n4), .Q(DataOut[0]) );
  INVX0 U2 ( .INP(eth_top_test_point_11887_in), .ZN(n4) );
  AO22X1 U3 ( .IN1(DataIn[0]), .IN2(n1), .IN3(n2), .IN4(DataOut[0]), .Q(n28)
         );
  AO22X1 U4 ( .IN1(DataIn[1]), .IN2(n1), .IN3(n2), .IN4(DataOut[1]), .Q(n27)
         );
  AO22X1 U5 ( .IN1(DataIn[2]), .IN2(n1), .IN3(n2), .IN4(DataOut[2]), .Q(n26)
         );
  AO22X1 U6 ( .IN1(DataIn[3]), .IN2(n1), .IN3(n2), .IN4(DataOut[3]), .Q(n25)
         );
  AO22X1 U7 ( .IN1(DataIn[4]), .IN2(n1), .IN3(n2), .IN4(DataOut[4]), .Q(n24)
         );
  AO22X1 U8 ( .IN1(DataIn[5]), .IN2(n1), .IN3(n2), .IN4(DataOut[5]), .Q(n23)
         );
  AO22X1 U9 ( .IN1(DataIn[6]), .IN2(n1), .IN3(n2), .IN4(DataOut[6]), .Q(n22)
         );
  AO22X1 U10 ( .IN1(DataIn[7]), .IN2(n1), .IN3(n2), .IN4(DataOut[7]), .Q(n21)
         );
  NOR2X0 U11 ( .IN1(n1), .IN2(SyncReset), .QN(n2) );
  NOR2X0 U12 ( .IN1(n3), .IN2(SyncReset), .QN(n1) );
  INVX0 U13 ( .INP(Write), .ZN(n3) );
endmodule


module eth_register_8_00_test_3 ( DataIn, DataOut, Write, Clk, Reset, 
        SyncReset, eth_top_test_point_11887_in, test_si, test_se );
  input [7:0] DataIn;
  output [7:0] DataOut;
  input Write, Clk, Reset, SyncReset, eth_top_test_point_11887_in, test_si,
         test_se;
  wire   n21, n22, n23, n24, n25, n26, n27, n28, n1, n2, n3, n4;

  SDFFARX1 \DataOut_reg[7]  ( .D(n21), .SI(DataOut[6]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[7]) );
  SDFFARX1 \DataOut_reg[6]  ( .D(n22), .SI(DataOut[5]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[6]) );
  SDFFARX1 \DataOut_reg[5]  ( .D(n23), .SI(DataOut[4]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[5]) );
  SDFFARX1 \DataOut_reg[4]  ( .D(n24), .SI(DataOut[3]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[4]) );
  SDFFARX1 \DataOut_reg[3]  ( .D(n25), .SI(DataOut[2]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[3]) );
  SDFFARX1 \DataOut_reg[2]  ( .D(n26), .SI(DataOut[1]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[2]) );
  SDFFARX1 \DataOut_reg[1]  ( .D(n27), .SI(DataOut[0]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[1]) );
  SDFFARX1 \DataOut_reg[0]  ( .D(n28), .SI(test_si), .SE(test_se), .CLK(Clk), 
        .RSTB(n4), .Q(DataOut[0]) );
  INVX0 U2 ( .INP(eth_top_test_point_11887_in), .ZN(n4) );
  AO22X1 U3 ( .IN1(DataIn[0]), .IN2(n1), .IN3(n2), .IN4(DataOut[0]), .Q(n28)
         );
  AO22X1 U4 ( .IN1(DataIn[1]), .IN2(n1), .IN3(n2), .IN4(DataOut[1]), .Q(n27)
         );
  AO22X1 U5 ( .IN1(DataIn[2]), .IN2(n1), .IN3(n2), .IN4(DataOut[2]), .Q(n26)
         );
  AO22X1 U6 ( .IN1(DataIn[3]), .IN2(n1), .IN3(n2), .IN4(DataOut[3]), .Q(n25)
         );
  AO22X1 U7 ( .IN1(DataIn[4]), .IN2(n1), .IN3(n2), .IN4(DataOut[4]), .Q(n24)
         );
  AO22X1 U8 ( .IN1(DataIn[5]), .IN2(n1), .IN3(n2), .IN4(DataOut[5]), .Q(n23)
         );
  AO22X1 U9 ( .IN1(DataIn[6]), .IN2(n1), .IN3(n2), .IN4(DataOut[6]), .Q(n22)
         );
  AO22X1 U10 ( .IN1(DataIn[7]), .IN2(n1), .IN3(n2), .IN4(DataOut[7]), .Q(n21)
         );
  NOR2X0 U11 ( .IN1(n1), .IN2(SyncReset), .QN(n2) );
  NOR2X0 U12 ( .IN1(n3), .IN2(SyncReset), .QN(n1) );
  INVX0 U13 ( .INP(Write), .ZN(n3) );
endmodule


module eth_register_8_00_test_2 ( DataIn, DataOut, Write, Clk, Reset, 
        SyncReset, eth_top_test_point_11887_in, test_si, test_se );
  input [7:0] DataIn;
  output [7:0] DataOut;
  input Write, Clk, Reset, SyncReset, eth_top_test_point_11887_in, test_si,
         test_se;
  wire   n21, n22, n23, n24, n25, n26, n27, n28, n1, n2, n3, n4;

  SDFFARX1 \DataOut_reg[7]  ( .D(n21), .SI(DataOut[6]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[7]) );
  SDFFARX1 \DataOut_reg[6]  ( .D(n22), .SI(DataOut[5]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[6]) );
  SDFFARX1 \DataOut_reg[5]  ( .D(n23), .SI(DataOut[4]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[5]) );
  SDFFARX1 \DataOut_reg[4]  ( .D(n24), .SI(DataOut[3]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[4]) );
  SDFFARX1 \DataOut_reg[3]  ( .D(n25), .SI(DataOut[2]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[3]) );
  SDFFARX1 \DataOut_reg[2]  ( .D(n26), .SI(DataOut[1]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[2]) );
  SDFFARX1 \DataOut_reg[1]  ( .D(n27), .SI(DataOut[0]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[1]) );
  SDFFARX1 \DataOut_reg[0]  ( .D(n28), .SI(test_si), .SE(test_se), .CLK(Clk), 
        .RSTB(n4), .Q(DataOut[0]) );
  INVX0 U2 ( .INP(eth_top_test_point_11887_in), .ZN(n4) );
  AO22X1 U3 ( .IN1(DataIn[0]), .IN2(n1), .IN3(n2), .IN4(DataOut[0]), .Q(n28)
         );
  AO22X1 U4 ( .IN1(DataIn[1]), .IN2(n1), .IN3(n2), .IN4(DataOut[1]), .Q(n27)
         );
  AO22X1 U5 ( .IN1(DataIn[2]), .IN2(n1), .IN3(n2), .IN4(DataOut[2]), .Q(n26)
         );
  AO22X1 U6 ( .IN1(DataIn[3]), .IN2(n1), .IN3(n2), .IN4(DataOut[3]), .Q(n25)
         );
  AO22X1 U7 ( .IN1(DataIn[4]), .IN2(n1), .IN3(n2), .IN4(DataOut[4]), .Q(n24)
         );
  AO22X1 U8 ( .IN1(DataIn[5]), .IN2(n1), .IN3(n2), .IN4(DataOut[5]), .Q(n23)
         );
  AO22X1 U9 ( .IN1(DataIn[6]), .IN2(n1), .IN3(n2), .IN4(DataOut[6]), .Q(n22)
         );
  AO22X1 U10 ( .IN1(DataIn[7]), .IN2(n1), .IN3(n2), .IN4(DataOut[7]), .Q(n21)
         );
  NOR2X0 U11 ( .IN1(n1), .IN2(SyncReset), .QN(n2) );
  NOR2X0 U12 ( .IN1(n3), .IN2(SyncReset), .QN(n1) );
  INVX0 U13 ( .INP(Write), .ZN(n3) );
endmodule


module eth_register_8_00_test_1 ( DataIn, DataOut, Write, Clk, Reset, 
        SyncReset, eth_top_test_point_11887_in, test_si, test_se );
  input [7:0] DataIn;
  output [7:0] DataOut;
  input Write, Clk, Reset, SyncReset, eth_top_test_point_11887_in, test_si,
         test_se;
  wire   n21, n22, n23, n24, n25, n26, n27, n28, n1, n2, n3, n4;

  SDFFARX1 \DataOut_reg[7]  ( .D(n21), .SI(DataOut[6]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[7]) );
  SDFFARX1 \DataOut_reg[6]  ( .D(n22), .SI(DataOut[5]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[6]) );
  SDFFARX1 \DataOut_reg[5]  ( .D(n23), .SI(DataOut[4]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[5]) );
  SDFFARX1 \DataOut_reg[4]  ( .D(n24), .SI(DataOut[3]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[4]) );
  SDFFARX1 \DataOut_reg[3]  ( .D(n25), .SI(DataOut[2]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[3]) );
  SDFFARX1 \DataOut_reg[2]  ( .D(n26), .SI(DataOut[1]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[2]) );
  SDFFARX1 \DataOut_reg[1]  ( .D(n27), .SI(DataOut[0]), .SE(test_se), .CLK(Clk), .RSTB(n4), .Q(DataOut[1]) );
  SDFFARX1 \DataOut_reg[0]  ( .D(n28), .SI(test_si), .SE(test_se), .CLK(Clk), 
        .RSTB(n4), .Q(DataOut[0]) );
  INVX0 U2 ( .INP(eth_top_test_point_11887_in), .ZN(n4) );
  AO22X1 U3 ( .IN1(DataIn[0]), .IN2(n1), .IN3(n2), .IN4(DataOut[0]), .Q(n28)
         );
  AO22X1 U4 ( .IN1(DataIn[1]), .IN2(n1), .IN3(n2), .IN4(DataOut[1]), .Q(n27)
         );
  AO22X1 U5 ( .IN1(DataIn[2]), .IN2(n1), .IN3(n2), .IN4(DataOut[2]), .Q(n26)
         );
  AO22X1 U6 ( .IN1(DataIn[3]), .IN2(n1), .IN3(n2), .IN4(DataOut[3]), .Q(n25)
         );
  AO22X1 U7 ( .IN1(DataIn[4]), .IN2(n1), .IN3(n2), .IN4(DataOut[4]), .Q(n24)
         );
  AO22X1 U8 ( .IN1(DataIn[5]), .IN2(n1), .IN3(n2), .IN4(DataOut[5]), .Q(n23)
         );
  AO22X1 U9 ( .IN1(DataIn[6]), .IN2(n1), .IN3(n2), .IN4(DataOut[6]), .Q(n22)
         );
  AO22X1 U10 ( .IN1(DataIn[7]), .IN2(n1), .IN3(n2), .IN4(DataOut[7]), .Q(n21)
         );
  NOR2X0 U11 ( .IN1(n1), .IN2(SyncReset), .QN(n2) );
  NOR2X0 U12 ( .IN1(n3), .IN2(SyncReset), .QN(n1) );
  INVX0 U13 ( .INP(Write), .ZN(n3) );
endmodule


module eth_register_1_0_test_1 ( DataIn, DataOut, Write, Clk, Reset, SyncReset, 
        eth_top_test_point_11887_in, test_si, test_se );
  input [0:0] DataIn;
  output [0:0] DataOut;
  input Write, Clk, Reset, SyncReset, eth_top_test_point_11887_in, test_si,
         test_se;
  wire   n6, n1, n2, n3;

  SDFFARX1 \DataOut_reg[0]  ( .D(n6), .SI(test_si), .SE(test_se), .CLK(Clk), 
        .RSTB(n3), .Q(DataOut[0]) );
  INVX0 U2 ( .INP(eth_top_test_point_11887_in), .ZN(n3) );
  NOR2X0 U3 ( .IN1(SyncReset), .IN2(n1), .QN(n6) );
  INVX0 U4 ( .INP(n2), .ZN(n1) );
  MUX21X1 U5 ( .IN1(DataOut[0]), .IN2(DataIn[0]), .S(Write), .Q(n2) );
endmodule


module eth_registers_test_1 ( DataIn, Address, Rw, Cs, Clk, Reset, DataOut, 
        r_RecSmall, r_Pad, r_HugEn, r_CrcEn, r_DlyCrcEn, r_FullD, r_ExDfrEn, 
        r_NoBckof, r_LoopBck, r_IFG, r_Pro, r_Iam, r_Bro, r_NoPre, r_TxEn, 
        r_RxEn, TxB_IRQ, TxE_IRQ, RxB_IRQ, RxE_IRQ, Busy_IRQ, r_IPGT, r_IPGR1, 
        r_IPGR2, r_MinFL, r_MaxFL, r_MaxRet, r_CollValid, r_TxFlow, r_RxFlow, 
        r_PassAll, r_MiiNoPre, r_ClkDiv, r_WCtrlData, r_RStat, r_ScanStat, 
        r_RGAD, r_FIAD, r_CtrlData, NValid_stat, Busy_stat, LinkFail, r_MAC, 
        WCtrlDataStart, RStatStart, UpdateMIIRX_DATAReg, Prsd, r_TxBDNum, 
        int_o, r_HASH0, r_HASH1, r_TxPauseTV, r_TxPauseRq, RstTxPauseRq, 
        TxCtrlEndFrm, StartTxDone, TxClk, RxClk, SetPauseTimer, 
        eth_top_test_point_11887_in, test_si, test_so, test_se );
  input [31:0] DataIn;
  input [7:0] Address;
  input [3:0] Cs;
  output [31:0] DataOut;
  output [6:0] r_IPGT;
  output [6:0] r_IPGR1;
  output [6:0] r_IPGR2;
  output [15:0] r_MinFL;
  output [15:0] r_MaxFL;
  output [3:0] r_MaxRet;
  output [5:0] r_CollValid;
  output [7:0] r_ClkDiv;
  output [4:0] r_RGAD;
  output [4:0] r_FIAD;
  output [15:0] r_CtrlData;
  output [47:0] r_MAC;
  input [15:0] Prsd;
  output [7:0] r_TxBDNum;
  output [31:0] r_HASH0;
  output [31:0] r_HASH1;
  output [15:0] r_TxPauseTV;
  input Rw, Clk, Reset, TxB_IRQ, TxE_IRQ, RxB_IRQ, RxE_IRQ, Busy_IRQ,
         NValid_stat, Busy_stat, LinkFail, WCtrlDataStart, RStatStart,
         UpdateMIIRX_DATAReg, RstTxPauseRq, TxCtrlEndFrm, StartTxDone, TxClk,
         RxClk, SetPauseTimer, eth_top_test_point_11887_in, test_si, test_se;
  output r_RecSmall, r_Pad, r_HugEn, r_CrcEn, r_DlyCrcEn, r_FullD, r_ExDfrEn,
         r_NoBckof, r_LoopBck, r_IFG, r_Pro, r_Iam, r_Bro, r_NoPre, r_TxEn,
         r_RxEn, r_TxFlow, r_RxFlow, r_PassAll, r_MiiNoPre, r_WCtrlData,
         r_RStat, r_ScanStat, int_o, r_TxPauseRq, test_so;
  wire   \INT_MASK_Wr[0] , \IPGT_Wr[0] , \IPGR1_Wr[0] , \IPGR2_Wr[0] ,
         \COLLCONF_Wr[2] , COLLCONF_Wr_0, \CTRLMODER_Wr[0] ,
         \MIICOMMAND_Wr[0] , \TX_BD_NUM_Wr[0] , MODEROut_11, SetTxCIrq_txclk,
         ResetTxCIrq_sync2, SetTxCIrq_sync1, SetTxCIrq_sync2, SetTxCIrq_sync3,
         N179, SetRxCIrq_rxclk, ResetRxCIrq_sync2, SetRxCIrq_sync1,
         SetRxCIrq_sync2, SetRxCIrq_sync3, N185, ResetRxCIrq_sync1, n30, n31,
         n32, n33, n241, n242, n243, n244, n245, n246, n247, n248, n249, n1,
         n2, n3, n4, n5, n6, n27, n265, n266, n270, n271, n272, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n28, n29, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240;
  wire   [2:0] MODER_Wr;
  wire   [3:0] PACKETLEN_Wr;
  wire   [1:0] MIIMODER_Wr;
  wire   [1:0] MIIADDRESS_Wr;
  wire   [1:0] MIITX_DATA_Wr;
  wire   [3:0] MAC_ADDR0_Wr;
  wire   [1:0] MAC_ADDR1_Wr;
  wire   [3:0] HASH0_Wr;
  wire   [3:0] HASH1_Wr;
  wire   [2:0] TXCTRL_Wr;
  wire   [1:0] MODEROut;
  wire   [6:0] INT_MASKOut;
  wire   [15:0] MIIRX_DATAOut;
  assign test_so = n3;

  SDFFARX1 ResetTxCIrq_sync2_reg ( .D(SetTxCIrq_sync1), .SI(n272), .SE(test_se), .CLK(TxClk), .RSTB(n240), .Q(ResetTxCIrq_sync2) );
  SDFFARX1 SetTxCIrq_txclk_reg ( .D(n249), .SI(SetTxCIrq_sync3), .SE(test_se), 
        .CLK(TxClk), .RSTB(n240), .Q(SetTxCIrq_txclk), .QN(n30) );
  SDFFARX1 SetTxCIrq_sync1_reg ( .D(SetTxCIrq_txclk), .SI(n270), .SE(test_se), 
        .CLK(n12), .RSTB(n240), .Q(SetTxCIrq_sync1) );
  SDFFARX1 SetTxCIrq_sync2_reg ( .D(SetTxCIrq_sync1), .SI(SetTxCIrq_sync1), 
        .SE(test_se), .CLK(n12), .RSTB(n240), .Q(SetTxCIrq_sync2), .QN(n31) );
  SDFFARX1 SetTxCIrq_sync3_reg ( .D(SetTxCIrq_sync2), .SI(SetTxCIrq_sync2), 
        .SE(test_se), .CLK(n12), .RSTB(n240), .Q(SetTxCIrq_sync3) );
  SDFFARX1 SetTxCIrq_reg ( .D(N179), .SI(SetRxCIrq_sync3), .SE(test_se), .CLK(
        n12), .RSTB(n240), .Q(n270), .QN(n266) );
  SDFFARX1 ResetRxCIrq_sync3_reg ( .D(ResetRxCIrq_sync2), .SI(
        ResetRxCIrq_sync2), .SE(test_se), .CLK(RxClk), .RSTB(n240), .Q(n272), 
        .QN(n33) );
  SDFFARX1 SetRxCIrq_rxclk_reg ( .D(n248), .SI(n271), .SE(test_se), .CLK(RxClk), .RSTB(n240), .Q(SetRxCIrq_rxclk) );
  SDFFARX1 SetRxCIrq_sync1_reg ( .D(SetRxCIrq_rxclk), .SI(SetRxCIrq_rxclk), 
        .SE(test_se), .CLK(n12), .RSTB(n240), .Q(SetRxCIrq_sync1) );
  SDFFARX1 SetRxCIrq_sync2_reg ( .D(SetRxCIrq_sync1), .SI(SetRxCIrq_sync1), 
        .SE(test_se), .CLK(n12), .RSTB(n240), .Q(SetRxCIrq_sync2), .QN(n32) );
  SDFFARX1 SetRxCIrq_sync3_reg ( .D(SetRxCIrq_sync2), .SI(SetRxCIrq_sync2), 
        .SE(test_se), .CLK(n12), .RSTB(n240), .Q(SetRxCIrq_sync3) );
  SDFFARX1 ResetRxCIrq_sync1_reg ( .D(SetRxCIrq_sync2), .SI(r_HASH1[31]), .SE(
        test_se), .CLK(RxClk), .RSTB(n240), .Q(ResetRxCIrq_sync1) );
  SDFFARX1 ResetRxCIrq_sync2_reg ( .D(ResetRxCIrq_sync1), .SI(
        ResetRxCIrq_sync1), .SE(test_se), .CLK(RxClk), .RSTB(n240), .Q(
        ResetRxCIrq_sync2) );
  SDFFARX1 SetRxCIrq_reg ( .D(N185), .SI(ResetTxCIrq_sync2), .SE(test_se), 
        .CLK(n12), .RSTB(n240), .Q(n271), .QN(n265) );
  SDFFARX1 irq_txb_reg ( .D(n247), .SI(n2), .SE(test_se), .CLK(n12), .RSTB(
        n240), .Q(n6) );
  SDFFARX1 irq_txe_reg ( .D(n246), .SI(n4), .SE(test_se), .CLK(n12), .RSTB(
        n240), .Q(n3) );
  SDFFARX1 irq_rxb_reg ( .D(n245), .SI(n1), .SE(test_se), .CLK(n12), .RSTB(
        n240), .Q(n5) );
  SDFFARX1 irq_rxe_reg ( .D(n244), .SI(n27), .SE(test_se), .CLK(n12), .RSTB(
        n240), .Q(n2) );
  SDFFARX1 irq_busy_reg ( .D(n243), .SI(r_TxBDNum[7]), .SE(test_se), .CLK(n12), 
        .RSTB(n240), .Q(n1) );
  SDFFARX1 irq_txc_reg ( .D(n242), .SI(n6), .SE(test_se), .CLK(n12), .RSTB(
        n240), .Q(n4), .QN(n239) );
  SDFFARX1 irq_rxc_reg ( .D(n241), .SI(n5), .SE(test_se), .CLK(n12), .RSTB(
        n240), .Q(n27), .QN(n238) );
  eth_register_8_00_test_0 MODER_0 ( .DataIn(DataIn[7:0]), .DataOut({r_LoopBck, 
        r_IFG, r_Pro, r_Iam, r_Bro, r_NoPre, MODEROut}), .Write(MODER_Wr[0]), 
        .Clk(n8), .Reset(Reset), .SyncReset(1'b0), 
        .eth_top_test_point_11887_in(eth_top_test_point_11887_in), .test_si(
        r_CtrlData[15]), .test_se(test_se) );
  eth_register_8_a0_test_1 MODER_1 ( .DataIn(DataIn[15:8]), .DataOut({r_Pad, 
        r_HugEn, r_CrcEn, r_DlyCrcEn, MODEROut_11, r_FullD, r_ExDfrEn, 
        r_NoBckof}), .Write(MODER_Wr[1]), .Clk(n7), .Reset(Reset), .SyncReset(
        1'b0), .eth_top_test_point_11887_in(eth_top_test_point_11887_in), 
        .test_si(r_LoopBck), .test_se(test_se) );
  eth_register_1_0_test_0 MODER_2 ( .DataIn(DataIn[16]), .DataOut(r_RecSmall), 
        .Write(MODER_Wr[2]), .Clk(n12), .Reset(Reset), .SyncReset(1'b0), 
        .eth_top_test_point_11887_in(eth_top_test_point_11887_in), .test_si(
        r_Pad), .test_se(test_se) );
  eth_register_7_00_test_1 INT_MASK_0 ( .DataIn(DataIn[6:0]), .DataOut(
        INT_MASKOut), .Write(\INT_MASK_Wr[0] ), .Clk(n12), .Reset(Reset), 
        .SyncReset(1'b0), .eth_top_test_point_11887_in(
        eth_top_test_point_11887_in), .test_si(r_TxFlow), .test_se(test_se) );
  eth_register_7_12_test_0 IPGT_0 ( .DataIn(DataIn[6:0]), .DataOut(r_IPGT), 
        .Write(\IPGT_Wr[0] ), .Clk(n11), .Reset(Reset), .SyncReset(1'b0), 
        .eth_top_test_point_11887_in(eth_top_test_point_11887_in), .test_si(
        r_IPGR2[6]), .test_se(test_se) );
  eth_register_7_0c_test_1 IPGR1_0 ( .DataIn(DataIn[6:0]), .DataOut(r_IPGR1), 
        .Write(\IPGR1_Wr[0] ), .Clk(n12), .Reset(Reset), .SyncReset(1'b0), 
        .eth_top_test_point_11887_in(eth_top_test_point_11887_in), .test_si(
        INT_MASKOut[6]), .test_se(test_se) );
  eth_register_7_12_test_1 IPGR2_0 ( .DataIn(DataIn[6:0]), .DataOut(r_IPGR2), 
        .Write(\IPGR2_Wr[0] ), .Clk(n11), .Reset(Reset), .SyncReset(1'b0), 
        .eth_top_test_point_11887_in(eth_top_test_point_11887_in), .test_si(
        r_IPGR1[6]), .test_se(test_se) );
  eth_register_8_00_test_20 PACKETLEN_0 ( .DataIn(DataIn[7:0]), .DataOut(
        r_MaxFL[7:0]), .Write(PACKETLEN_Wr[0]), .Clk(n11), .Reset(Reset), 
        .SyncReset(1'b0), .eth_top_test_point_11887_in(
        eth_top_test_point_11887_in), .test_si(r_RecSmall), .test_se(test_se)
         );
  eth_register_8_06_test_1 PACKETLEN_1 ( .DataIn(DataIn[15:8]), .DataOut(
        r_MaxFL[15:8]), .Write(PACKETLEN_Wr[1]), .Clk(n7), .Reset(Reset), 
        .SyncReset(1'b0), .eth_top_test_point_11887_in(
        eth_top_test_point_11887_in), .test_si(r_MaxFL[7]), .test_se(test_se)
         );
  eth_register_8_40_test_0 PACKETLEN_2 ( .DataIn(DataIn[23:16]), .DataOut(
        r_MinFL[7:0]), .Write(PACKETLEN_Wr[2]), .Clk(n8), .Reset(Reset), 
        .SyncReset(1'b0), .eth_top_test_point_11887_in(
        eth_top_test_point_11887_in), .test_si(r_MaxFL[15]), .test_se(test_se)
         );
  eth_register_8_00_test_19 PACKETLEN_3 ( .DataIn(DataIn[31:24]), .DataOut(
        r_MinFL[15:8]), .Write(PACKETLEN_Wr[3]), .Clk(n11), .Reset(Reset), 
        .SyncReset(1'b0), .eth_top_test_point_11887_in(
        eth_top_test_point_11887_in), .test_si(r_MinFL[7]), .test_se(test_se)
         );
  eth_register_6_3f_test_1 COLLCONF_0 ( .DataIn(DataIn[5:0]), .DataOut(
        r_CollValid), .Write(COLLCONF_Wr_0), .Clk(n11), .Reset(Reset), 
        .SyncReset(1'b0), .eth_top_test_point_11887_in(
        eth_top_test_point_11887_in), .test_si(test_si), .test_se(test_se) );
  eth_register_4_f_test_1 COLLCONF_2 ( .DataIn(DataIn[19:16]), .DataOut(
        r_MaxRet), .Write(\COLLCONF_Wr[2] ), .Clk(n10), .Reset(Reset), 
        .SyncReset(1'b0), .eth_top_test_point_11887_in(
        eth_top_test_point_11887_in), .test_si(r_CollValid[5]), .test_se(
        test_se) );
  eth_register_8_40_test_1 TX_BD_NUM_0 ( .DataIn(DataIn[7:0]), .DataOut(
        r_TxBDNum), .Write(\TX_BD_NUM_Wr[0] ), .Clk(n7), .Reset(Reset), 
        .SyncReset(1'b0), .eth_top_test_point_11887_in(
        eth_top_test_point_11887_in), .test_si(r_TxPauseRq), .test_se(test_se)
         );
  eth_register_3_0_test_1 CTRLMODER_0 ( .DataIn(DataIn[2:0]), .DataOut({
        r_TxFlow, r_RxFlow, r_PassAll}), .Write(\CTRLMODER_Wr[0] ), .Clk(n12), 
        .Reset(Reset), .SyncReset(1'b0), .eth_top_test_point_11887_in(
        eth_top_test_point_11887_in), .test_si(r_MaxRet[3]), .test_se(test_se)
         );
  eth_register_8_64_test_1 MIIMODER_0 ( .DataIn(DataIn[7:0]), .DataOut(
        r_ClkDiv), .Write(MIIMODER_Wr[0]), .Clk(n7), .Reset(Reset), 
        .SyncReset(1'b0), .eth_top_test_point_11887_in(
        eth_top_test_point_11887_in), .test_si(r_WCtrlData), .test_se(test_se)
         );
  eth_register_1_0_test_2 MIIMODER_1 ( .DataIn(DataIn[8]), .DataOut(r_MiiNoPre), .Write(MIIMODER_Wr[1]), .Clk(n12), .Reset(Reset), .SyncReset(1'b0), 
        .eth_top_test_point_11887_in(eth_top_test_point_11887_in), .test_si(
        r_ClkDiv[7]), .test_se(test_se) );
  eth_register_WIDTH1_RESET_VALUE0_test_0 MIICOMMAND0 ( .DataIn(DataIn[0]), 
        .DataOut(r_ScanStat), .Write(\MIICOMMAND_Wr[0] ), .Clk(n12), .Reset(
        Reset), .SyncReset(1'b0), .eth_top_test_point_11887_in(
        eth_top_test_point_11887_in), .test_si(r_RGAD[4]), .test_se(test_se)
         );
  eth_register_WIDTH1_RESET_VALUE0_test_2 MIICOMMAND1 ( .DataIn(DataIn[1]), 
        .DataOut(r_RStat), .Write(\MIICOMMAND_Wr[0] ), .Clk(n12), .Reset(Reset), .SyncReset(RStatStart), .eth_top_test_point_11887_in(
        eth_top_test_point_11887_in), .test_si(r_ScanStat), .test_se(test_se)
         );
  eth_register_WIDTH1_RESET_VALUE0_test_1 MIICOMMAND2 ( .DataIn(DataIn[2]), 
        .DataOut(r_WCtrlData), .Write(\MIICOMMAND_Wr[0] ), .Clk(n12), .Reset(
        Reset), .SyncReset(WCtrlDataStart), .eth_top_test_point_11887_in(
        eth_top_test_point_11887_in), .test_si(r_RStat), .test_se(test_se) );
  eth_register_5_00_test_0 MIIADDRESS_0 ( .DataIn(DataIn[4:0]), .DataOut(
        r_FIAD), .Write(MIIADDRESS_Wr[0]), .Clk(n9), .Reset(Reset), 
        .SyncReset(1'b0), .eth_top_test_point_11887_in(
        eth_top_test_point_11887_in), .test_si(r_MAC[47]), .test_se(test_se)
         );
  eth_register_5_00_test_1 MIIADDRESS_1 ( .DataIn(DataIn[12:8]), .DataOut(
        r_RGAD), .Write(MIIADDRESS_Wr[1]), .Clk(n8), .Reset(Reset), 
        .SyncReset(1'b0), .eth_top_test_point_11887_in(
        eth_top_test_point_11887_in), .test_si(r_FIAD[4]), .test_se(test_se)
         );
  eth_register_8_00_test_18 MIITX_DATA_0 ( .DataIn(DataIn[7:0]), .DataOut(
        r_CtrlData[7:0]), .Write(MIITX_DATA_Wr[0]), .Clk(n11), .Reset(Reset), 
        .SyncReset(1'b0), .eth_top_test_point_11887_in(
        eth_top_test_point_11887_in), .test_si(MIIRX_DATAOut[15]), .test_se(
        test_se) );
  eth_register_8_00_test_17 MIITX_DATA_1 ( .DataIn(DataIn[15:8]), .DataOut(
        r_CtrlData[15:8]), .Write(MIITX_DATA_Wr[1]), .Clk(n10), .Reset(Reset), 
        .SyncReset(1'b0), .eth_top_test_point_11887_in(
        eth_top_test_point_11887_in), .test_si(r_CtrlData[7]), .test_se(
        test_se) );
  eth_register_16_0000_test_1 MIIRX_DATA ( .DataIn(Prsd), .DataOut(
        MIIRX_DATAOut), .Write(UpdateMIIRX_DATAReg), .Clk(n7), .Reset(Reset), 
        .SyncReset(1'b0), .eth_top_test_point_11887_in(
        eth_top_test_point_11887_in), .test_si(r_MiiNoPre), .test_se(test_se)
         );
  eth_register_8_00_test_16 MAC_ADDR0_0 ( .DataIn(DataIn[7:0]), .DataOut(
        r_MAC[7:0]), .Write(MAC_ADDR0_Wr[0]), .Clk(n10), .Reset(Reset), 
        .SyncReset(1'b0), .eth_top_test_point_11887_in(
        eth_top_test_point_11887_in), .test_si(r_IPGT[6]), .test_se(test_se)
         );
  eth_register_8_00_test_15 MAC_ADDR0_1 ( .DataIn(DataIn[15:8]), .DataOut(
        r_MAC[15:8]), .Write(MAC_ADDR0_Wr[1]), .Clk(n11), .Reset(Reset), 
        .SyncReset(1'b0), .eth_top_test_point_11887_in(
        eth_top_test_point_11887_in), .test_si(r_MAC[7]), .test_se(test_se) );
  eth_register_8_00_test_14 MAC_ADDR0_2 ( .DataIn(DataIn[23:16]), .DataOut(
        r_MAC[23:16]), .Write(MAC_ADDR0_Wr[2]), .Clk(n10), .Reset(Reset), 
        .SyncReset(1'b0), .eth_top_test_point_11887_in(
        eth_top_test_point_11887_in), .test_si(r_MAC[15]), .test_se(test_se)
         );
  eth_register_8_00_test_13 MAC_ADDR0_3 ( .DataIn(DataIn[31:24]), .DataOut(
        r_MAC[31:24]), .Write(MAC_ADDR0_Wr[3]), .Clk(n10), .Reset(Reset), 
        .SyncReset(1'b0), .eth_top_test_point_11887_in(
        eth_top_test_point_11887_in), .test_si(r_MAC[23]), .test_se(test_se)
         );
  eth_register_8_00_test_12 MAC_ADDR1_0 ( .DataIn(DataIn[7:0]), .DataOut(
        r_MAC[39:32]), .Write(MAC_ADDR1_Wr[0]), .Clk(n10), .Reset(Reset), 
        .SyncReset(1'b0), .eth_top_test_point_11887_in(
        eth_top_test_point_11887_in), .test_si(r_MAC[31]), .test_se(test_se)
         );
  eth_register_8_00_test_11 MAC_ADDR1_1 ( .DataIn(DataIn[15:8]), .DataOut(
        r_MAC[47:40]), .Write(MAC_ADDR1_Wr[1]), .Clk(n9), .Reset(Reset), 
        .SyncReset(1'b0), .eth_top_test_point_11887_in(
        eth_top_test_point_11887_in), .test_si(r_MAC[39]), .test_se(test_se)
         );
  eth_register_8_00_test_10 RXHASH0_0 ( .DataIn(DataIn[7:0]), .DataOut(
        r_HASH0[7:0]), .Write(HASH0_Wr[0]), .Clk(n9), .Reset(Reset), 
        .SyncReset(1'b0), .eth_top_test_point_11887_in(
        eth_top_test_point_11887_in), .test_si(r_MinFL[15]), .test_se(test_se)
         );
  eth_register_8_00_test_9 RXHASH0_1 ( .DataIn(DataIn[15:8]), .DataOut(
        r_HASH0[15:8]), .Write(HASH0_Wr[1]), .Clk(n9), .Reset(Reset), 
        .SyncReset(1'b0), .eth_top_test_point_11887_in(
        eth_top_test_point_11887_in), .test_si(r_HASH0[7]), .test_se(test_se)
         );
  eth_register_8_00_test_8 RXHASH0_2 ( .DataIn(DataIn[23:16]), .DataOut(
        r_HASH0[23:16]), .Write(HASH0_Wr[2]), .Clk(n9), .Reset(Reset), 
        .SyncReset(1'b0), .eth_top_test_point_11887_in(
        eth_top_test_point_11887_in), .test_si(r_HASH0[15]), .test_se(test_se)
         );
  eth_register_8_00_test_7 RXHASH0_3 ( .DataIn(DataIn[31:24]), .DataOut(
        r_HASH0[31:24]), .Write(HASH0_Wr[3]), .Clk(n9), .Reset(Reset), 
        .SyncReset(1'b0), .eth_top_test_point_11887_in(
        eth_top_test_point_11887_in), .test_si(r_HASH0[23]), .test_se(test_se)
         );
  eth_register_8_00_test_6 RXHASH1_0 ( .DataIn(DataIn[7:0]), .DataOut(
        r_HASH1[7:0]), .Write(HASH1_Wr[0]), .Clk(n8), .Reset(Reset), 
        .SyncReset(1'b0), .eth_top_test_point_11887_in(
        eth_top_test_point_11887_in), .test_si(r_HASH0[31]), .test_se(test_se)
         );
  eth_register_8_00_test_5 RXHASH1_1 ( .DataIn(DataIn[15:8]), .DataOut(
        r_HASH1[15:8]), .Write(HASH1_Wr[1]), .Clk(n8), .Reset(Reset), 
        .SyncReset(1'b0), .eth_top_test_point_11887_in(
        eth_top_test_point_11887_in), .test_si(r_HASH1[7]), .test_se(test_se)
         );
  eth_register_8_00_test_4 RXHASH1_2 ( .DataIn(DataIn[23:16]), .DataOut(
        r_HASH1[23:16]), .Write(HASH1_Wr[2]), .Clk(n8), .Reset(Reset), 
        .SyncReset(1'b0), .eth_top_test_point_11887_in(
        eth_top_test_point_11887_in), .test_si(r_HASH1[15]), .test_se(test_se)
         );
  eth_register_8_00_test_3 RXHASH1_3 ( .DataIn(DataIn[31:24]), .DataOut(
        r_HASH1[31:24]), .Write(HASH1_Wr[3]), .Clk(n10), .Reset(Reset), 
        .SyncReset(1'b0), .eth_top_test_point_11887_in(
        eth_top_test_point_11887_in), .test_si(r_HASH1[23]), .test_se(test_se)
         );
  eth_register_8_00_test_2 TXCTRL_0 ( .DataIn(DataIn[7:0]), .DataOut(
        r_TxPauseTV[7:0]), .Write(TXCTRL_Wr[0]), .Clk(n9), .Reset(Reset), 
        .SyncReset(1'b0), .eth_top_test_point_11887_in(
        eth_top_test_point_11887_in), .test_si(SetTxCIrq_txclk), .test_se(
        test_se) );
  eth_register_8_00_test_1 TXCTRL_1 ( .DataIn(DataIn[15:8]), .DataOut(
        r_TxPauseTV[15:8]), .Write(TXCTRL_Wr[1]), .Clk(n8), .Reset(Reset), 
        .SyncReset(1'b0), .eth_top_test_point_11887_in(
        eth_top_test_point_11887_in), .test_si(r_TxPauseTV[7]), .test_se(
        test_se) );
  eth_register_1_0_test_1 TXCTRL_2 ( .DataIn(DataIn[16]), .DataOut(r_TxPauseRq), .Write(TXCTRL_Wr[2]), .Clk(n12), .Reset(Reset), .SyncReset(RstTxPauseRq), 
        .eth_top_test_point_11887_in(eth_top_test_point_11887_in), .test_si(
        r_TxPauseTV[15]), .test_se(test_se) );
  NBUFFX4 U3 ( .INP(Clk), .Z(n8) );
  NBUFFX4 U4 ( .INP(Clk), .Z(n9) );
  NBUFFX4 U5 ( .INP(Clk), .Z(n11) );
  NBUFFX4 U6 ( .INP(Clk), .Z(n10) );
  NBUFFX4 U7 ( .INP(Clk), .Z(n7) );
  NBUFFX4 U8 ( .INP(Clk), .Z(n12) );
  OA21X1 U9 ( .IN1(n13), .IN2(n14), .IN3(MODEROut[1]), .Q(r_TxEn) );
  OR4X1 U10 ( .IN1(r_TxBDNum[0]), .IN2(r_TxBDNum[1]), .IN3(r_TxBDNum[2]), 
        .IN4(r_TxBDNum[3]), .Q(n14) );
  OR4X1 U11 ( .IN1(r_TxBDNum[4]), .IN2(r_TxBDNum[5]), .IN3(r_TxBDNum[6]), 
        .IN4(r_TxBDNum[7]), .Q(n13) );
  NOR2X0 U12 ( .IN1(r_TxBDNum[7]), .IN2(n15), .QN(r_RxEn) );
  INVX0 U13 ( .INP(MODEROut[0]), .ZN(n15) );
  INVX0 U14 ( .INP(eth_top_test_point_11887_in), .ZN(n240) );
  OAI21X1 U15 ( .IN1(n30), .IN2(ResetTxCIrq_sync2), .IN3(n16), .QN(n249) );
  NAND3X0 U16 ( .IN1(TxCtrlEndFrm), .IN2(StartTxDone), .IN3(r_TxFlow), .QN(n16) );
  AO22X1 U17 ( .IN1(r_RxFlow), .IN2(SetPauseTimer), .IN3(n17), .IN4(
        SetRxCIrq_rxclk), .Q(n248) );
  NAND2X0 U18 ( .IN1(n33), .IN2(ResetRxCIrq_sync2), .QN(n17) );
  AO21X1 U19 ( .IN1(n6), .IN2(n18), .IN3(TxB_IRQ), .Q(n247) );
  NAND2X0 U20 ( .IN1(DataIn[0]), .IN2(n19), .QN(n18) );
  AO21X1 U21 ( .IN1(n3), .IN2(n20), .IN3(TxE_IRQ), .Q(n246) );
  NAND2X0 U22 ( .IN1(DataIn[1]), .IN2(n19), .QN(n20) );
  AO21X1 U23 ( .IN1(n5), .IN2(n21), .IN3(RxB_IRQ), .Q(n245) );
  NAND2X0 U24 ( .IN1(DataIn[2]), .IN2(n19), .QN(n21) );
  AO21X1 U25 ( .IN1(n22), .IN2(n2), .IN3(RxE_IRQ), .Q(n244) );
  NAND2X0 U26 ( .IN1(DataIn[3]), .IN2(n19), .QN(n22) );
  AO21X1 U27 ( .IN1(n23), .IN2(n1), .IN3(Busy_IRQ), .Q(n243) );
  NAND2X0 U28 ( .IN1(DataIn[4]), .IN2(n19), .QN(n23) );
  NAND2X0 U29 ( .IN1(n266), .IN2(n24), .QN(n242) );
  AO21X1 U30 ( .IN1(DataIn[5]), .IN2(n19), .IN3(n239), .Q(n24) );
  NAND2X0 U31 ( .IN1(n265), .IN2(n25), .QN(n241) );
  AO21X1 U32 ( .IN1(DataIn[6]), .IN2(n19), .IN3(n238), .Q(n25) );
  NOR2X0 U33 ( .IN1(n26), .IN2(n28), .QN(n19) );
  NAND3X0 U34 ( .IN1(n29), .IN2(n34), .IN3(n35), .QN(int_o) );
  AOI222X1 U35 ( .IN1(n27), .IN2(INT_MASKOut[6]), .IN3(n1), .IN4(
        INT_MASKOut[4]), .IN5(n4), .IN6(INT_MASKOut[5]), .QN(n35) );
  AOI22X1 U36 ( .IN1(n6), .IN2(INT_MASKOut[0]), .IN3(n3), .IN4(INT_MASKOut[1]), 
        .QN(n34) );
  AOI22X1 U37 ( .IN1(n5), .IN2(INT_MASKOut[2]), .IN3(n2), .IN4(INT_MASKOut[3]), 
        .QN(n29) );
  AND4X1 U38 ( .IN1(n36), .IN2(n37), .IN3(n38), .IN4(n39), .Q(
        \TX_BD_NUM_Wr[0] ) );
  NOR4X0 U39 ( .IN1(n40), .IN2(DataIn[27]), .IN3(DataIn[29]), .IN4(DataIn[28]), 
        .QN(n39) );
  OR4X1 U40 ( .IN1(DataIn[31]), .IN2(DataIn[30]), .IN3(DataIn[9]), .IN4(
        DataIn[8]), .Q(n40) );
  NOR4X0 U41 ( .IN1(n41), .IN2(DataIn[20]), .IN3(DataIn[22]), .IN4(DataIn[21]), 
        .QN(n38) );
  OR4X1 U42 ( .IN1(DataIn[24]), .IN2(DataIn[23]), .IN3(DataIn[26]), .IN4(
        DataIn[25]), .Q(n41) );
  NOR4X0 U43 ( .IN1(n42), .IN2(DataIn[13]), .IN3(DataIn[15]), .IN4(DataIn[14]), 
        .QN(n37) );
  OR4X1 U44 ( .IN1(DataIn[17]), .IN2(DataIn[16]), .IN3(DataIn[19]), .IN4(
        DataIn[18]), .Q(n42) );
  NOR4X0 U45 ( .IN1(n43), .IN2(DataIn[10]), .IN3(DataIn[12]), .IN4(DataIn[11]), 
        .QN(n36) );
  NAND3X0 U46 ( .IN1(n44), .IN2(n45), .IN3(n46), .QN(n43) );
  NAND2X0 U47 ( .IN1(DataIn[7]), .IN2(n47), .QN(n45) );
  OR4X1 U48 ( .IN1(DataIn[1]), .IN2(DataIn[2]), .IN3(DataIn[0]), .IN4(n48), 
        .Q(n47) );
  OR4X1 U49 ( .IN1(DataIn[6]), .IN2(DataIn[5]), .IN3(DataIn[4]), .IN4(
        DataIn[3]), .Q(n48) );
  NOR3X0 U50 ( .IN1(n49), .IN2(n50), .IN3(n51), .QN(TXCTRL_Wr[2]) );
  NOR2X0 U51 ( .IN1(n51), .IN2(n52), .QN(TXCTRL_Wr[1]) );
  NOR2X0 U52 ( .IN1(n53), .IN2(n51), .QN(TXCTRL_Wr[0]) );
  NOR2X0 U53 ( .IN1(n54), .IN2(n55), .QN(PACKETLEN_Wr[3]) );
  NOR2X0 U54 ( .IN1(n49), .IN2(n54), .QN(PACKETLEN_Wr[2]) );
  NOR2X0 U55 ( .IN1(n56), .IN2(n54), .QN(PACKETLEN_Wr[1]) );
  NOR2X0 U56 ( .IN1(n57), .IN2(n54), .QN(PACKETLEN_Wr[0]) );
  OR2X1 U57 ( .IN1(n58), .IN2(n59), .Q(n54) );
  NOR2X0 U58 ( .IN1(n32), .IN2(SetRxCIrq_sync3), .QN(N185) );
  NOR2X0 U59 ( .IN1(n31), .IN2(SetTxCIrq_sync3), .QN(N179) );
  NOR3X0 U60 ( .IN1(n49), .IN2(n28), .IN3(n60), .QN(MODER_Wr[2]) );
  NOR3X0 U61 ( .IN1(n56), .IN2(n28), .IN3(n60), .QN(MODER_Wr[1]) );
  NOR2X0 U62 ( .IN1(n28), .IN2(n61), .QN(MODER_Wr[0]) );
  NOR3X0 U63 ( .IN1(n62), .IN2(n63), .IN3(n56), .QN(MIITX_DATA_Wr[1]) );
  NOR2X0 U64 ( .IN1(n26), .IN2(n62), .QN(MIITX_DATA_Wr[0]) );
  NOR2X0 U65 ( .IN1(n52), .IN2(n64), .QN(MIIMODER_Wr[1]) );
  NOR2X0 U66 ( .IN1(n53), .IN2(n64), .QN(MIIMODER_Wr[0]) );
  INVX0 U67 ( .INP(n65), .ZN(n64) );
  AND2X1 U68 ( .IN1(n44), .IN2(n66), .Q(\MIICOMMAND_Wr[0] ) );
  INVX0 U69 ( .INP(n53), .ZN(n44) );
  NOR3X0 U70 ( .IN1(n62), .IN2(n60), .IN3(n56), .QN(MIIADDRESS_Wr[1]) );
  NOR2X0 U71 ( .IN1(n61), .IN2(n62), .QN(MIIADDRESS_Wr[0]) );
  NAND2X0 U72 ( .IN1(n67), .IN2(n68), .QN(n62) );
  NOR2X0 U73 ( .IN1(n52), .IN2(n69), .QN(MAC_ADDR1_Wr[1]) );
  OR2X1 U74 ( .IN1(n56), .IN2(n50), .Q(n52) );
  NOR2X0 U75 ( .IN1(n53), .IN2(n69), .QN(MAC_ADDR1_Wr[0]) );
  INVX0 U76 ( .INP(n70), .ZN(n69) );
  NAND2X0 U77 ( .IN1(n71), .IN2(n72), .QN(n53) );
  NOR2X0 U78 ( .IN1(n55), .IN2(n73), .QN(MAC_ADDR0_Wr[3]) );
  NOR2X0 U79 ( .IN1(n49), .IN2(n73), .QN(MAC_ADDR0_Wr[2]) );
  NOR2X0 U80 ( .IN1(n56), .IN2(n73), .QN(MAC_ADDR0_Wr[1]) );
  NOR2X0 U81 ( .IN1(n57), .IN2(n73), .QN(MAC_ADDR0_Wr[0]) );
  NOR3X0 U82 ( .IN1(n74), .IN2(n57), .IN3(n28), .QN(\IPGT_Wr[0] ) );
  NOR2X0 U83 ( .IN1(n26), .IN2(n58), .QN(\IPGR2_Wr[0] ) );
  NOR2X0 U84 ( .IN1(n58), .IN2(n61), .QN(\IPGR1_Wr[0] ) );
  NAND2X0 U85 ( .IN1(n75), .IN2(n72), .QN(n61) );
  NOR3X0 U86 ( .IN1(n59), .IN2(n57), .IN3(n28), .QN(\INT_MASK_Wr[0] ) );
  NAND2X0 U87 ( .IN1(n76), .IN2(n68), .QN(n28) );
  NOR2X0 U88 ( .IN1(n55), .IN2(n77), .QN(HASH1_Wr[3]) );
  NOR2X0 U89 ( .IN1(n49), .IN2(n77), .QN(HASH1_Wr[2]) );
  NOR2X0 U90 ( .IN1(n56), .IN2(n77), .QN(HASH1_Wr[1]) );
  NOR2X0 U91 ( .IN1(n57), .IN2(n77), .QN(HASH1_Wr[0]) );
  NOR2X0 U92 ( .IN1(n55), .IN2(n78), .QN(HASH0_Wr[3]) );
  NAND2X0 U93 ( .IN1(Cs[3]), .IN2(Rw), .QN(n55) );
  NOR2X0 U94 ( .IN1(n49), .IN2(n78), .QN(HASH0_Wr[2]) );
  NOR2X0 U95 ( .IN1(n56), .IN2(n78), .QN(HASH0_Wr[1]) );
  NAND2X0 U96 ( .IN1(Cs[1]), .IN2(Rw), .QN(n56) );
  NOR2X0 U97 ( .IN1(n57), .IN2(n78), .QN(HASH0_Wr[0]) );
  AO22X1 U98 ( .IN1(r_MaxFL[9]), .IN2(n79), .IN3(n80), .IN4(n81), .Q(
        DataOut[9]) );
  OR2X1 U99 ( .IN1(n82), .IN2(n83), .Q(n81) );
  AO221X1 U100 ( .IN1(r_HASH0[9]), .IN2(n84), .IN3(r_HASH1[9]), .IN4(n85), 
        .IN5(n86), .Q(n83) );
  AO22X1 U101 ( .IN1(r_TxPauseTV[9]), .IN2(n87), .IN3(r_MAC[9]), .IN4(n88), 
        .Q(n86) );
  AO221X1 U102 ( .IN1(MIIRX_DATAOut[9]), .IN2(n89), .IN3(r_ExDfrEn), .IN4(n90), 
        .IN5(n91), .Q(n82) );
  AO222X1 U103 ( .IN1(r_MAC[41]), .IN2(n70), .IN3(r_RGAD[1]), .IN4(n92), .IN5(
        r_CtrlData[9]), .IN6(n93), .Q(n91) );
  AO22X1 U104 ( .IN1(r_MaxFL[8]), .IN2(n79), .IN3(n80), .IN4(n94), .Q(
        DataOut[8]) );
  OR2X1 U105 ( .IN1(n95), .IN2(n96), .Q(n94) );
  AO221X1 U106 ( .IN1(r_MAC[8]), .IN2(n88), .IN3(r_TxPauseTV[8]), .IN4(n87), 
        .IN5(n97), .Q(n96) );
  AO222X1 U107 ( .IN1(r_HASH0[8]), .IN2(n84), .IN3(r_NoBckof), .IN4(n90), 
        .IN5(r_HASH1[8]), .IN6(n85), .Q(n97) );
  AO221X1 U108 ( .IN1(r_CtrlData[8]), .IN2(n93), .IN3(MIIRX_DATAOut[8]), .IN4(
        n89), .IN5(n98), .Q(n95) );
  AO222X1 U109 ( .IN1(r_MiiNoPre), .IN2(n65), .IN3(r_RGAD[0]), .IN4(n92), 
        .IN5(r_MAC[40]), .IN6(n70), .Q(n98) );
  AO22X1 U110 ( .IN1(r_MaxFL[7]), .IN2(n79), .IN3(n80), .IN4(n99), .Q(
        DataOut[7]) );
  OR2X1 U111 ( .IN1(n100), .IN2(n101), .Q(n99) );
  AO221X1 U112 ( .IN1(r_MAC[7]), .IN2(n88), .IN3(r_TxPauseTV[7]), .IN4(n87), 
        .IN5(n102), .Q(n101) );
  AO222X1 U113 ( .IN1(r_HASH0[7]), .IN2(n84), .IN3(r_LoopBck), .IN4(n90), 
        .IN5(r_HASH1[7]), .IN6(n85), .Q(n102) );
  AO221X1 U114 ( .IN1(r_CtrlData[7]), .IN2(n93), .IN3(MIIRX_DATAOut[7]), .IN4(
        n89), .IN5(n103), .Q(n100) );
  AO222X1 U115 ( .IN1(r_TxBDNum[7]), .IN2(n46), .IN3(r_ClkDiv[7]), .IN4(n65), 
        .IN5(r_MAC[39]), .IN6(n70), .Q(n103) );
  AO22X1 U116 ( .IN1(r_MaxFL[6]), .IN2(n79), .IN3(n80), .IN4(n104), .Q(
        DataOut[6]) );
  OR4X1 U117 ( .IN1(n105), .IN2(n106), .IN3(n107), .IN4(n108), .Q(n104) );
  AO221X1 U118 ( .IN1(r_TxBDNum[6]), .IN2(n46), .IN3(r_MAC[38]), .IN4(n70), 
        .IN5(n109), .Q(n108) );
  AO22X1 U119 ( .IN1(r_IPGR1[6]), .IN2(n110), .IN3(n111), .IN4(n27), .Q(n109)
         );
  AO221X1 U120 ( .IN1(r_ClkDiv[6]), .IN2(n65), .IN3(r_IPGT[6]), .IN4(n112), 
        .IN5(n113), .Q(n107) );
  AO22X1 U121 ( .IN1(n114), .IN2(INT_MASKOut[6]), .IN3(r_IPGR2[6]), .IN4(n115), 
        .Q(n113) );
  AO222X1 U122 ( .IN1(r_MAC[6]), .IN2(n88), .IN3(r_HASH1[6]), .IN4(n85), .IN5(
        r_TxPauseTV[6]), .IN6(n87), .Q(n106) );
  AO221X1 U123 ( .IN1(r_CtrlData[6]), .IN2(n93), .IN3(MIIRX_DATAOut[6]), .IN4(
        n89), .IN5(n116), .Q(n105) );
  AO22X1 U124 ( .IN1(r_HASH0[6]), .IN2(n84), .IN3(r_IFG), .IN4(n90), .Q(n116)
         );
  AO22X1 U125 ( .IN1(r_MaxFL[5]), .IN2(n79), .IN3(n80), .IN4(n117), .Q(
        DataOut[5]) );
  OR4X1 U126 ( .IN1(n118), .IN2(n119), .IN3(n120), .IN4(n121), .Q(n117) );
  AO221X1 U127 ( .IN1(r_TxBDNum[5]), .IN2(n46), .IN3(r_MAC[37]), .IN4(n70), 
        .IN5(n122), .Q(n121) );
  AO22X1 U128 ( .IN1(r_IPGR1[5]), .IN2(n110), .IN3(n111), .IN4(n4), .Q(n122)
         );
  AO221X1 U129 ( .IN1(r_ClkDiv[5]), .IN2(n65), .IN3(r_IPGT[5]), .IN4(n112), 
        .IN5(n123), .Q(n120) );
  AO22X1 U130 ( .IN1(n114), .IN2(INT_MASKOut[5]), .IN3(r_IPGR2[5]), .IN4(n115), 
        .Q(n123) );
  AO221X1 U131 ( .IN1(r_HASH0[5]), .IN2(n84), .IN3(r_HASH1[5]), .IN4(n85), 
        .IN5(n124), .Q(n119) );
  AO22X1 U132 ( .IN1(r_TxPauseTV[5]), .IN2(n87), .IN3(r_MAC[5]), .IN4(n88), 
        .Q(n124) );
  AO221X1 U133 ( .IN1(r_CollValid[5]), .IN2(n125), .IN3(r_CtrlData[5]), .IN4(
        n93), .IN5(n126), .Q(n118) );
  AO22X1 U134 ( .IN1(r_Pro), .IN2(n90), .IN3(MIIRX_DATAOut[5]), .IN4(n89), .Q(
        n126) );
  AO22X1 U135 ( .IN1(r_MaxFL[4]), .IN2(n79), .IN3(n80), .IN4(n127), .Q(
        DataOut[4]) );
  OR4X1 U136 ( .IN1(n128), .IN2(n129), .IN3(n130), .IN4(n131), .Q(n127) );
  AO221X1 U137 ( .IN1(r_TxBDNum[4]), .IN2(n46), .IN3(r_MAC[36]), .IN4(n70), 
        .IN5(n132), .Q(n131) );
  AO22X1 U138 ( .IN1(r_IPGR1[4]), .IN2(n110), .IN3(n111), .IN4(n1), .Q(n132)
         );
  AO221X1 U139 ( .IN1(r_IPGR2[4]), .IN2(n115), .IN3(n114), .IN4(INT_MASKOut[4]), .IN5(n133), .Q(n130) );
  AO222X1 U140 ( .IN1(r_ClkDiv[4]), .IN2(n65), .IN3(r_FIAD[4]), .IN4(n92), 
        .IN5(r_IPGT[4]), .IN6(n112), .Q(n133) );
  AO221X1 U141 ( .IN1(r_HASH0[4]), .IN2(n84), .IN3(r_HASH1[4]), .IN4(n85), 
        .IN5(n134), .Q(n129) );
  AO22X1 U142 ( .IN1(r_TxPauseTV[4]), .IN2(n87), .IN3(r_MAC[4]), .IN4(n88), 
        .Q(n134) );
  AO221X1 U143 ( .IN1(r_CollValid[4]), .IN2(n125), .IN3(r_CtrlData[4]), .IN4(
        n93), .IN5(n135), .Q(n128) );
  AO22X1 U144 ( .IN1(r_Iam), .IN2(n90), .IN3(MIIRX_DATAOut[4]), .IN4(n89), .Q(
        n135) );
  AO22X1 U145 ( .IN1(r_MaxFL[3]), .IN2(n79), .IN3(n80), .IN4(n136), .Q(
        DataOut[3]) );
  OR4X1 U146 ( .IN1(n137), .IN2(n138), .IN3(n139), .IN4(n140), .Q(n136) );
  AO221X1 U147 ( .IN1(r_TxBDNum[3]), .IN2(n46), .IN3(r_MAC[35]), .IN4(n70), 
        .IN5(n141), .Q(n140) );
  AO22X1 U148 ( .IN1(r_IPGR1[3]), .IN2(n110), .IN3(n111), .IN4(n2), .Q(n141)
         );
  AO221X1 U149 ( .IN1(r_IPGR2[3]), .IN2(n115), .IN3(n114), .IN4(INT_MASKOut[3]), .IN5(n142), .Q(n139) );
  AO222X1 U150 ( .IN1(r_ClkDiv[3]), .IN2(n65), .IN3(r_FIAD[3]), .IN4(n92), 
        .IN5(r_IPGT[3]), .IN6(n112), .Q(n142) );
  AO221X1 U151 ( .IN1(r_HASH0[3]), .IN2(n84), .IN3(r_HASH1[3]), .IN4(n85), 
        .IN5(n143), .Q(n138) );
  AO22X1 U152 ( .IN1(r_TxPauseTV[3]), .IN2(n87), .IN3(r_MAC[3]), .IN4(n88), 
        .Q(n143) );
  AO221X1 U153 ( .IN1(r_CollValid[3]), .IN2(n125), .IN3(r_CtrlData[3]), .IN4(
        n93), .IN5(n144), .Q(n137) );
  AO22X1 U154 ( .IN1(r_Bro), .IN2(n90), .IN3(MIIRX_DATAOut[3]), .IN4(n89), .Q(
        n144) );
  AO221X1 U155 ( .IN1(r_HASH1[31]), .IN2(n145), .IN3(r_MAC[31]), .IN4(n146), 
        .IN5(n147), .Q(DataOut[31]) );
  AO22X1 U156 ( .IN1(r_MinFL[15]), .IN2(n79), .IN3(r_HASH0[31]), .IN4(n148), 
        .Q(n147) );
  AO221X1 U157 ( .IN1(r_HASH1[30]), .IN2(n145), .IN3(r_MAC[30]), .IN4(n146), 
        .IN5(n149), .Q(DataOut[30]) );
  AO22X1 U158 ( .IN1(r_MinFL[14]), .IN2(n79), .IN3(r_HASH0[30]), .IN4(n148), 
        .Q(n149) );
  AO22X1 U159 ( .IN1(r_MaxFL[2]), .IN2(n79), .IN3(n80), .IN4(n150), .Q(
        DataOut[2]) );
  OR4X1 U160 ( .IN1(n151), .IN2(n152), .IN3(n153), .IN4(n154), .Q(n150) );
  AO221X1 U161 ( .IN1(n111), .IN2(n5), .IN3(r_IPGR1[2]), .IN4(n110), .IN5(n155), .Q(n154) );
  AO222X1 U162 ( .IN1(r_IPGR2[2]), .IN2(n115), .IN3(r_IPGT[2]), .IN4(n112), 
        .IN5(n114), .IN6(INT_MASKOut[2]), .Q(n155) );
  AO221X1 U163 ( .IN1(r_FIAD[2]), .IN2(n92), .IN3(r_ClkDiv[2]), .IN4(n65), 
        .IN5(n156), .Q(n153) );
  AO222X1 U164 ( .IN1(r_WCtrlData), .IN2(n66), .IN3(NValid_stat), .IN4(n157), 
        .IN5(n158), .IN6(r_TxFlow), .Q(n156) );
  AO221X1 U165 ( .IN1(r_MAC[2]), .IN2(n88), .IN3(r_TxPauseTV[2]), .IN4(n87), 
        .IN5(n159), .Q(n152) );
  AO222X1 U166 ( .IN1(r_HASH0[2]), .IN2(n84), .IN3(r_NoPre), .IN4(n90), .IN5(
        r_HASH1[2]), .IN6(n85), .Q(n159) );
  AO221X1 U167 ( .IN1(r_CtrlData[2]), .IN2(n93), .IN3(MIIRX_DATAOut[2]), .IN4(
        n89), .IN5(n160), .Q(n151) );
  AO222X1 U168 ( .IN1(r_MAC[34]), .IN2(n70), .IN3(r_TxBDNum[2]), .IN4(n46), 
        .IN5(r_CollValid[2]), .IN6(n125), .Q(n160) );
  AO221X1 U169 ( .IN1(r_HASH1[29]), .IN2(n145), .IN3(r_MAC[29]), .IN4(n146), 
        .IN5(n161), .Q(DataOut[29]) );
  AO22X1 U170 ( .IN1(r_MinFL[13]), .IN2(n79), .IN3(r_HASH0[29]), .IN4(n148), 
        .Q(n161) );
  AO221X1 U171 ( .IN1(r_HASH1[28]), .IN2(n145), .IN3(r_MAC[28]), .IN4(n146), 
        .IN5(n162), .Q(DataOut[28]) );
  AO22X1 U172 ( .IN1(r_MinFL[12]), .IN2(n79), .IN3(r_HASH0[28]), .IN4(n148), 
        .Q(n162) );
  AO221X1 U173 ( .IN1(r_HASH1[27]), .IN2(n145), .IN3(r_MAC[27]), .IN4(n146), 
        .IN5(n163), .Q(DataOut[27]) );
  AO22X1 U174 ( .IN1(r_MinFL[11]), .IN2(n79), .IN3(r_HASH0[27]), .IN4(n148), 
        .Q(n163) );
  AO221X1 U175 ( .IN1(r_HASH1[26]), .IN2(n145), .IN3(r_MAC[26]), .IN4(n146), 
        .IN5(n164), .Q(DataOut[26]) );
  AO22X1 U176 ( .IN1(r_MinFL[10]), .IN2(n79), .IN3(r_HASH0[26]), .IN4(n148), 
        .Q(n164) );
  AO221X1 U177 ( .IN1(r_HASH1[25]), .IN2(n145), .IN3(r_MAC[25]), .IN4(n146), 
        .IN5(n165), .Q(DataOut[25]) );
  AO22X1 U178 ( .IN1(r_MinFL[9]), .IN2(n79), .IN3(r_HASH0[25]), .IN4(n148), 
        .Q(n165) );
  AO221X1 U179 ( .IN1(r_HASH1[24]), .IN2(n145), .IN3(r_MAC[24]), .IN4(n146), 
        .IN5(n166), .Q(DataOut[24]) );
  AO22X1 U180 ( .IN1(r_MinFL[8]), .IN2(n79), .IN3(r_HASH0[24]), .IN4(n148), 
        .Q(n166) );
  AO221X1 U181 ( .IN1(r_HASH1[23]), .IN2(n145), .IN3(r_MAC[23]), .IN4(n146), 
        .IN5(n167), .Q(DataOut[23]) );
  AO22X1 U182 ( .IN1(r_MinFL[7]), .IN2(n79), .IN3(r_HASH0[23]), .IN4(n148), 
        .Q(n167) );
  AO221X1 U183 ( .IN1(r_HASH1[22]), .IN2(n145), .IN3(r_MAC[22]), .IN4(n146), 
        .IN5(n168), .Q(DataOut[22]) );
  AO22X1 U184 ( .IN1(r_MinFL[6]), .IN2(n79), .IN3(r_HASH0[22]), .IN4(n148), 
        .Q(n168) );
  AO221X1 U185 ( .IN1(r_HASH1[21]), .IN2(n145), .IN3(r_MAC[21]), .IN4(n146), 
        .IN5(n169), .Q(DataOut[21]) );
  AO22X1 U186 ( .IN1(r_MinFL[5]), .IN2(n79), .IN3(r_HASH0[21]), .IN4(n148), 
        .Q(n169) );
  AO221X1 U187 ( .IN1(r_HASH1[20]), .IN2(n145), .IN3(r_MAC[20]), .IN4(n146), 
        .IN5(n170), .Q(DataOut[20]) );
  AO22X1 U188 ( .IN1(r_MinFL[4]), .IN2(n79), .IN3(r_HASH0[20]), .IN4(n148), 
        .Q(n170) );
  AO22X1 U189 ( .IN1(r_MaxFL[1]), .IN2(n79), .IN3(n80), .IN4(n171), .Q(
        DataOut[1]) );
  OR4X1 U190 ( .IN1(n172), .IN2(n173), .IN3(n174), .IN4(n175), .Q(n171) );
  AO221X1 U191 ( .IN1(n111), .IN2(n3), .IN3(r_IPGR1[1]), .IN4(n110), .IN5(n176), .Q(n175) );
  AO222X1 U192 ( .IN1(r_IPGR2[1]), .IN2(n115), .IN3(r_IPGT[1]), .IN4(n112), 
        .IN5(n114), .IN6(INT_MASKOut[1]), .Q(n176) );
  AO221X1 U193 ( .IN1(r_FIAD[1]), .IN2(n92), .IN3(r_ClkDiv[1]), .IN4(n65), 
        .IN5(n177), .Q(n174) );
  AO222X1 U194 ( .IN1(r_RStat), .IN2(n66), .IN3(Busy_stat), .IN4(n157), .IN5(
        n158), .IN6(r_RxFlow), .Q(n177) );
  AO221X1 U195 ( .IN1(r_MAC[1]), .IN2(n88), .IN3(r_TxPauseTV[1]), .IN4(n87), 
        .IN5(n178), .Q(n173) );
  AO222X1 U196 ( .IN1(r_HASH0[1]), .IN2(n84), .IN3(n90), .IN4(MODEROut[1]), 
        .IN5(r_HASH1[1]), .IN6(n85), .Q(n178) );
  AO221X1 U197 ( .IN1(r_CtrlData[1]), .IN2(n93), .IN3(MIIRX_DATAOut[1]), .IN4(
        n89), .IN5(n179), .Q(n172) );
  AO222X1 U198 ( .IN1(r_MAC[33]), .IN2(n70), .IN3(r_TxBDNum[1]), .IN4(n46), 
        .IN5(r_CollValid[1]), .IN6(n125), .Q(n179) );
  AO221X1 U199 ( .IN1(r_HASH0[19]), .IN2(n148), .IN3(r_MinFL[3]), .IN4(n79), 
        .IN5(n180), .Q(DataOut[19]) );
  AO222X1 U200 ( .IN1(r_HASH1[19]), .IN2(n145), .IN3(r_MaxRet[3]), .IN4(n181), 
        .IN5(r_MAC[19]), .IN6(n146), .Q(n180) );
  AO221X1 U201 ( .IN1(r_HASH0[18]), .IN2(n148), .IN3(r_MinFL[2]), .IN4(n79), 
        .IN5(n182), .Q(DataOut[18]) );
  AO222X1 U202 ( .IN1(r_HASH1[18]), .IN2(n145), .IN3(r_MaxRet[2]), .IN4(n181), 
        .IN5(r_MAC[18]), .IN6(n146), .Q(n182) );
  AO221X1 U203 ( .IN1(r_HASH0[17]), .IN2(n148), .IN3(r_MinFL[1]), .IN4(n79), 
        .IN5(n183), .Q(DataOut[17]) );
  AO222X1 U204 ( .IN1(r_HASH1[17]), .IN2(n145), .IN3(r_MaxRet[1]), .IN4(n181), 
        .IN5(r_MAC[17]), .IN6(n146), .Q(n183) );
  AND2X1 U205 ( .IN1(n125), .IN2(n80), .Q(n181) );
  AO221X1 U206 ( .IN1(r_HASH0[16]), .IN2(n148), .IN3(r_MinFL[0]), .IN4(n79), 
        .IN5(n184), .Q(DataOut[16]) );
  AO222X1 U207 ( .IN1(r_HASH1[16]), .IN2(n145), .IN3(n80), .IN4(n185), .IN5(
        r_MAC[16]), .IN6(n146), .Q(n184) );
  NOR2X0 U208 ( .IN1(n186), .IN2(n73), .QN(n146) );
  NAND2X0 U209 ( .IN1(n88), .IN2(n71), .QN(n73) );
  AO222X1 U210 ( .IN1(r_RecSmall), .IN2(n90), .IN3(r_MaxRet[0]), .IN4(n125), 
        .IN5(r_TxPauseRq), .IN6(n87), .Q(n185) );
  NOR2X0 U211 ( .IN1(n186), .IN2(n77), .QN(n145) );
  NAND2X0 U212 ( .IN1(n85), .IN2(n71), .QN(n77) );
  NOR2X0 U213 ( .IN1(n186), .IN2(n78), .QN(n148) );
  NAND2X0 U214 ( .IN1(n84), .IN2(n71), .QN(n78) );
  AO22X1 U215 ( .IN1(r_MaxFL[15]), .IN2(n79), .IN3(n80), .IN4(n187), .Q(
        DataOut[15]) );
  OR2X1 U216 ( .IN1(n188), .IN2(n189), .Q(n187) );
  AO221X1 U217 ( .IN1(r_HASH0[15]), .IN2(n84), .IN3(r_HASH1[15]), .IN4(n85), 
        .IN5(n190), .Q(n189) );
  AO22X1 U218 ( .IN1(r_TxPauseTV[15]), .IN2(n87), .IN3(r_MAC[15]), .IN4(n88), 
        .Q(n190) );
  AO221X1 U219 ( .IN1(r_MAC[47]), .IN2(n70), .IN3(r_CtrlData[15]), .IN4(n93), 
        .IN5(n191), .Q(n188) );
  AO22X1 U220 ( .IN1(r_Pad), .IN2(n90), .IN3(MIIRX_DATAOut[15]), .IN4(n89), 
        .Q(n191) );
  AO22X1 U221 ( .IN1(r_MaxFL[14]), .IN2(n79), .IN3(n80), .IN4(n192), .Q(
        DataOut[14]) );
  OR2X1 U222 ( .IN1(n193), .IN2(n194), .Q(n192) );
  AO221X1 U223 ( .IN1(r_HASH0[14]), .IN2(n84), .IN3(r_HASH1[14]), .IN4(n85), 
        .IN5(n195), .Q(n194) );
  AO22X1 U224 ( .IN1(r_TxPauseTV[14]), .IN2(n87), .IN3(r_MAC[14]), .IN4(n88), 
        .Q(n195) );
  AO221X1 U225 ( .IN1(r_MAC[46]), .IN2(n70), .IN3(r_CtrlData[14]), .IN4(n93), 
        .IN5(n196), .Q(n193) );
  AO22X1 U226 ( .IN1(r_HugEn), .IN2(n90), .IN3(MIIRX_DATAOut[14]), .IN4(n89), 
        .Q(n196) );
  AO22X1 U227 ( .IN1(r_MaxFL[13]), .IN2(n79), .IN3(n80), .IN4(n197), .Q(
        DataOut[13]) );
  OR2X1 U228 ( .IN1(n198), .IN2(n199), .Q(n197) );
  AO221X1 U229 ( .IN1(r_HASH0[13]), .IN2(n84), .IN3(r_HASH1[13]), .IN4(n85), 
        .IN5(n200), .Q(n199) );
  AO22X1 U230 ( .IN1(r_TxPauseTV[13]), .IN2(n87), .IN3(r_MAC[13]), .IN4(n88), 
        .Q(n200) );
  AO221X1 U231 ( .IN1(r_MAC[45]), .IN2(n70), .IN3(r_CtrlData[13]), .IN4(n93), 
        .IN5(n201), .Q(n198) );
  AO22X1 U232 ( .IN1(r_CrcEn), .IN2(n90), .IN3(MIIRX_DATAOut[13]), .IN4(n89), 
        .Q(n201) );
  AO22X1 U233 ( .IN1(r_MaxFL[12]), .IN2(n79), .IN3(n80), .IN4(n202), .Q(
        DataOut[12]) );
  OR2X1 U234 ( .IN1(n203), .IN2(n204), .Q(n202) );
  AO221X1 U235 ( .IN1(r_HASH0[12]), .IN2(n84), .IN3(r_HASH1[12]), .IN4(n85), 
        .IN5(n205), .Q(n204) );
  AO22X1 U236 ( .IN1(r_TxPauseTV[12]), .IN2(n87), .IN3(r_MAC[12]), .IN4(n88), 
        .Q(n205) );
  AO221X1 U237 ( .IN1(MIIRX_DATAOut[12]), .IN2(n89), .IN3(r_DlyCrcEn), .IN4(
        n90), .IN5(n206), .Q(n203) );
  AO222X1 U238 ( .IN1(r_MAC[44]), .IN2(n70), .IN3(r_RGAD[4]), .IN4(n92), .IN5(
        r_CtrlData[12]), .IN6(n93), .Q(n206) );
  AO22X1 U239 ( .IN1(r_MaxFL[11]), .IN2(n79), .IN3(n80), .IN4(n207), .Q(
        DataOut[11]) );
  OR2X1 U240 ( .IN1(n208), .IN2(n209), .Q(n207) );
  AO221X1 U241 ( .IN1(r_HASH0[11]), .IN2(n84), .IN3(r_HASH1[11]), .IN4(n85), 
        .IN5(n210), .Q(n209) );
  AO22X1 U242 ( .IN1(r_TxPauseTV[11]), .IN2(n87), .IN3(r_MAC[11]), .IN4(n88), 
        .Q(n210) );
  AO221X1 U243 ( .IN1(MIIRX_DATAOut[11]), .IN2(n89), .IN3(MODEROut_11), .IN4(
        n90), .IN5(n211), .Q(n208) );
  AO222X1 U244 ( .IN1(r_MAC[43]), .IN2(n70), .IN3(r_RGAD[3]), .IN4(n92), .IN5(
        r_CtrlData[11]), .IN6(n93), .Q(n211) );
  AO22X1 U245 ( .IN1(r_MaxFL[10]), .IN2(n79), .IN3(n80), .IN4(n212), .Q(
        DataOut[10]) );
  OR2X1 U246 ( .IN1(n213), .IN2(n214), .Q(n212) );
  AO221X1 U247 ( .IN1(r_HASH0[10]), .IN2(n84), .IN3(r_HASH1[10]), .IN4(n85), 
        .IN5(n215), .Q(n214) );
  AO22X1 U248 ( .IN1(r_TxPauseTV[10]), .IN2(n87), .IN3(r_MAC[10]), .IN4(n88), 
        .Q(n215) );
  AO221X1 U249 ( .IN1(MIIRX_DATAOut[10]), .IN2(n89), .IN3(r_FullD), .IN4(n90), 
        .IN5(n216), .Q(n213) );
  AO222X1 U250 ( .IN1(r_MAC[42]), .IN2(n70), .IN3(r_RGAD[2]), .IN4(n92), .IN5(
        r_CtrlData[10]), .IN6(n93), .Q(n216) );
  AO22X1 U251 ( .IN1(r_MaxFL[0]), .IN2(n79), .IN3(n80), .IN4(n217), .Q(
        DataOut[0]) );
  OR4X1 U252 ( .IN1(n218), .IN2(n219), .IN3(n220), .IN4(n221), .Q(n217) );
  AO221X1 U253 ( .IN1(n111), .IN2(n6), .IN3(r_IPGR1[0]), .IN4(n110), .IN5(n222), .Q(n221) );
  AO222X1 U254 ( .IN1(r_IPGR2[0]), .IN2(n115), .IN3(r_IPGT[0]), .IN4(n112), 
        .IN5(n114), .IN6(INT_MASKOut[0]), .Q(n222) );
  AND2X1 U255 ( .IN1(n223), .IN2(n76), .Q(n114) );
  AND2X1 U256 ( .IN1(n224), .IN2(n76), .Q(n112) );
  AND2X1 U257 ( .IN1(n225), .IN2(n226), .Q(n115) );
  AND2X1 U258 ( .IN1(n227), .IN2(n226), .Q(n110) );
  AND2X1 U259 ( .IN1(n225), .IN2(n76), .Q(n111) );
  AO221X1 U260 ( .IN1(r_FIAD[0]), .IN2(n92), .IN3(r_ClkDiv[0]), .IN4(n65), 
        .IN5(n228), .Q(n220) );
  AO222X1 U261 ( .IN1(r_ScanStat), .IN2(n66), .IN3(LinkFail), .IN4(n157), 
        .IN5(r_PassAll), .IN6(n158), .Q(n228) );
  AND3X1 U262 ( .IN1(Address[3]), .IN2(n229), .IN3(n225), .Q(n158) );
  AND2X1 U263 ( .IN1(n224), .IN2(n67), .Q(n157) );
  NOR2X0 U264 ( .IN1(n74), .IN2(n230), .QN(n66) );
  NOR2X0 U265 ( .IN1(n59), .IN2(n230), .QN(n65) );
  AND2X1 U266 ( .IN1(n227), .IN2(n67), .Q(n92) );
  AO221X1 U267 ( .IN1(r_MAC[0]), .IN2(n88), .IN3(r_TxPauseTV[0]), .IN4(n87), 
        .IN5(n231), .Q(n219) );
  AO222X1 U268 ( .IN1(r_HASH0[0]), .IN2(n84), .IN3(n90), .IN4(MODEROut[0]), 
        .IN5(r_HASH1[0]), .IN6(n85), .Q(n231) );
  NOR2X0 U269 ( .IN1(n232), .IN2(n74), .QN(n85) );
  AND2X1 U270 ( .IN1(n227), .IN2(n76), .Q(n90) );
  NOR2X0 U271 ( .IN1(n60), .IN2(Address[4]), .QN(n227) );
  NOR2X0 U272 ( .IN1(n232), .IN2(n59), .QN(n84) );
  INVX0 U273 ( .INP(n51), .ZN(n87) );
  NAND3X0 U274 ( .IN1(n226), .IN2(n75), .IN3(Address[4]), .QN(n51) );
  NOR2X0 U275 ( .IN1(n232), .IN2(n60), .QN(n88) );
  AO221X1 U276 ( .IN1(r_CtrlData[0]), .IN2(n93), .IN3(MIIRX_DATAOut[0]), .IN4(
        n89), .IN5(n233), .Q(n218) );
  AO222X1 U277 ( .IN1(r_MAC[32]), .IN2(n70), .IN3(r_TxBDNum[0]), .IN4(n46), 
        .IN5(r_CollValid[0]), .IN6(n125), .Q(n233) );
  AND2X1 U278 ( .IN1(n224), .IN2(n226), .Q(n125) );
  NOR2X0 U279 ( .IN1(n74), .IN2(Address[4]), .QN(n224) );
  NOR2X0 U280 ( .IN1(n60), .IN2(n230), .QN(n46) );
  INVX0 U281 ( .INP(n75), .ZN(n60) );
  NOR2X0 U282 ( .IN1(Address[0]), .IN2(Address[1]), .QN(n75) );
  NOR2X0 U283 ( .IN1(n232), .IN2(n63), .QN(n70) );
  NAND2X0 U284 ( .IN1(Address[4]), .IN2(n76), .QN(n232) );
  NOR2X0 U285 ( .IN1(Address[2]), .IN2(Address[3]), .QN(n76) );
  AND2X1 U286 ( .IN1(n223), .IN2(n67), .Q(n89) );
  AND2X1 U287 ( .IN1(n225), .IN2(n67), .Q(n93) );
  NOR2X0 U288 ( .IN1(n229), .IN2(n234), .QN(n67) );
  NOR2X0 U289 ( .IN1(n63), .IN2(Address[4]), .QN(n225) );
  INVX0 U290 ( .INP(n235), .ZN(n63) );
  AND3X1 U291 ( .IN1(n223), .IN2(n226), .IN3(n80), .Q(n79) );
  NOR2X0 U292 ( .IN1(n186), .IN2(n50), .QN(n80) );
  OR2X1 U293 ( .IN1(Rw), .IN2(n236), .Q(n186) );
  NOR4X0 U294 ( .IN1(Cs[0]), .IN2(Cs[1]), .IN3(Cs[2]), .IN4(Cs[3]), .QN(n236)
         );
  NOR2X0 U295 ( .IN1(n59), .IN2(Address[4]), .QN(n223) );
  NAND2X0 U296 ( .IN1(Address[1]), .IN2(n237), .QN(n59) );
  NOR3X0 U297 ( .IN1(n26), .IN2(n50), .IN3(n230), .QN(\CTRLMODER_Wr[0] ) );
  OR3X1 U298 ( .IN1(Address[2]), .IN2(Address[4]), .IN3(n234), .Q(n230) );
  INVX0 U299 ( .INP(Address[3]), .ZN(n234) );
  NAND2X0 U300 ( .IN1(n235), .IN2(n72), .QN(n26) );
  INVX0 U301 ( .INP(n57), .ZN(n72) );
  NOR2X0 U302 ( .IN1(n237), .IN2(Address[1]), .QN(n235) );
  INVX0 U303 ( .INP(Address[0]), .ZN(n237) );
  NOR3X0 U304 ( .IN1(n74), .IN2(n57), .IN3(n58), .QN(COLLCONF_Wr_0) );
  NAND2X0 U305 ( .IN1(Rw), .IN2(Cs[0]), .QN(n57) );
  NOR3X0 U306 ( .IN1(n74), .IN2(n49), .IN3(n58), .QN(\COLLCONF_Wr[2] ) );
  NAND2X0 U307 ( .IN1(n226), .IN2(n68), .QN(n58) );
  NOR2X0 U308 ( .IN1(n50), .IN2(Address[4]), .QN(n68) );
  INVX0 U309 ( .INP(n71), .ZN(n50) );
  NOR3X0 U310 ( .IN1(Address[7]), .IN2(Address[6]), .IN3(Address[5]), .QN(n71)
         );
  NOR2X0 U311 ( .IN1(n229), .IN2(Address[3]), .QN(n226) );
  INVX0 U312 ( .INP(Address[2]), .ZN(n229) );
  NAND2X0 U313 ( .IN1(Cs[2]), .IN2(Rw), .QN(n49) );
  NAND2X0 U314 ( .IN1(Address[1]), .IN2(Address[0]), .QN(n74) );
endmodule


module eth_receivecontrol_DW01_dec_0 ( A, SUM );
  input [15:0] A;
  output [15:0] SUM;
  wire   n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42;

  AO21X1 U15 ( .IN1(A[9]), .IN2(n35), .IN3(n15), .Q(SUM[9]) );
  AO21X1 U16 ( .IN1(A[8]), .IN2(n36), .IN3(n16), .Q(SUM[8]) );
  AO21X1 U17 ( .IN1(A[7]), .IN2(n37), .IN3(n17), .Q(SUM[7]) );
  AO21X1 U18 ( .IN1(A[6]), .IN2(n38), .IN3(n18), .Q(SUM[6]) );
  AO21X1 U19 ( .IN1(A[5]), .IN2(n39), .IN3(n19), .Q(SUM[5]) );
  AO21X1 U20 ( .IN1(A[4]), .IN2(n40), .IN3(n20), .Q(SUM[4]) );
  AO21X1 U21 ( .IN1(A[3]), .IN2(n41), .IN3(n21), .Q(SUM[3]) );
  AO21X1 U22 ( .IN1(A[2]), .IN2(n42), .IN3(n22), .Q(SUM[2]) );
  AO21X1 U23 ( .IN1(A[1]), .IN2(A[0]), .IN3(n23), .Q(SUM[1]) );
  XOR2X1 U24 ( .IN1(A[15]), .IN2(n24), .Q(SUM[15]) );
  XNOR2X1 U26 ( .IN1(A[14]), .IN2(n30), .Q(SUM[14]) );
  AO21X1 U27 ( .IN1(A[13]), .IN2(n31), .IN3(n25), .Q(SUM[13]) );
  AO21X1 U29 ( .IN1(A[12]), .IN2(n32), .IN3(n26), .Q(SUM[12]) );
  AO21X1 U31 ( .IN1(A[11]), .IN2(n33), .IN3(n27), .Q(SUM[11]) );
  AO21X1 U33 ( .IN1(A[10]), .IN2(n34), .IN3(n28), .Q(SUM[10]) );
  INVX0 U1 ( .INP(n25), .ZN(n30) );
  INVX0 U2 ( .INP(n23), .ZN(n42) );
  INVX0 U3 ( .INP(n27), .ZN(n32) );
  INVX0 U4 ( .INP(n26), .ZN(n31) );
  INVX0 U5 ( .INP(n22), .ZN(n41) );
  INVX0 U6 ( .INP(n21), .ZN(n40) );
  INVX0 U7 ( .INP(n20), .ZN(n39) );
  INVX0 U8 ( .INP(n19), .ZN(n38) );
  INVX0 U9 ( .INP(n18), .ZN(n37) );
  INVX0 U10 ( .INP(n17), .ZN(n36) );
  INVX0 U11 ( .INP(n16), .ZN(n35) );
  INVX0 U12 ( .INP(n15), .ZN(n34) );
  INVX0 U13 ( .INP(n28), .ZN(n33) );
  NOR2X0 U14 ( .IN1(A[1]), .IN2(A[0]), .QN(n23) );
  NOR2X0 U25 ( .IN1(A[14]), .IN2(n30), .QN(n24) );
  INVX0 U28 ( .INP(A[0]), .ZN(SUM[0]) );
  NOR2X0 U30 ( .IN1(n33), .IN2(A[11]), .QN(n27) );
  NOR2X0 U32 ( .IN1(n32), .IN2(A[12]), .QN(n26) );
  NOR2X0 U34 ( .IN1(n31), .IN2(A[13]), .QN(n25) );
  NOR2X0 U35 ( .IN1(n42), .IN2(A[2]), .QN(n22) );
  NOR2X0 U36 ( .IN1(n41), .IN2(A[3]), .QN(n21) );
  NOR2X0 U37 ( .IN1(n40), .IN2(A[4]), .QN(n20) );
  NOR2X0 U38 ( .IN1(n39), .IN2(A[5]), .QN(n19) );
  NOR2X0 U39 ( .IN1(n38), .IN2(A[6]), .QN(n18) );
  NOR2X0 U40 ( .IN1(n37), .IN2(A[7]), .QN(n17) );
  NOR2X0 U41 ( .IN1(n36), .IN2(A[8]), .QN(n16) );
  NOR2X0 U42 ( .IN1(n35), .IN2(A[9]), .QN(n15) );
  NOR2X0 U43 ( .IN1(n34), .IN2(A[10]), .QN(n28) );
endmodule


module eth_receivecontrol_test_1 ( MTxClk, MRxClk, TxReset, RxReset, RxData, 
        RxValid, RxStartFrm, RxEndFrm, RxFlow, ReceiveEnd, MAC, DlyCrcEn, 
        TxDoneIn, TxAbortIn, TxStartFrmOut, ReceivedLengthOK, 
        ReceivedPacketGood, TxUsedDataOutDetected, Pause, ReceivedPauseFrm, 
        AddressOK, RxStatusWriteLatched_sync2, r_PassAll, SetPauseTimer, 
        eth_top_data_sourcea_in, eth_top_test_mode_in, 
        eth_top_test_point_11887_in, test_so, test_se );
  input [7:0] RxData;
  input [47:0] MAC;
  input MTxClk, MRxClk, TxReset, RxReset, RxValid, RxStartFrm, RxEndFrm,
         RxFlow, ReceiveEnd, DlyCrcEn, TxDoneIn, TxAbortIn, TxStartFrmOut,
         ReceivedLengthOK, ReceivedPacketGood, TxUsedDataOutDetected,
         RxStatusWriteLatched_sync2, r_PassAll, eth_top_data_sourcea_in,
         eth_top_test_mode_in, eth_top_test_point_11887_in, test_se;
  output Pause, ReceivedPauseFrm, AddressOK, SetPauseTimer, test_so;
  wire   N143, N144, N145, N146, N147, N148, N149, N150, N151, N152, N153,
         N154, N155, N156, N157, N158, PauseTimerEq0_sync1, N183, n195, n212,
         n213, n214, n216, n218, n220, n222, n224, n226, n228, n230, n232,
         n234, n236, n238, n240, n242, n244, n246, n247, n248, n249, n250,
         n260, n333, n334, n336, n337, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n1, n2, n3, n4, n5,
         n6, n7, n8, n152, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n198, n199,
         n200, n201, n202, n203, n204, n205, n211, n297, n314, n332, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n153, n193, n194, n196, n197, n206, n207, n208, n209, n210,
         n215, n217, n219, n223;
  wire   [15:0] PauseTimer;
  assign test_so = n187;

  SDFFARX1 \DlyCrcCnt_reg[0]  ( .D(n406), .SI(n154), .SE(test_se), .CLK(n9), 
        .RSTB(n211), .Q(n191), .QN(n6) );
  SDFFARX1 \DlyCrcCnt_reg[2]  ( .D(n405), .SI(n190), .SE(test_se), .CLK(n9), 
        .RSTB(n211), .Q(n189), .QN(n8) );
  SDFFARX1 \DlyCrcCnt_reg[1]  ( .D(n404), .SI(n191), .SE(test_se), .CLK(n9), 
        .RSTB(n211), .Q(n190), .QN(n297) );
  SDFFARX1 \ByteCnt_reg[0]  ( .D(n403), .SI(n178), .SE(test_se), .CLK(n11), 
        .RSTB(n211), .Q(n3), .QN(n336) );
  SDFFASX1 DetectionWindow_reg ( .D(n401), .SI(n205), .SE(test_se), .CLK(n9), 
        .SETB(n211), .Q(n188), .QN(n314) );
  SDFFARX1 \ByteCnt_reg[4]  ( .D(n402), .SI(n2), .SE(test_se), .CLK(n9), 
        .RSTB(n211), .Q(n205), .QN(n219) );
  SDFFARX1 \ByteCnt_reg[1]  ( .D(n400), .SI(n3), .SE(test_se), .CLK(n11), 
        .RSTB(n211), .Q(n4), .QN(n217) );
  SDFFARX1 \ByteCnt_reg[2]  ( .D(n399), .SI(n4), .SE(test_se), .CLK(n11), 
        .RSTB(n211), .Q(n1), .QN(n334) );
  SDFFARX1 \ByteCnt_reg[3]  ( .D(n398), .SI(n1), .SE(test_se), .CLK(n11), 
        .RSTB(n211), .Q(n2), .QN(n333) );
  SDFFARX1 \AssembledTimerValue_reg[7]  ( .D(n386), .SI(n185), .SE(test_se), 
        .CLK(n10), .RSTB(n211), .Q(n186) );
  SDFFARX1 \AssembledTimerValue_reg[6]  ( .D(n387), .SI(n184), .SE(test_se), 
        .CLK(n10), .RSTB(n211), .Q(n185) );
  SDFFARX1 \AssembledTimerValue_reg[5]  ( .D(n388), .SI(n183), .SE(test_se), 
        .CLK(n11), .RSTB(n211), .Q(n184) );
  SDFFARX1 \AssembledTimerValue_reg[4]  ( .D(n389), .SI(n182), .SE(test_se), 
        .CLK(n10), .RSTB(n211), .Q(n183) );
  SDFFARX1 \AssembledTimerValue_reg[3]  ( .D(n390), .SI(n181), .SE(test_se), 
        .CLK(n10), .RSTB(n211), .Q(n182) );
  SDFFARX1 \AssembledTimerValue_reg[2]  ( .D(n391), .SI(n180), .SE(test_se), 
        .CLK(n10), .RSTB(n211), .Q(n181) );
  SDFFARX1 \AssembledTimerValue_reg[1]  ( .D(n392), .SI(n179), .SE(test_se), 
        .CLK(n10), .RSTB(n211), .Q(n180) );
  SDFFARX1 \AssembledTimerValue_reg[0]  ( .D(n393), .SI(AddressOK), .SE(
        test_se), .CLK(n10), .RSTB(n211), .Q(n179) );
  SDFFARX1 TypeLengthOK_reg ( .D(n396), .SI(n198), .SE(test_se), .CLK(n9), 
        .RSTB(n211), .Q(n187), .QN(n5) );
  SDFFARX1 OpCodeOK_reg ( .D(n397), .SI(n170), .SE(test_se), .CLK(n13), .RSTB(
        n211), .Q(n204), .QN(n215) );
  SDFFARX1 \AssembledTimerValue_reg[15]  ( .D(n378), .SI(n177), .SE(test_se), 
        .CLK(n11), .RSTB(n211), .Q(n178) );
  SDFFARX1 \AssembledTimerValue_reg[14]  ( .D(n379), .SI(n176), .SE(test_se), 
        .CLK(n11), .RSTB(n211), .Q(n177) );
  SDFFARX1 \AssembledTimerValue_reg[13]  ( .D(n380), .SI(n175), .SE(test_se), 
        .CLK(n11), .RSTB(n211), .Q(n176) );
  SDFFARX1 \AssembledTimerValue_reg[12]  ( .D(n381), .SI(n174), .SE(test_se), 
        .CLK(n10), .RSTB(n211), .Q(n175) );
  SDFFARX1 \AssembledTimerValue_reg[11]  ( .D(n382), .SI(n173), .SE(test_se), 
        .CLK(n10), .RSTB(n211), .Q(n174) );
  SDFFARX1 \AssembledTimerValue_reg[10]  ( .D(n383), .SI(n172), .SE(test_se), 
        .CLK(n10), .RSTB(n211), .Q(n173) );
  SDFFARX1 \AssembledTimerValue_reg[9]  ( .D(n384), .SI(n171), .SE(test_se), 
        .CLK(n10), .RSTB(n211), .Q(n172) );
  SDFFARX1 \AssembledTimerValue_reg[8]  ( .D(n385), .SI(n186), .SE(test_se), 
        .CLK(n10), .RSTB(n211), .Q(n171) );
  SDFFARX1 AddressOK_reg ( .D(n395), .SI(TxUsedDataOutDetected), .SE(test_se), 
        .CLK(n11), .RSTB(n211), .Q(AddressOK), .QN(n195) );
  SDFFARX1 ReceivedPauseFrmWAddr_reg ( .D(n394), .SI(Pause), .SE(test_se), 
        .CLK(n13), .RSTB(n211), .Q(n192), .QN(n7) );
  SDFFARX1 \LatchedTimerValue_reg[15]  ( .D(n362), .SI(n169), .SE(test_se), 
        .CLK(n13), .RSTB(n211), .Q(n170) );
  SDFFARX1 \LatchedTimerValue_reg[14]  ( .D(n363), .SI(n168), .SE(test_se), 
        .CLK(n12), .RSTB(n211), .Q(n169) );
  SDFFARX1 \LatchedTimerValue_reg[13]  ( .D(n364), .SI(n167), .SE(test_se), 
        .CLK(n12), .RSTB(n211), .Q(n168) );
  SDFFARX1 \LatchedTimerValue_reg[12]  ( .D(n365), .SI(n166), .SE(test_se), 
        .CLK(n12), .RSTB(n211), .Q(n167) );
  SDFFARX1 \LatchedTimerValue_reg[11]  ( .D(n366), .SI(n165), .SE(test_se), 
        .CLK(n12), .RSTB(n211), .Q(n166) );
  SDFFARX1 \LatchedTimerValue_reg[10]  ( .D(n367), .SI(n164), .SE(test_se), 
        .CLK(n12), .RSTB(n211), .Q(n165) );
  SDFFARX1 \LatchedTimerValue_reg[9]  ( .D(n368), .SI(n163), .SE(test_se), 
        .CLK(n12), .RSTB(n211), .Q(n164) );
  SDFFARX1 \LatchedTimerValue_reg[8]  ( .D(n369), .SI(n162), .SE(test_se), 
        .CLK(n12), .RSTB(n211), .Q(n163) );
  SDFFARX1 \LatchedTimerValue_reg[7]  ( .D(n370), .SI(n161), .SE(test_se), 
        .CLK(n12), .RSTB(n211), .Q(n162) );
  SDFFARX1 \LatchedTimerValue_reg[6]  ( .D(n371), .SI(n160), .SE(test_se), 
        .CLK(n12), .RSTB(n211), .Q(n161) );
  SDFFARX1 \LatchedTimerValue_reg[5]  ( .D(n372), .SI(n159), .SE(test_se), 
        .CLK(n12), .RSTB(n211), .Q(n160) );
  SDFFARX1 \LatchedTimerValue_reg[4]  ( .D(n373), .SI(n158), .SE(test_se), 
        .CLK(n12), .RSTB(n211), .Q(n159) );
  SDFFARX1 \LatchedTimerValue_reg[3]  ( .D(n374), .SI(n157), .SE(test_se), 
        .CLK(n12), .RSTB(n211), .Q(n158) );
  SDFFARX1 \LatchedTimerValue_reg[2]  ( .D(n375), .SI(n156), .SE(test_se), 
        .CLK(n12), .RSTB(n211), .Q(n157) );
  SDFFARX1 \LatchedTimerValue_reg[1]  ( .D(n376), .SI(n155), .SE(test_se), 
        .CLK(n11), .RSTB(n211), .Q(n156) );
  SDFFARX1 \LatchedTimerValue_reg[0]  ( .D(n377), .SI(n189), .SE(test_se), 
        .CLK(n11), .RSTB(n211), .Q(n155) );
  SDFFARX1 \SlotTimer_reg[0]  ( .D(n361), .SI(ReceivedPauseFrm), .SE(test_se), 
        .CLK(n9), .RSTB(n211), .Q(n203), .QN(n212) );
  SDFFARX1 \PauseTimer_reg[0]  ( .D(n359), .SI(n152), .SE(test_se), .CLK(n11), 
        .RSTB(n211), .Q(PauseTimer[0]), .QN(n214) );
  SDFFARX1 \PauseTimer_reg[1]  ( .D(n358), .SI(PauseTimer[0]), .SE(test_se), 
        .CLK(n13), .RSTB(n211), .Q(PauseTimer[1]), .QN(n216) );
  SDFFARX1 \PauseTimer_reg[2]  ( .D(n357), .SI(PauseTimer[1]), .SE(test_se), 
        .CLK(n13), .RSTB(n211), .Q(PauseTimer[2]), .QN(n218) );
  SDFFARX1 \PauseTimer_reg[3]  ( .D(n356), .SI(PauseTimer[2]), .SE(test_se), 
        .CLK(n13), .RSTB(n211), .Q(PauseTimer[3]), .QN(n220) );
  SDFFARX1 \PauseTimer_reg[4]  ( .D(n355), .SI(PauseTimer[3]), .SE(test_se), 
        .CLK(n13), .RSTB(n211), .Q(PauseTimer[4]), .QN(n222) );
  SDFFARX1 \PauseTimer_reg[5]  ( .D(n354), .SI(PauseTimer[4]), .SE(test_se), 
        .CLK(n13), .RSTB(n211), .Q(PauseTimer[5]), .QN(n224) );
  SDFFARX1 \PauseTimer_reg[6]  ( .D(n353), .SI(PauseTimer[5]), .SE(test_se), 
        .CLK(n13), .RSTB(n211), .Q(PauseTimer[6]), .QN(n226) );
  SDFFARX1 \PauseTimer_reg[7]  ( .D(n352), .SI(PauseTimer[6]), .SE(test_se), 
        .CLK(n13), .RSTB(n211), .Q(PauseTimer[7]), .QN(n228) );
  SDFFARX1 \PauseTimer_reg[8]  ( .D(n351), .SI(PauseTimer[7]), .SE(test_se), 
        .CLK(n13), .RSTB(n211), .Q(PauseTimer[8]), .QN(n230) );
  SDFFARX1 \PauseTimer_reg[9]  ( .D(n350), .SI(PauseTimer[8]), .SE(test_se), 
        .CLK(n13), .RSTB(n211), .Q(PauseTimer[9]), .QN(n232) );
  SDFFARX1 \PauseTimer_reg[10]  ( .D(n349), .SI(PauseTimer[9]), .SE(test_se), 
        .CLK(n13), .RSTB(n211), .Q(PauseTimer[10]), .QN(n234) );
  SDFFARX1 \PauseTimer_reg[11]  ( .D(n348), .SI(PauseTimer[10]), .SE(test_se), 
        .CLK(n14), .RSTB(n211), .Q(PauseTimer[11]), .QN(n236) );
  SDFFARX1 \PauseTimer_reg[12]  ( .D(n347), .SI(PauseTimer[11]), .SE(test_se), 
        .CLK(n14), .RSTB(n211), .Q(PauseTimer[12]), .QN(n238) );
  SDFFARX1 \PauseTimer_reg[13]  ( .D(n346), .SI(PauseTimer[12]), .SE(test_se), 
        .CLK(n14), .RSTB(n211), .Q(PauseTimer[13]), .QN(n240) );
  SDFFARX1 \PauseTimer_reg[14]  ( .D(n345), .SI(PauseTimer[13]), .SE(test_se), 
        .CLK(n14), .RSTB(n211), .Q(PauseTimer[14]), .QN(n242) );
  SDFFARX1 \PauseTimer_reg[15]  ( .D(n344), .SI(PauseTimer[14]), .SE(test_se), 
        .CLK(n9), .RSTB(n211), .Q(PauseTimer[15]), .QN(n244) );
  SDFFASX1 PauseTimerEq0_sync1_reg ( .D(n407), .SI(n204), .SE(test_se), .CLK(
        MTxClk), .SETB(n223), .Q(PauseTimerEq0_sync1) );
  SDFFASX1 PauseTimerEq0_sync2_reg ( .D(PauseTimerEq0_sync1), .SI(
        PauseTimerEq0_sync1), .SE(test_se), .CLK(MTxClk), .SETB(n223), .Q(n152) );
  SDFFARX1 Pause_reg ( .D(n260), .SI(PauseTimer[15]), .SE(test_se), .CLK(
        MTxClk), .RSTB(n223), .Q(Pause), .QN(n337) );
  SDFFARX1 Divider2_reg ( .D(N183), .SI(n188), .SE(test_se), .CLK(n11), .RSTB(
        n211), .Q(n154), .QN(n332) );
  SDFFARX1 \SlotTimer_reg[5]  ( .D(n360), .SI(n199), .SE(test_se), .CLK(n9), 
        .RSTB(n211), .Q(n198), .QN(n213) );
  SDFFARX1 \SlotTimer_reg[1]  ( .D(n343), .SI(n203), .SE(test_se), .CLK(n9), 
        .RSTB(n211), .Q(n202), .QN(n246) );
  SDFFARX1 \SlotTimer_reg[2]  ( .D(n342), .SI(n202), .SE(test_se), .CLK(n10), 
        .RSTB(n211), .Q(n201), .QN(n247) );
  SDFFARX1 \SlotTimer_reg[3]  ( .D(n341), .SI(n201), .SE(test_se), .CLK(n9), 
        .RSTB(n211), .Q(n200), .QN(n248) );
  SDFFARX1 \SlotTimer_reg[4]  ( .D(n340), .SI(n200), .SE(test_se), .CLK(n9), 
        .RSTB(n211), .Q(n199), .QN(n249) );
  SDFFARX1 ReceivedPauseFrm_reg ( .D(n339), .SI(n192), .SE(test_se), .CLK(n9), 
        .RSTB(n211), .Q(ReceivedPauseFrm), .QN(n250) );
  eth_receivecontrol_DW01_dec_0 sub_358 ( .A(PauseTimer), .SUM({N158, N157, 
        N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, 
        N144, N143}) );
  INVX2 U3 ( .INP(n197), .ZN(n211) );
  NBUFFX2 U4 ( .INP(MRxClk), .Z(n9) );
  NBUFFX2 U5 ( .INP(MRxClk), .Z(n12) );
  NBUFFX2 U6 ( .INP(MRxClk), .Z(n13) );
  NBUFFX2 U7 ( .INP(MRxClk), .Z(n10) );
  NBUFFX2 U8 ( .INP(MRxClk), .Z(n11) );
  NBUFFX2 U9 ( .INP(MRxClk), .Z(n14) );
  INVX0 U10 ( .INP(eth_top_test_point_11887_in), .ZN(n223) );
  MUX21X1 U11 ( .IN1(n15), .IN2(n16), .S(n6), .Q(n406) );
  AND2X1 U12 ( .IN1(n17), .IN2(n18), .Q(n15) );
  AO22X1 U13 ( .IN1(n19), .IN2(n189), .IN3(n20), .IN4(n16), .Q(n405) );
  NOR2X0 U14 ( .IN1(n6), .IN2(n297), .QN(n20) );
  MUX21X1 U15 ( .IN1(n19), .IN2(n21), .S(n297), .Q(n404) );
  NOR2X0 U16 ( .IN1(n6), .IN2(n17), .QN(n21) );
  INVX0 U17 ( .INP(n16), .ZN(n17) );
  MUX21X1 U18 ( .IN1(n18), .IN2(n6), .S(n16), .Q(n19) );
  NOR3X0 U19 ( .IN1(n22), .IN2(RxEndFrm), .IN3(n189), .QN(n16) );
  NAND2X0 U20 ( .IN1(RxEndFrm), .IN2(RxValid), .QN(n18) );
  MUX21X1 U21 ( .IN1(n23), .IN2(n24), .S(n3), .Q(n403) );
  MUX21X1 U22 ( .IN1(n25), .IN2(n26), .S(n219), .Q(n402) );
  NOR3X0 U23 ( .IN1(n27), .IN2(n333), .IN3(n28), .QN(n26) );
  AO21X1 U24 ( .IN1(n23), .IN2(n333), .IN3(n29), .Q(n25) );
  OA21X1 U25 ( .IN1(ReceiveEnd), .IN2(n188), .IN3(n30), .Q(n401) );
  MUX21X1 U26 ( .IN1(n31), .IN2(n32), .S(n4), .Q(n400) );
  NOR2X0 U27 ( .IN1(n336), .IN2(n28), .QN(n31) );
  MUX21X1 U28 ( .IN1(n33), .IN2(n34), .S(n1), .Q(n399) );
  AO21X1 U29 ( .IN1(n217), .IN2(n23), .IN3(n32), .Q(n34) );
  AO21X1 U30 ( .IN1(n23), .IN2(n336), .IN3(n24), .Q(n32) );
  AND3X1 U31 ( .IN1(n23), .IN2(n4), .IN3(n3), .Q(n33) );
  MUX21X1 U32 ( .IN1(n35), .IN2(n29), .S(n2), .Q(n398) );
  AO21X1 U33 ( .IN1(n23), .IN2(n27), .IN3(n24), .Q(n29) );
  NOR2X0 U34 ( .IN1(n23), .IN2(RxEndFrm), .QN(n24) );
  INVX0 U35 ( .INP(n28), .ZN(n23) );
  NOR2X0 U36 ( .IN1(n28), .IN2(n27), .QN(n35) );
  NAND3X0 U37 ( .IN1(n3), .IN2(n4), .IN3(n1), .QN(n27) );
  NAND4X0 U38 ( .IN1(RxValid), .IN2(n36), .IN3(n37), .IN4(n30), .QN(n28) );
  NOR2X0 U39 ( .IN1(n314), .IN2(RxEndFrm), .QN(n37) );
  NAND2X0 U40 ( .IN1(DlyCrcEn), .IN2(n8), .QN(n36) );
  OAI21X1 U41 ( .IN1(n215), .IN2(n38), .IN3(n39), .QN(n397) );
  NAND4X0 U42 ( .IN1(n40), .IN2(n41), .IN3(n336), .IN4(n42), .QN(n39) );
  OA22X1 U43 ( .IN1(n336), .IN2(n43), .IN3(n44), .IN4(n41), .Q(n38) );
  AND4X1 U44 ( .IN1(n45), .IN2(n2), .IN3(n1), .IN4(n4), .Q(n41) );
  INVX0 U45 ( .INP(n46), .ZN(n44) );
  MUX21X1 U46 ( .IN1(n47), .IN2(n48), .S(n49), .Q(n396) );
  NOR2X0 U47 ( .IN1(n333), .IN2(n50), .QN(n49) );
  NOR2X0 U48 ( .IN1(n51), .IN2(n52), .QN(n48) );
  NAND4X0 U49 ( .IN1(n53), .IN2(RxData[3]), .IN3(n42), .IN4(n54), .QN(n52) );
  MUX21X1 U50 ( .IN1(RxData[7]), .IN2(n55), .S(n3), .Q(n53) );
  NOR2X0 U51 ( .IN1(RxData[7]), .IN2(n5), .QN(n55) );
  OR4X1 U52 ( .IN1(RxData[2]), .IN2(RxData[4]), .IN3(RxData[5]), .IN4(
        RxData[6]), .Q(n51) );
  NOR2X0 U53 ( .IN1(n5), .IN2(ReceiveEnd), .QN(n47) );
  AO22X1 U54 ( .IN1(n56), .IN2(AddressOK), .IN3(n57), .IN4(n58), .Q(n395) );
  NAND2X0 U55 ( .IN1(n59), .IN2(n43), .QN(n58) );
  AO221X1 U56 ( .IN1(n60), .IN2(n42), .IN3(n61), .IN4(n62), .IN5(n63), .Q(n56)
         );
  MUX21X1 U57 ( .IN1(n64), .IN2(n65), .S(n66), .Q(n63) );
  NOR4X0 U58 ( .IN1(n61), .IN2(n67), .IN3(n68), .IN4(n69), .QN(n66) );
  NOR2X0 U59 ( .IN1(ReceiveEnd), .IN2(n57), .QN(n65) );
  INVX0 U60 ( .INP(n59), .ZN(n64) );
  NAND4X0 U61 ( .IN1(n70), .IN2(n71), .IN3(n72), .IN4(n73), .QN(n59) );
  NOR4X0 U62 ( .IN1(n74), .IN2(n75), .IN3(n76), .IN4(n77), .QN(n73) );
  XNOR2X1 U63 ( .IN1(RxData[3]), .IN2(n78), .Q(n77) );
  NOR2X0 U64 ( .IN1(n79), .IN2(n80), .QN(n78) );
  AO222X1 U65 ( .IN1(MAC[11]), .IN2(n81), .IN3(MAC[35]), .IN4(n67), .IN5(
        MAC[19]), .IN6(n82), .Q(n80) );
  AO222X1 U66 ( .IN1(MAC[43]), .IN2(n57), .IN3(MAC[3]), .IN4(n83), .IN5(
        MAC[27]), .IN6(n68), .Q(n79) );
  XNOR2X1 U67 ( .IN1(RxData[2]), .IN2(n84), .Q(n76) );
  NOR2X0 U68 ( .IN1(n85), .IN2(n86), .QN(n84) );
  AO222X1 U69 ( .IN1(MAC[10]), .IN2(n81), .IN3(MAC[34]), .IN4(n67), .IN5(
        MAC[18]), .IN6(n82), .Q(n86) );
  AO222X1 U70 ( .IN1(MAC[42]), .IN2(n57), .IN3(MAC[2]), .IN4(n83), .IN5(
        MAC[26]), .IN6(n68), .Q(n85) );
  XNOR2X1 U71 ( .IN1(RxData[1]), .IN2(n87), .Q(n75) );
  NOR2X0 U72 ( .IN1(n88), .IN2(n89), .QN(n87) );
  AO222X1 U73 ( .IN1(MAC[9]), .IN2(n81), .IN3(MAC[33]), .IN4(n67), .IN5(
        MAC[17]), .IN6(n82), .Q(n89) );
  AO222X1 U74 ( .IN1(MAC[41]), .IN2(n57), .IN3(MAC[1]), .IN4(n83), .IN5(
        MAC[25]), .IN6(n68), .Q(n88) );
  XNOR2X1 U75 ( .IN1(RxData[0]), .IN2(n90), .Q(n74) );
  NOR2X0 U76 ( .IN1(n91), .IN2(n92), .QN(n90) );
  AO222X1 U77 ( .IN1(MAC[8]), .IN2(n81), .IN3(MAC[32]), .IN4(n67), .IN5(
        MAC[16]), .IN6(n82), .Q(n92) );
  AO222X1 U78 ( .IN1(MAC[40]), .IN2(n57), .IN3(MAC[0]), .IN4(n83), .IN5(
        MAC[24]), .IN6(n68), .Q(n91) );
  NOR2X0 U79 ( .IN1(n93), .IN2(n94), .QN(n72) );
  XNOR2X1 U80 ( .IN1(RxData[5]), .IN2(n95), .Q(n94) );
  NOR2X0 U81 ( .IN1(n96), .IN2(n97), .QN(n95) );
  AO222X1 U82 ( .IN1(MAC[13]), .IN2(n81), .IN3(MAC[37]), .IN4(n67), .IN5(
        MAC[21]), .IN6(n82), .Q(n97) );
  AO222X1 U83 ( .IN1(MAC[45]), .IN2(n57), .IN3(MAC[5]), .IN4(n83), .IN5(
        MAC[29]), .IN6(n68), .Q(n96) );
  XNOR2X1 U84 ( .IN1(RxData[4]), .IN2(n98), .Q(n93) );
  NOR2X0 U85 ( .IN1(n99), .IN2(n100), .QN(n98) );
  AO222X1 U86 ( .IN1(MAC[12]), .IN2(n81), .IN3(MAC[36]), .IN4(n67), .IN5(
        MAC[20]), .IN6(n82), .Q(n100) );
  AO222X1 U87 ( .IN1(MAC[44]), .IN2(n57), .IN3(MAC[4]), .IN4(n83), .IN5(
        MAC[28]), .IN6(n68), .Q(n99) );
  XOR2X1 U88 ( .IN1(RxData[6]), .IN2(n101), .Q(n71) );
  NOR2X0 U89 ( .IN1(n102), .IN2(n103), .QN(n101) );
  AO222X1 U90 ( .IN1(MAC[14]), .IN2(n81), .IN3(MAC[38]), .IN4(n67), .IN5(
        MAC[22]), .IN6(n82), .Q(n103) );
  AO222X1 U91 ( .IN1(MAC[46]), .IN2(n57), .IN3(MAC[6]), .IN4(n83), .IN5(
        MAC[30]), .IN6(n68), .Q(n102) );
  XNOR2X1 U92 ( .IN1(n104), .IN2(n105), .Q(n70) );
  NOR2X0 U93 ( .IN1(n106), .IN2(n107), .QN(n105) );
  AO222X1 U94 ( .IN1(MAC[15]), .IN2(n81), .IN3(MAC[39]), .IN4(n67), .IN5(
        MAC[23]), .IN6(n82), .Q(n107) );
  AO222X1 U95 ( .IN1(MAC[47]), .IN2(n57), .IN3(MAC[7]), .IN4(n83), .IN5(
        MAC[31]), .IN6(n68), .Q(n106) );
  NOR4X0 U96 ( .IN1(n69), .IN2(n68), .IN3(n67), .IN4(n57), .QN(n83) );
  INVX0 U97 ( .INP(n108), .ZN(n67) );
  INVX0 U98 ( .INP(n109), .ZN(n68) );
  AND3X1 U99 ( .IN1(n217), .IN2(n336), .IN3(n110), .Q(n57) );
  INVX0 U100 ( .INP(n43), .ZN(n62) );
  NAND2X0 U101 ( .IN1(RxData[0]), .IN2(n40), .QN(n43) );
  NOR3X0 U102 ( .IN1(n2), .IN2(n336), .IN3(n50), .QN(n61) );
  INVX0 U103 ( .INP(RxData[0]), .ZN(n42) );
  AO22X1 U104 ( .IN1(n40), .IN2(n69), .IN3(n111), .IN4(n112), .Q(n60) );
  MUX21X1 U105 ( .IN1(n113), .IN2(n114), .S(RxData[6]), .Q(n112) );
  NOR2X0 U106 ( .IN1(n109), .IN2(n54), .QN(n114) );
  INVX0 U107 ( .INP(RxData[1]), .ZN(n54) );
  NAND3X0 U108 ( .IN1(n336), .IN2(n4), .IN3(n110), .QN(n109) );
  NOR2X0 U109 ( .IN1(RxData[1]), .IN2(n108), .QN(n113) );
  NAND3X0 U110 ( .IN1(n217), .IN2(n3), .IN3(n110), .QN(n108) );
  NOR2X0 U111 ( .IN1(n115), .IN2(n104), .QN(n111) );
  INVX0 U112 ( .INP(RxData[7]), .ZN(n104) );
  OR2X1 U113 ( .IN1(n82), .IN2(n81), .Q(n69) );
  NOR3X0 U114 ( .IN1(n3), .IN2(n2), .IN3(n50), .QN(n81) );
  NAND3X0 U115 ( .IN1(n217), .IN2(n1), .IN3(n45), .QN(n50) );
  AND3X1 U116 ( .IN1(n3), .IN2(n4), .IN3(n110), .Q(n82) );
  AND3X1 U117 ( .IN1(n334), .IN2(n333), .IN3(n45), .Q(n110) );
  AND3X1 U118 ( .IN1(RxValid), .IN2(n188), .IN3(n219), .Q(n45) );
  NOR4X0 U119 ( .IN1(n115), .IN2(RxData[1]), .IN3(RxData[6]), .IN4(RxData[7]), 
        .QN(n40) );
  OR4X1 U120 ( .IN1(RxData[2]), .IN2(RxData[3]), .IN3(RxData[4]), .IN4(
        RxData[5]), .Q(n115) );
  MUX21X1 U121 ( .IN1(n116), .IN2(n192), .S(n117), .Q(n394) );
  NOR2X0 U122 ( .IN1(n118), .IN2(ReceiveEnd), .QN(n117) );
  NOR4X0 U123 ( .IN1(n215), .IN2(n5), .IN3(n195), .IN4(n46), .QN(n118) );
  AO22X1 U124 ( .IN1(n119), .IN2(n179), .IN3(n120), .IN4(RxData[0]), .Q(n393)
         );
  AO22X1 U125 ( .IN1(n119), .IN2(n180), .IN3(n120), .IN4(RxData[1]), .Q(n392)
         );
  AO22X1 U126 ( .IN1(n119), .IN2(n181), .IN3(n120), .IN4(RxData[2]), .Q(n391)
         );
  AO22X1 U127 ( .IN1(n119), .IN2(n182), .IN3(n120), .IN4(RxData[3]), .Q(n390)
         );
  AO22X1 U128 ( .IN1(n119), .IN2(n183), .IN3(n120), .IN4(RxData[4]), .Q(n389)
         );
  AO22X1 U129 ( .IN1(n119), .IN2(n184), .IN3(n120), .IN4(RxData[5]), .Q(n388)
         );
  AO22X1 U130 ( .IN1(n119), .IN2(n185), .IN3(n120), .IN4(RxData[6]), .Q(n387)
         );
  AO22X1 U131 ( .IN1(n119), .IN2(n186), .IN3(n120), .IN4(RxData[7]), .Q(n386)
         );
  NOR2X0 U132 ( .IN1(n119), .IN2(RxStartFrm), .QN(n120) );
  AND2X1 U133 ( .IN1(n121), .IN2(n122), .Q(n119) );
  NAND4X0 U134 ( .IN1(n217), .IN2(n123), .IN3(n188), .IN4(n3), .QN(n121) );
  AO22X1 U135 ( .IN1(n124), .IN2(n171), .IN3(n125), .IN4(RxData[0]), .Q(n385)
         );
  AO22X1 U136 ( .IN1(n124), .IN2(n172), .IN3(n125), .IN4(RxData[1]), .Q(n384)
         );
  AO22X1 U137 ( .IN1(n124), .IN2(n173), .IN3(n125), .IN4(RxData[2]), .Q(n383)
         );
  AO22X1 U138 ( .IN1(n124), .IN2(n174), .IN3(n125), .IN4(RxData[3]), .Q(n382)
         );
  AO22X1 U139 ( .IN1(n124), .IN2(n175), .IN3(n125), .IN4(RxData[4]), .Q(n381)
         );
  AO22X1 U140 ( .IN1(n124), .IN2(n176), .IN3(n125), .IN4(RxData[5]), .Q(n380)
         );
  AO22X1 U141 ( .IN1(n124), .IN2(n177), .IN3(n125), .IN4(RxData[6]), .Q(n379)
         );
  AO22X1 U142 ( .IN1(n124), .IN2(n178), .IN3(n125), .IN4(RxData[7]), .Q(n378)
         );
  NOR2X0 U143 ( .IN1(n124), .IN2(RxStartFrm), .QN(n125) );
  OA21X1 U144 ( .IN1(n46), .IN2(n314), .IN3(n122), .Q(n124) );
  INVX0 U145 ( .INP(RxStartFrm), .ZN(n122) );
  AO22X1 U146 ( .IN1(n126), .IN2(n179), .IN3(n127), .IN4(n155), .Q(n377) );
  AO22X1 U147 ( .IN1(n126), .IN2(n180), .IN3(n127), .IN4(n156), .Q(n376) );
  AO22X1 U148 ( .IN1(n126), .IN2(n181), .IN3(n127), .IN4(n157), .Q(n375) );
  AO22X1 U149 ( .IN1(n126), .IN2(n182), .IN3(n127), .IN4(n158), .Q(n374) );
  AO22X1 U150 ( .IN1(n126), .IN2(n183), .IN3(n127), .IN4(n159), .Q(n373) );
  AO22X1 U151 ( .IN1(n126), .IN2(n184), .IN3(n127), .IN4(n160), .Q(n372) );
  AO22X1 U152 ( .IN1(n126), .IN2(n185), .IN3(n127), .IN4(n161), .Q(n371) );
  AO22X1 U153 ( .IN1(n126), .IN2(n186), .IN3(n127), .IN4(n162), .Q(n370) );
  AO22X1 U154 ( .IN1(n126), .IN2(n171), .IN3(n127), .IN4(n163), .Q(n369) );
  AO22X1 U155 ( .IN1(n126), .IN2(n172), .IN3(n127), .IN4(n164), .Q(n368) );
  AO22X1 U156 ( .IN1(n126), .IN2(n173), .IN3(n127), .IN4(n165), .Q(n367) );
  AO22X1 U157 ( .IN1(n126), .IN2(n174), .IN3(n127), .IN4(n166), .Q(n366) );
  AO22X1 U158 ( .IN1(n126), .IN2(n175), .IN3(n127), .IN4(n167), .Q(n365) );
  AO22X1 U159 ( .IN1(n126), .IN2(n176), .IN3(n127), .IN4(n168), .Q(n364) );
  AO22X1 U160 ( .IN1(n126), .IN2(n177), .IN3(n127), .IN4(n169), .Q(n363) );
  AO22X1 U161 ( .IN1(n126), .IN2(n178), .IN3(n127), .IN4(n170), .Q(n362) );
  NOR2X0 U162 ( .IN1(n126), .IN2(ReceiveEnd), .QN(n127) );
  NOR2X0 U163 ( .IN1(n30), .IN2(n7), .QN(n126) );
  NAND4X0 U164 ( .IN1(n336), .IN2(n123), .IN3(n188), .IN4(n4), .QN(n30) );
  MUX21X1 U165 ( .IN1(n128), .IN2(n129), .S(n212), .Q(n361) );
  MUX21X1 U166 ( .IN1(n130), .IN2(n131), .S(n213), .Q(n360) );
  AND2X1 U167 ( .IN1(n129), .IN2(n132), .Q(n131) );
  AO21X1 U168 ( .IN1(n249), .IN2(n129), .IN3(n133), .Q(n130) );
  AO222X1 U169 ( .IN1(N143), .IN2(n134), .IN3(n135), .IN4(PauseTimer[0]), 
        .IN5(SetPauseTimer), .IN6(n155), .Q(n359) );
  AO222X1 U170 ( .IN1(N144), .IN2(n134), .IN3(n135), .IN4(PauseTimer[1]), 
        .IN5(SetPauseTimer), .IN6(n156), .Q(n358) );
  AO222X1 U171 ( .IN1(N145), .IN2(n134), .IN3(n135), .IN4(PauseTimer[2]), 
        .IN5(SetPauseTimer), .IN6(n157), .Q(n357) );
  AO222X1 U172 ( .IN1(N146), .IN2(n134), .IN3(n135), .IN4(PauseTimer[3]), 
        .IN5(SetPauseTimer), .IN6(n158), .Q(n356) );
  AO222X1 U173 ( .IN1(N147), .IN2(n134), .IN3(n135), .IN4(PauseTimer[4]), 
        .IN5(SetPauseTimer), .IN6(n159), .Q(n355) );
  AO222X1 U174 ( .IN1(N148), .IN2(n134), .IN3(n135), .IN4(PauseTimer[5]), 
        .IN5(SetPauseTimer), .IN6(n160), .Q(n354) );
  AO222X1 U175 ( .IN1(N149), .IN2(n134), .IN3(n135), .IN4(PauseTimer[6]), 
        .IN5(SetPauseTimer), .IN6(n161), .Q(n353) );
  AO222X1 U176 ( .IN1(N150), .IN2(n134), .IN3(n135), .IN4(PauseTimer[7]), 
        .IN5(SetPauseTimer), .IN6(n162), .Q(n352) );
  AO222X1 U177 ( .IN1(N151), .IN2(n134), .IN3(n135), .IN4(PauseTimer[8]), 
        .IN5(SetPauseTimer), .IN6(n163), .Q(n351) );
  AO222X1 U178 ( .IN1(N152), .IN2(n134), .IN3(n135), .IN4(PauseTimer[9]), 
        .IN5(SetPauseTimer), .IN6(n164), .Q(n350) );
  AO222X1 U179 ( .IN1(N153), .IN2(n134), .IN3(n135), .IN4(PauseTimer[10]), 
        .IN5(SetPauseTimer), .IN6(n165), .Q(n349) );
  AO222X1 U180 ( .IN1(N154), .IN2(n134), .IN3(n135), .IN4(PauseTimer[11]), 
        .IN5(SetPauseTimer), .IN6(n166), .Q(n348) );
  AO222X1 U181 ( .IN1(N155), .IN2(n134), .IN3(n135), .IN4(PauseTimer[12]), 
        .IN5(SetPauseTimer), .IN6(n167), .Q(n347) );
  AO222X1 U182 ( .IN1(N156), .IN2(n134), .IN3(n135), .IN4(PauseTimer[13]), 
        .IN5(SetPauseTimer), .IN6(n168), .Q(n346) );
  AO222X1 U183 ( .IN1(N157), .IN2(n134), .IN3(n135), .IN4(PauseTimer[14]), 
        .IN5(SetPauseTimer), .IN6(n169), .Q(n345) );
  AO222X1 U184 ( .IN1(N158), .IN2(n134), .IN3(n135), .IN4(PauseTimer[15]), 
        .IN5(SetPauseTimer), .IN6(n170), .Q(n344) );
  NOR2X0 U185 ( .IN1(SetPauseTimer), .IN2(n134), .QN(n135) );
  INVX0 U186 ( .INP(n136), .ZN(SetPauseTimer) );
  AND4X1 U187 ( .IN1(RxFlow), .IN2(n136), .IN3(n132), .IN4(n137), .Q(n134) );
  NOR4X0 U188 ( .IN1(n337), .IN2(n332), .IN3(n213), .IN4(n407), .QN(n137) );
  NOR3X0 U189 ( .IN1(n248), .IN2(n249), .IN3(n138), .QN(n132) );
  NAND4X0 U190 ( .IN1(RxFlow), .IN2(ReceivedPacketGood), .IN3(n139), .IN4(
        ReceivedLengthOK), .QN(n136) );
  NOR2X0 U191 ( .IN1(n7), .IN2(n116), .QN(n139) );
  INVX0 U192 ( .INP(ReceiveEnd), .ZN(n116) );
  MUX21X1 U193 ( .IN1(n140), .IN2(n141), .S(n246), .Q(n343) );
  NOR2X0 U194 ( .IN1(n212), .IN2(n142), .QN(n141) );
  MUX21X1 U195 ( .IN1(n143), .IN2(n144), .S(n247), .Q(n342) );
  NOR3X0 U196 ( .IN1(n142), .IN2(n246), .IN3(n212), .QN(n144) );
  AO21X1 U197 ( .IN1(n246), .IN2(n129), .IN3(n140), .Q(n143) );
  AO21X1 U198 ( .IN1(n212), .IN2(n129), .IN3(n128), .Q(n140) );
  MUX21X1 U199 ( .IN1(n145), .IN2(n146), .S(n248), .Q(n341) );
  NOR2X0 U200 ( .IN1(n142), .IN2(n138), .QN(n146) );
  MUX21X1 U201 ( .IN1(n133), .IN2(n147), .S(n249), .Q(n340) );
  NOR3X0 U202 ( .IN1(n138), .IN2(n248), .IN3(n142), .QN(n147) );
  INVX0 U203 ( .INP(n129), .ZN(n142) );
  AO21X1 U204 ( .IN1(n248), .IN2(n129), .IN3(n145), .Q(n133) );
  AO21X1 U205 ( .IN1(n129), .IN2(n138), .IN3(n128), .Q(n145) );
  NOR2X0 U206 ( .IN1(n129), .IN2(RxReset), .QN(n128) );
  OR3X1 U207 ( .IN1(n246), .IN2(n247), .IN3(n212), .Q(n138) );
  NOR4X0 U208 ( .IN1(n148), .IN2(RxReset), .IN3(n332), .IN4(n337), .QN(n129)
         );
  MUX21X1 U209 ( .IN1(n149), .IN2(n150), .S(n250), .Q(n339) );
  NOR4X0 U210 ( .IN1(n215), .IN2(n5), .IN3(n151), .IN4(n46), .QN(n150) );
  NAND3X0 U211 ( .IN1(n336), .IN2(n123), .IN3(n217), .QN(n46) );
  NOR4X0 U212 ( .IN1(n1), .IN2(n2), .IN3(n22), .IN4(n219), .QN(n123) );
  INVX0 U213 ( .INP(RxValid), .ZN(n22) );
  AND2X1 U214 ( .IN1(RxStatusWriteLatched_sync2), .IN2(r_PassAll), .Q(n151) );
  NOR2X0 U215 ( .IN1(RxStatusWriteLatched_sync2), .IN2(n153), .QN(n149) );
  INVX0 U216 ( .INP(r_PassAll), .ZN(n153) );
  MUX21X1 U217 ( .IN1(Pause), .IN2(n193), .S(n194), .Q(n260) );
  AOI21X1 U218 ( .IN1(n196), .IN2(TxUsedDataOutDetected), .IN3(TxStartFrmOut), 
        .QN(n194) );
  NOR2X0 U219 ( .IN1(TxDoneIn), .IN2(TxAbortIn), .QN(n196) );
  NOR2X0 U220 ( .IN1(n148), .IN2(n152), .QN(n193) );
  INVX0 U221 ( .INP(RxFlow), .ZN(n148) );
  MUX21X1 U222 ( .IN1(RxReset), .IN2(eth_top_data_sourcea_in), .S(
        eth_top_test_mode_in), .Q(n197) );
  AND3X1 U223 ( .IN1(n332), .IN2(n206), .IN3(RxFlow), .Q(N183) );
  INVX0 U224 ( .INP(n407), .ZN(n206) );
  NOR4X0 U225 ( .IN1(n207), .IN2(n208), .IN3(n209), .IN4(n210), .QN(n407) );
  NAND4X0 U226 ( .IN1(n228), .IN2(n226), .IN3(n224), .IN4(n222), .QN(n210) );
  NAND4X0 U227 ( .IN1(n220), .IN2(n218), .IN3(n216), .IN4(n214), .QN(n209) );
  NAND4X0 U228 ( .IN1(n244), .IN2(n242), .IN3(n240), .IN4(n238), .QN(n208) );
  NAND4X0 U229 ( .IN1(n236), .IN2(n234), .IN3(n232), .IN4(n230), .QN(n207) );
endmodule


module eth_transmitcontrol_test_1 ( MTxClk, TxReset, TxUsedDataIn, 
        TxUsedDataOut, TxDoneIn, TxAbortIn, TxStartFrmIn, TPauseRq, 
        TxUsedDataOutDetected, TxFlow, DlyCrcEn, TxPauseTV, MAC, 
        TxCtrlStartFrm, TxCtrlEndFrm, SendingCtrlFrm, CtrlMux, ControlData, 
        WillSendControlFrame, BlockTxDone, eth_top_test_point_11887_in, 
        test_si, test_se );
  input [15:0] TxPauseTV;
  input [47:0] MAC;
  output [7:0] ControlData;
  input MTxClk, TxReset, TxUsedDataIn, TxUsedDataOut, TxDoneIn, TxAbortIn,
         TxStartFrmIn, TPauseRq, TxUsedDataOutDetected, TxFlow, DlyCrcEn,
         eth_top_test_point_11887_in, test_si, test_se;
  output TxCtrlStartFrm, TxCtrlEndFrm, SendingCtrlFrm, CtrlMux,
         WillSendControlFrame, BlockTxDone;
  wire   N31, n38, n39, n41, n42, n45, n46, n48, n49, n50, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n1, n2, n3, n4, n5,
         n32, n33, n169, n171, n172, n175, n176, n177, n178, n179, n160, n162,
         n163, n165, n167, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n34, n35, n36, n37, n40, n43, n44, n47, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n154;

  SDFFARX1 TxUsedDataIn_q_reg ( .D(TxUsedDataIn), .SI(TxCtrlStartFrm), .SE(
        test_se), .CLK(MTxClk), .RSTB(n154), .Q(n175), .QN(n129) );
  SDFFARX1 \ByteCnt_reg[0]  ( .D(n153), .SI(BlockTxDone), .SE(test_se), .CLK(
        MTxClk), .RSTB(n154), .Q(n32), .QN(n50) );
  SDFFX1 ControlEnd_q_reg ( .D(n131), .SI(ControlData[7]), .SE(test_se), .CLK(
        MTxClk), .Q(n179), .QN(n172) );
  SDFFARX1 TxCtrlEndFrm_reg ( .D(N31), .SI(SendingCtrlFrm), .SE(test_se), 
        .CLK(MTxClk), .RSTB(n154), .Q(TxCtrlEndFrm), .QN(n169) );
  SDFFARX1 WillSendControlFrame_reg ( .D(n151), .SI(n175), .SE(test_se), .CLK(
        MTxClk), .RSTB(n154), .Q(WillSendControlFrame) );
  SDFFARX1 CtrlMux_reg ( .D(n150), .SI(n179), .SE(test_se), .CLK(MTxClk), 
        .RSTB(n154), .Q(CtrlMux), .QN(n171) );
  SDFFARX1 TxCtrlStartFrm_reg ( .D(n149), .SI(n176), .SE(test_se), .CLK(MTxClk), .RSTB(n154), .Q(TxCtrlStartFrm) );
  SDFFX1 TxCtrlStartFrm_q_reg ( .D(TxCtrlStartFrm), .SI(TxCtrlEndFrm), .SE(
        test_se), .CLK(MTxClk), .Q(n176), .QN(n38) );
  SDFFARX1 BlockTxDone_reg ( .D(n148), .SI(test_si), .SE(test_se), .CLK(MTxClk), .RSTB(n154), .Q(BlockTxDone) );
  SDFFARX1 SendingCtrlFrm_reg ( .D(n140), .SI(n33), .SE(test_se), .CLK(MTxClk), 
        .RSTB(n154), .Q(SendingCtrlFrm) );
  SDFFARX1 \DlyCrcCnt_reg[0]  ( .D(n147), .SI(CtrlMux), .SE(test_se), .CLK(
        MTxClk), .RSTB(n154), .Q(n178), .QN(n42) );
  SDFFARX1 \DlyCrcCnt_reg[1]  ( .D(n146), .SI(n178), .SE(test_se), .CLK(MTxClk), .RSTB(n154), .Q(n177), .QN(n41) );
  SDFFARX1 \DlyCrcCnt_reg[2]  ( .D(n145), .SI(n177), .SE(test_se), .CLK(MTxClk), .RSTB(n154), .Q(n33), .QN(n39) );
  SDFFARX1 \ByteCnt_reg[4]  ( .D(n141), .SI(n5), .SE(test_se), .CLK(MTxClk), 
        .RSTB(n154), .Q(n3), .QN(n46) );
  SDFFARX1 \ByteCnt_reg[1]  ( .D(n144), .SI(n32), .SE(test_se), .CLK(MTxClk), 
        .RSTB(n154), .Q(n4), .QN(n49) );
  SDFFARX1 \ByteCnt_reg[2]  ( .D(n143), .SI(n4), .SE(test_se), .CLK(MTxClk), 
        .RSTB(n154), .Q(n2), .QN(n48) );
  SDFFARX1 \ByteCnt_reg[3]  ( .D(n142), .SI(n2), .SE(test_se), .CLK(MTxClk), 
        .RSTB(n154), .Q(n5), .QN(n130) );
  SDFFARX1 \ByteCnt_reg[5]  ( .D(n152), .SI(n3), .SE(test_se), .CLK(MTxClk), 
        .RSTB(n154), .Q(n1), .QN(n45) );
  SDFFARX1 \ControlData_reg[7]  ( .D(n139), .SI(ControlData[6]), .SE(test_se), 
        .CLK(MTxClk), .RSTB(n154), .Q(ControlData[7]), .QN(n160) );
  SDFFARX1 \ControlData_reg[6]  ( .D(n138), .SI(ControlData[5]), .SE(test_se), 
        .CLK(MTxClk), .RSTB(n154), .Q(ControlData[6]) );
  SDFFARX1 \ControlData_reg[5]  ( .D(n137), .SI(ControlData[4]), .SE(test_se), 
        .CLK(MTxClk), .RSTB(n154), .Q(ControlData[5]), .QN(n162) );
  SDFFARX1 \ControlData_reg[4]  ( .D(n136), .SI(ControlData[3]), .SE(test_se), 
        .CLK(MTxClk), .RSTB(n154), .Q(ControlData[4]), .QN(n163) );
  SDFFARX1 \ControlData_reg[3]  ( .D(n135), .SI(ControlData[2]), .SE(test_se), 
        .CLK(MTxClk), .RSTB(n154), .Q(ControlData[3]) );
  SDFFARX1 \ControlData_reg[2]  ( .D(n134), .SI(ControlData[1]), .SE(test_se), 
        .CLK(MTxClk), .RSTB(n154), .Q(ControlData[2]), .QN(n165) );
  SDFFARX1 \ControlData_reg[1]  ( .D(n133), .SI(ControlData[0]), .SE(test_se), 
        .CLK(MTxClk), .RSTB(n154), .Q(ControlData[1]) );
  SDFFARX1 \ControlData_reg[0]  ( .D(n132), .SI(n1), .SE(test_se), .CLK(MTxClk), .RSTB(n154), .Q(ControlData[0]), .QN(n167) );
  INVX0 U3 ( .INP(eth_top_test_point_11887_in), .ZN(n154) );
  MUX21X1 U4 ( .IN1(n6), .IN2(n7), .S(n50), .Q(n153) );
  NOR2X0 U5 ( .IN1(n8), .IN2(n9), .QN(n7) );
  AO21X1 U6 ( .IN1(n8), .IN2(n10), .IN3(n11), .Q(n6) );
  INVX0 U7 ( .INP(n12), .ZN(n8) );
  MUX21X1 U8 ( .IN1(n13), .IN2(n14), .S(n45), .Q(n152) );
  NOR3X0 U9 ( .IN1(n15), .IN2(n46), .IN3(n9), .QN(n14) );
  AO21X1 U10 ( .IN1(n10), .IN2(n46), .IN3(n16), .Q(n13) );
  OA22X1 U11 ( .IN1(n17), .IN2(WillSendControlFrame), .IN3(n169), .IN4(n171), 
        .Q(n151) );
  AND2X1 U12 ( .IN1(TxFlow), .IN2(TPauseRq), .Q(n17) );
  AO22X1 U13 ( .IN1(n18), .IN2(WillSendControlFrame), .IN3(n19), .IN4(CtrlMux), 
        .Q(n150) );
  MUX21X1 U14 ( .IN1(n20), .IN2(TxCtrlStartFrm), .S(n21), .Q(n149) );
  OA21X1 U15 ( .IN1(n129), .IN2(n171), .IN3(n22), .Q(n21) );
  NAND3X0 U16 ( .IN1(n18), .IN2(WillSendControlFrame), .IN3(n23), .QN(n22) );
  NAND3X0 U17 ( .IN1(n24), .IN2(n25), .IN3(TxUsedDataOutDetected), .QN(n23) );
  INVX0 U18 ( .INP(TxUsedDataOut), .ZN(n18) );
  OR2X1 U19 ( .IN1(n129), .IN2(n171), .Q(n20) );
  AO21X1 U20 ( .IN1(n25), .IN2(BlockTxDone), .IN3(TxCtrlStartFrm), .Q(n148) );
  INVX0 U21 ( .INP(TxStartFrmIn), .ZN(n25) );
  MUX21X1 U22 ( .IN1(n26), .IN2(n27), .S(n42), .Q(n147) );
  NOR2X0 U23 ( .IN1(n27), .IN2(n28), .QN(n26) );
  MUX21X1 U24 ( .IN1(n29), .IN2(n30), .S(n41), .Q(n146) );
  NOR2X0 U25 ( .IN1(n42), .IN2(n31), .QN(n30) );
  AO22X1 U26 ( .IN1(n29), .IN2(n33), .IN3(n34), .IN4(n27), .Q(n145) );
  INVX0 U27 ( .INP(n31), .ZN(n27) );
  NOR2X0 U28 ( .IN1(n42), .IN2(n41), .QN(n34) );
  MUX21X1 U29 ( .IN1(n42), .IN2(n35), .S(n31), .Q(n29) );
  NAND4X0 U30 ( .IN1(n39), .IN2(n35), .IN3(TxUsedDataIn), .IN4(CtrlMux), .QN(
        n31) );
  AO22X1 U31 ( .IN1(n11), .IN2(n4), .IN3(n36), .IN4(n10), .Q(n144) );
  XOR3X1 U32 ( .IN1(n12), .IN2(n4), .IN3(n37), .Q(n36) );
  MUX21X1 U33 ( .IN1(n40), .IN2(n43), .S(n48), .Q(n143) );
  NOR2X0 U34 ( .IN1(n9), .IN2(n44), .QN(n43) );
  MUX21X1 U35 ( .IN1(n47), .IN2(n51), .S(n130), .Q(n142) );
  NOR3X0 U36 ( .IN1(n44), .IN2(n48), .IN3(n9), .QN(n51) );
  AO21X1 U37 ( .IN1(n10), .IN2(n48), .IN3(n40), .Q(n47) );
  AO21X1 U38 ( .IN1(n10), .IN2(n44), .IN3(n11), .Q(n40) );
  MUX21X1 U39 ( .IN1(n16), .IN2(n52), .S(n46), .Q(n141) );
  NOR2X0 U40 ( .IN1(n9), .IN2(n15), .QN(n52) );
  AO21X1 U41 ( .IN1(n10), .IN2(n15), .IN3(n11), .Q(n16) );
  NOR2X0 U42 ( .IN1(n28), .IN2(n10), .QN(n11) );
  INVX0 U43 ( .INP(n35), .ZN(n28) );
  OR3X1 U44 ( .IN1(n48), .IN2(n130), .IN3(n44), .Q(n15) );
  AO21X1 U45 ( .IN1(n37), .IN2(n12), .IN3(n49), .Q(n44) );
  NAND2X0 U46 ( .IN1(n32), .IN2(n12), .QN(n37) );
  NAND2X0 U47 ( .IN1(n53), .IN2(TxUsedDataIn), .QN(n12) );
  INVX0 U48 ( .INP(n9), .ZN(n10) );
  NAND4X0 U49 ( .IN1(n35), .IN2(n54), .IN3(n55), .IN4(CtrlMux), .QN(n9) );
  AO21X1 U50 ( .IN1(TxUsedDataIn), .IN2(n56), .IN3(n53), .Q(n55) );
  AND2X1 U51 ( .IN1(n38), .IN2(TxCtrlStartFrm), .Q(n53) );
  INVX0 U52 ( .INP(n57), .ZN(n54) );
  OA21X1 U53 ( .IN1(TxCtrlStartFrm), .IN2(n24), .IN3(n58), .Q(n35) );
  INVX0 U54 ( .INP(TxReset), .ZN(n58) );
  NOR2X0 U55 ( .IN1(TxAbortIn), .IN2(TxDoneIn), .QN(n24) );
  AO22X1 U56 ( .IN1(WillSendControlFrame), .IN2(TxCtrlStartFrm), .IN3(n19), 
        .IN4(SendingCtrlFrm), .Q(n140) );
  INVX0 U57 ( .INP(TxDoneIn), .ZN(n19) );
  NAND2X0 U58 ( .IN1(n59), .IN2(n60), .QN(n139) );
  NAND2X0 U59 ( .IN1(TxPauseTV[7]), .IN2(n131), .QN(n60) );
  MUX21X1 U60 ( .IN1(n160), .IN2(n61), .S(n50), .Q(n59) );
  NOR2X0 U61 ( .IN1(n62), .IN2(n63), .QN(n61) );
  AO221X1 U62 ( .IN1(MAC[39]), .IN2(n64), .IN3(MAC[47]), .IN4(n65), .IN5(n66), 
        .Q(n63) );
  AO22X1 U63 ( .IN1(MAC[7]), .IN2(n67), .IN3(MAC[15]), .IN4(n68), .Q(n66) );
  AO221X1 U64 ( .IN1(TxPauseTV[15]), .IN2(n69), .IN3(MAC[31]), .IN4(n70), 
        .IN5(n71), .Q(n62) );
  AO221X1 U65 ( .IN1(n72), .IN2(n45), .IN3(MAC[23]), .IN4(n73), .IN5(n74), .Q(
        n71) );
  OA21X1 U66 ( .IN1(n75), .IN2(n76), .IN3(n48), .Q(n72) );
  NOR3X0 U67 ( .IN1(n4), .IN2(n130), .IN3(n46), .QN(n75) );
  AO21X1 U68 ( .IN1(TxPauseTV[6]), .IN2(n131), .IN3(n77), .Q(n138) );
  MUX21X1 U69 ( .IN1(ControlData[6]), .IN2(n78), .S(n50), .Q(n77) );
  NAND4X0 U70 ( .IN1(n79), .IN2(n80), .IN3(n81), .IN4(n82), .QN(n78) );
  AOI221X1 U71 ( .IN1(MAC[38]), .IN2(n64), .IN3(MAC[46]), .IN4(n65), .IN5(n83), 
        .QN(n82) );
  AO22X1 U72 ( .IN1(MAC[6]), .IN2(n67), .IN3(MAC[14]), .IN4(n68), .Q(n83) );
  AOI22X1 U73 ( .IN1(TxPauseTV[14]), .IN2(n69), .IN3(MAC[30]), .IN4(n70), .QN(
        n81) );
  NAND2X0 U74 ( .IN1(MAC[22]), .IN2(n73), .QN(n79) );
  NAND2X0 U75 ( .IN1(n84), .IN2(n85), .QN(n137) );
  NAND2X0 U76 ( .IN1(TxPauseTV[5]), .IN2(n131), .QN(n85) );
  MUX21X1 U77 ( .IN1(n162), .IN2(n86), .S(n50), .Q(n84) );
  NOR2X0 U78 ( .IN1(n87), .IN2(n88), .QN(n86) );
  AO222X1 U79 ( .IN1(MAC[37]), .IN2(n64), .IN3(MAC[5]), .IN4(n67), .IN5(
        MAC[45]), .IN6(n65), .Q(n88) );
  AO221X1 U80 ( .IN1(MAC[29]), .IN2(n70), .IN3(MAC[13]), .IN4(n68), .IN5(n89), 
        .Q(n87) );
  AO22X1 U81 ( .IN1(TxPauseTV[13]), .IN2(n69), .IN3(MAC[21]), .IN4(n73), .Q(
        n89) );
  NAND2X0 U82 ( .IN1(n90), .IN2(n91), .QN(n136) );
  NAND2X0 U83 ( .IN1(TxPauseTV[4]), .IN2(n131), .QN(n91) );
  MUX21X1 U84 ( .IN1(n163), .IN2(n92), .S(n50), .Q(n90) );
  NOR2X0 U85 ( .IN1(n93), .IN2(n94), .QN(n92) );
  AO222X1 U86 ( .IN1(MAC[36]), .IN2(n64), .IN3(MAC[4]), .IN4(n67), .IN5(
        MAC[44]), .IN6(n65), .Q(n94) );
  AO221X1 U87 ( .IN1(MAC[28]), .IN2(n70), .IN3(MAC[12]), .IN4(n68), .IN5(n95), 
        .Q(n93) );
  AO22X1 U88 ( .IN1(TxPauseTV[12]), .IN2(n69), .IN3(MAC[20]), .IN4(n73), .Q(
        n95) );
  AO21X1 U89 ( .IN1(TxPauseTV[3]), .IN2(n131), .IN3(n96), .Q(n135) );
  MUX21X1 U90 ( .IN1(ControlData[3]), .IN2(n97), .S(n50), .Q(n96) );
  NAND4X0 U91 ( .IN1(n98), .IN2(n99), .IN3(n100), .IN4(n101), .QN(n97) );
  AOI221X1 U92 ( .IN1(MAC[35]), .IN2(n64), .IN3(MAC[43]), .IN4(n65), .IN5(n102), .QN(n101) );
  AO22X1 U93 ( .IN1(MAC[3]), .IN2(n67), .IN3(MAC[11]), .IN4(n68), .Q(n102) );
  AOI22X1 U94 ( .IN1(TxPauseTV[11]), .IN2(n69), .IN3(MAC[27]), .IN4(n70), .QN(
        n100) );
  NAND3X0 U95 ( .IN1(n48), .IN2(n3), .IN3(n103), .QN(n99) );
  NAND2X0 U96 ( .IN1(MAC[19]), .IN2(n73), .QN(n98) );
  NAND2X0 U97 ( .IN1(n104), .IN2(n105), .QN(n134) );
  NAND2X0 U98 ( .IN1(TxPauseTV[2]), .IN2(n131), .QN(n105) );
  MUX21X1 U99 ( .IN1(n165), .IN2(n106), .S(n50), .Q(n104) );
  NOR2X0 U100 ( .IN1(n107), .IN2(n108), .QN(n106) );
  AO222X1 U101 ( .IN1(MAC[34]), .IN2(n64), .IN3(MAC[2]), .IN4(n67), .IN5(
        MAC[42]), .IN6(n65), .Q(n108) );
  AO221X1 U102 ( .IN1(MAC[26]), .IN2(n70), .IN3(MAC[10]), .IN4(n68), .IN5(n109), .Q(n107) );
  AO22X1 U103 ( .IN1(TxPauseTV[10]), .IN2(n69), .IN3(MAC[18]), .IN4(n73), .Q(
        n109) );
  AO21X1 U104 ( .IN1(TxPauseTV[1]), .IN2(n131), .IN3(n110), .Q(n133) );
  MUX21X1 U105 ( .IN1(ControlData[1]), .IN2(n111), .S(n50), .Q(n110) );
  NAND4X0 U106 ( .IN1(n112), .IN2(n80), .IN3(n113), .IN4(n114), .QN(n111) );
  AOI221X1 U107 ( .IN1(MAC[33]), .IN2(n64), .IN3(MAC[41]), .IN4(n65), .IN5(
        n115), .QN(n114) );
  AO22X1 U108 ( .IN1(MAC[1]), .IN2(n67), .IN3(MAC[9]), .IN4(n68), .Q(n115) );
  AOI22X1 U109 ( .IN1(TxPauseTV[9]), .IN2(n69), .IN3(MAC[25]), .IN4(n70), .QN(
        n113) );
  INVX0 U110 ( .INP(n74), .ZN(n80) );
  NOR3X0 U111 ( .IN1(n1), .IN2(n48), .IN3(n116), .QN(n74) );
  NAND2X0 U112 ( .IN1(MAC[17]), .IN2(n73), .QN(n112) );
  NAND2X0 U113 ( .IN1(n117), .IN2(n118), .QN(n132) );
  NAND2X0 U114 ( .IN1(TxPauseTV[0]), .IN2(n131), .QN(n118) );
  INVX0 U115 ( .INP(n56), .ZN(n131) );
  MUX21X1 U116 ( .IN1(n167), .IN2(n119), .S(n50), .Q(n117) );
  NOR2X0 U117 ( .IN1(n120), .IN2(n121), .QN(n119) );
  AO221X1 U118 ( .IN1(MAC[32]), .IN2(n64), .IN3(MAC[40]), .IN4(n65), .IN5(n122), .Q(n121) );
  AO22X1 U119 ( .IN1(MAC[0]), .IN2(n67), .IN3(MAC[8]), .IN4(n68), .Q(n122) );
  AND3X1 U120 ( .IN1(n49), .IN2(n2), .IN3(n123), .Q(n68) );
  AND3X1 U121 ( .IN1(n2), .IN2(n4), .IN3(n123), .Q(n67) );
  AND2X1 U122 ( .IN1(n124), .IN2(n49), .Q(n65) );
  AND2X1 U123 ( .IN1(n124), .IN2(n4), .Q(n64) );
  AND3X1 U124 ( .IN1(n46), .IN2(n2), .IN3(n103), .Q(n124) );
  AO221X1 U125 ( .IN1(TxPauseTV[8]), .IN2(n69), .IN3(MAC[24]), .IN4(n70), 
        .IN5(n125), .Q(n120) );
  AO221X1 U126 ( .IN1(n126), .IN2(n127), .IN3(MAC[16]), .IN4(n73), .IN5(n128), 
        .Q(n125) );
  NOR4X0 U127 ( .IN1(n57), .IN2(n2), .IN3(n1), .IN4(n116), .QN(n128) );
  OA21X1 U128 ( .IN1(n42), .IN2(n41), .IN3(DlyCrcEn), .Q(n57) );
  AND3X1 U129 ( .IN1(n48), .IN2(n4), .IN3(n123), .Q(n73) );
  XOR2X1 U130 ( .IN1(n3), .IN2(n48), .Q(n127) );
  AND2X1 U131 ( .IN1(n4), .IN2(n103), .Q(n126) );
  NOR2X0 U132 ( .IN1(n1), .IN2(n130), .QN(n103) );
  AND3X1 U133 ( .IN1(n49), .IN2(n48), .IN3(n123), .Q(n70) );
  NOR3X0 U134 ( .IN1(n5), .IN2(n46), .IN3(n1), .QN(n123) );
  NOR3X0 U135 ( .IN1(n2), .IN2(n45), .IN3(n116), .QN(n69) );
  NAND3X0 U136 ( .IN1(n130), .IN2(n46), .IN3(n49), .QN(n116) );
  NAND2X0 U137 ( .IN1(n172), .IN2(n56), .QN(N31) );
  NAND4X0 U138 ( .IN1(n50), .IN2(n48), .IN3(n76), .IN4(n1), .QN(n56) );
  NOR3X0 U139 ( .IN1(n3), .IN2(n49), .IN3(n5), .QN(n76) );
endmodule


module eth_maccontrol_test_1 ( MTxClk, MRxClk, TxReset, RxReset, TPauseRq, 
        TxDataIn, TxStartFrmIn, TxUsedDataIn, TxEndFrmIn, TxDoneIn, TxAbortIn, 
        RxData, RxValid, RxStartFrm, RxEndFrm, ReceiveEnd, ReceivedPacketGood, 
        ReceivedLengthOK, TxFlow, RxFlow, DlyCrcEn, TxPauseTV, MAC, PadIn, 
        PadOut, CrcEnIn, CrcEnOut, TxDataOut, TxStartFrmOut, TxEndFrmOut, 
        TxDoneOut, TxAbortOut, TxUsedDataOut, WillSendControlFrame, 
        TxCtrlEndFrm, ReceivedPauseFrm, ControlFrmAddressOK, SetPauseTimer, 
        r_PassAll, RxStatusWriteLatched_sync2, eth_top_data_sourcea_in, 
        eth_top_test_mode_in, eth_top_test_point_11887_in, test_si, test_se );
  input [7:0] TxDataIn;
  input [7:0] RxData;
  input [15:0] TxPauseTV;
  input [47:0] MAC;
  output [7:0] TxDataOut;
  input MTxClk, MRxClk, TxReset, RxReset, TPauseRq, TxStartFrmIn, TxUsedDataIn,
         TxEndFrmIn, TxDoneIn, TxAbortIn, RxValid, RxStartFrm, RxEndFrm,
         ReceiveEnd, ReceivedPacketGood, ReceivedLengthOK, TxFlow, RxFlow,
         DlyCrcEn, PadIn, CrcEnIn, r_PassAll, RxStatusWriteLatched_sync2,
         eth_top_data_sourcea_in, eth_top_test_mode_in,
         eth_top_test_point_11887_in, test_si, test_se;
  output PadOut, CrcEnOut, TxStartFrmOut, TxEndFrmOut, TxDoneOut, TxAbortOut,
         TxUsedDataOut, WillSendControlFrame, TxCtrlEndFrm, ReceivedPauseFrm,
         ControlFrmAddressOK, SetPauseTimer;
  wire   TxUsedDataOutDetected, TxAbortInLatched, TxDoneInLatched, BlockTxDone,
         CtrlMux, TxCtrlStartFrm, Pause, SendingCtrlFrm, n9, n28, n25, n29,
         n30, n14, n15, n1, n2, n3, n4, n5, n6, n7, n8, n10, n11, n12, n13,
         n16;
  wire   [7:0] ControlData;

  SDFFARX1 TxUsedDataOutDetected_reg ( .D(n28), .SI(TxDoneInLatched), .SE(
        test_se), .CLK(MTxClk), .RSTB(n16), .Q(TxUsedDataOutDetected), .QN(n9)
         );
  SDFFARX1 TxAbortInLatched_reg ( .D(TxAbortIn), .SI(n29), .SE(test_se), .CLK(
        MTxClk), .RSTB(n16), .Q(TxAbortInLatched) );
  SDFFARX1 TxDoneInLatched_reg ( .D(TxDoneIn), .SI(TxAbortInLatched), .SE(
        test_se), .CLK(MTxClk), .RSTB(n16), .Q(TxDoneInLatched) );
  SDFFARX1 MuxedAbort_reg ( .D(n14), .SI(test_si), .SE(test_se), .CLK(MTxClk), 
        .RSTB(n16), .Q(n30), .QN(n13) );
  SDFFARX1 MuxedDone_reg ( .D(n15), .SI(n30), .SE(test_se), .CLK(MTxClk), 
        .RSTB(n16), .Q(n29), .QN(n12) );
  eth_receivecontrol_test_1 receivecontrol1 ( .MTxClk(MTxClk), .MRxClk(MRxClk), 
        .TxReset(TxReset), .RxReset(RxReset), .RxData(RxData), .RxValid(
        RxValid), .RxStartFrm(RxStartFrm), .RxEndFrm(RxEndFrm), .RxFlow(RxFlow), .ReceiveEnd(ReceiveEnd), .MAC(MAC), .DlyCrcEn(DlyCrcEn), .TxDoneIn(TxDoneIn), 
        .TxAbortIn(TxAbortIn), .TxStartFrmOut(TxStartFrmOut), 
        .ReceivedLengthOK(ReceivedLengthOK), .ReceivedPacketGood(
        ReceivedPacketGood), .TxUsedDataOutDetected(TxUsedDataOutDetected), 
        .Pause(Pause), .ReceivedPauseFrm(ReceivedPauseFrm), .AddressOK(
        ControlFrmAddressOK), .RxStatusWriteLatched_sync2(
        RxStatusWriteLatched_sync2), .r_PassAll(r_PassAll), .SetPauseTimer(
        SetPauseTimer), .eth_top_data_sourcea_in(eth_top_data_sourcea_in), 
        .eth_top_test_mode_in(eth_top_test_mode_in), 
        .eth_top_test_point_11887_in(eth_top_test_point_11887_in), .test_so(
        n25), .test_se(test_se) );
  eth_transmitcontrol_test_1 transmitcontrol1 ( .MTxClk(MTxClk), .TxReset(
        TxReset), .TxUsedDataIn(TxUsedDataIn), .TxUsedDataOut(TxUsedDataOut), 
        .TxDoneIn(TxDoneIn), .TxAbortIn(TxAbortIn), .TxStartFrmIn(TxStartFrmIn), .TPauseRq(TPauseRq), .TxUsedDataOutDetected(TxUsedDataOutDetected), .TxFlow(
        TxFlow), .DlyCrcEn(DlyCrcEn), .TxPauseTV(TxPauseTV), .MAC(MAC), 
        .TxCtrlStartFrm(TxCtrlStartFrm), .TxCtrlEndFrm(TxCtrlEndFrm), 
        .SendingCtrlFrm(SendingCtrlFrm), .CtrlMux(CtrlMux), .ControlData(
        ControlData), .WillSendControlFrame(WillSendControlFrame), 
        .BlockTxDone(BlockTxDone), .eth_top_test_point_11887_in(
        eth_top_test_point_11887_in), .test_si(n25), .test_se(test_se) );
  INVX0 U3 ( .INP(eth_top_test_point_11887_in), .ZN(n16) );
  NOR3X0 U4 ( .IN1(n1), .IN2(TxDoneIn), .IN3(TxAbortIn), .QN(n28) );
  NOR2X0 U5 ( .IN1(TxUsedDataOut), .IN2(TxUsedDataOutDetected), .QN(n1) );
  OA21X1 U6 ( .IN1(n2), .IN2(n29), .IN3(n3), .Q(n15) );
  NOR3X0 U7 ( .IN1(TxDoneInLatched), .IN2(n9), .IN3(n4), .QN(n2) );
  OA21X1 U8 ( .IN1(n5), .IN2(n30), .IN3(n3), .Q(n14) );
  NOR3X0 U9 ( .IN1(TxAbortInLatched), .IN2(n9), .IN3(n6), .QN(n5) );
  NOR2X0 U10 ( .IN1(n7), .IN2(CtrlMux), .QN(TxUsedDataOut) );
  INVX0 U11 ( .INP(TxUsedDataIn), .ZN(n7) );
  MUX21X1 U12 ( .IN1(n8), .IN2(TxCtrlStartFrm), .S(CtrlMux), .Q(TxStartFrmOut)
         );
  NOR2X0 U13 ( .IN1(Pause), .IN2(n3), .QN(n8) );
  INVX0 U14 ( .INP(TxStartFrmIn), .ZN(n3) );
  MUX21X1 U15 ( .IN1(TxEndFrmIn), .IN2(TxCtrlEndFrm), .S(CtrlMux), .Q(
        TxEndFrmOut) );
  NOR3X0 U16 ( .IN1(n10), .IN2(TxStartFrmIn), .IN3(BlockTxDone), .QN(TxDoneOut) );
  MUX21X1 U17 ( .IN1(n4), .IN2(n12), .S(CtrlMux), .Q(n10) );
  INVX0 U18 ( .INP(TxDoneIn), .ZN(n4) );
  MUX21X1 U19 ( .IN1(TxDataIn[7]), .IN2(ControlData[7]), .S(CtrlMux), .Q(
        TxDataOut[7]) );
  MUX21X1 U20 ( .IN1(TxDataIn[6]), .IN2(ControlData[6]), .S(CtrlMux), .Q(
        TxDataOut[6]) );
  MUX21X1 U21 ( .IN1(TxDataIn[5]), .IN2(ControlData[5]), .S(CtrlMux), .Q(
        TxDataOut[5]) );
  MUX21X1 U22 ( .IN1(TxDataIn[4]), .IN2(ControlData[4]), .S(CtrlMux), .Q(
        TxDataOut[4]) );
  MUX21X1 U23 ( .IN1(TxDataIn[3]), .IN2(ControlData[3]), .S(CtrlMux), .Q(
        TxDataOut[3]) );
  MUX21X1 U24 ( .IN1(TxDataIn[2]), .IN2(ControlData[2]), .S(CtrlMux), .Q(
        TxDataOut[2]) );
  MUX21X1 U25 ( .IN1(TxDataIn[1]), .IN2(ControlData[1]), .S(CtrlMux), .Q(
        TxDataOut[1]) );
  MUX21X1 U26 ( .IN1(TxDataIn[0]), .IN2(ControlData[0]), .S(CtrlMux), .Q(
        TxDataOut[0]) );
  NOR3X0 U27 ( .IN1(n11), .IN2(TxStartFrmIn), .IN3(BlockTxDone), .QN(
        TxAbortOut) );
  MUX21X1 U28 ( .IN1(n6), .IN2(n13), .S(CtrlMux), .Q(n11) );
  INVX0 U29 ( .INP(TxAbortIn), .ZN(n6) );
  OR2X1 U30 ( .IN1(PadIn), .IN2(SendingCtrlFrm), .Q(PadOut) );
  OR2X1 U31 ( .IN1(CrcEnIn), .IN2(SendingCtrlFrm), .Q(CrcEnOut) );
endmodule


module eth_txcounters_DW01_inc_0 ( A, SUM );
  input [15:0] A;
  output [15:0] SUM;

  wire   [15:2] carry;

  HADDX1 U1_1_14 ( .A0(A[14]), .B0(carry[14]), .C1(carry[15]), .SO(SUM[14]) );
  HADDX1 U1_1_13 ( .A0(A[13]), .B0(carry[13]), .C1(carry[14]), .SO(SUM[13]) );
  HADDX1 U1_1_12 ( .A0(A[12]), .B0(carry[12]), .C1(carry[13]), .SO(SUM[12]) );
  HADDX1 U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1 U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1 U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1 U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  XOR2X1 U2 ( .IN1(carry[15]), .IN2(A[15]), .Q(SUM[15]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module eth_txcounters_DW01_dec_0 ( A, SUM );
  input [18:0] A;
  output [18:0] SUM;
  wire   n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44;

  AO21X1 U16 ( .IN1(A[9]), .IN2(n38), .IN3(n16), .Q(SUM[9]) );
  AO21X1 U17 ( .IN1(A[8]), .IN2(n39), .IN3(n17), .Q(SUM[8]) );
  AO21X1 U18 ( .IN1(A[7]), .IN2(n40), .IN3(n18), .Q(SUM[7]) );
  AO21X1 U19 ( .IN1(A[6]), .IN2(n41), .IN3(n19), .Q(SUM[6]) );
  AO21X1 U20 ( .IN1(A[5]), .IN2(n42), .IN3(n20), .Q(SUM[5]) );
  AO21X1 U21 ( .IN1(A[4]), .IN2(n43), .IN3(n21), .Q(SUM[4]) );
  AO21X1 U22 ( .IN1(A[3]), .IN2(n44), .IN3(n22), .Q(SUM[3]) );
  AO21X1 U23 ( .IN1(A[2]), .IN2(A[1]), .IN3(n23), .Q(SUM[2]) );
  OR2X1 U24 ( .IN1(A[18]), .IN2(n24), .Q(SUM[18]) );
  XOR2X1 U25 ( .IN1(A[18]), .IN2(n24), .Q(SUM[17]) );
  AO21X1 U26 ( .IN1(A[16]), .IN2(n31), .IN3(n24), .Q(SUM[16]) );
  AO21X1 U28 ( .IN1(A[15]), .IN2(n32), .IN3(n25), .Q(SUM[15]) );
  AO21X1 U30 ( .IN1(A[14]), .IN2(n33), .IN3(n26), .Q(SUM[14]) );
  AO21X1 U32 ( .IN1(A[13]), .IN2(n34), .IN3(n27), .Q(SUM[13]) );
  AO21X1 U34 ( .IN1(A[12]), .IN2(n35), .IN3(n28), .Q(SUM[12]) );
  AO21X1 U36 ( .IN1(A[11]), .IN2(n36), .IN3(n29), .Q(SUM[11]) );
  AO21X1 U38 ( .IN1(A[10]), .IN2(n37), .IN3(n30), .Q(SUM[10]) );
  INVX0 U1 ( .INP(n16), .ZN(n37) );
  NOR2X0 U2 ( .IN1(n38), .IN2(A[9]), .QN(n16) );
  INVX0 U3 ( .INP(n22), .ZN(n43) );
  INVX0 U4 ( .INP(n30), .ZN(n36) );
  INVX0 U5 ( .INP(n17), .ZN(n38) );
  INVX0 U6 ( .INP(n25), .ZN(n31) );
  INVX0 U7 ( .INP(n21), .ZN(n42) );
  INVX0 U8 ( .INP(n18), .ZN(n39) );
  INVX0 U9 ( .INP(n20), .ZN(n41) );
  INVX0 U10 ( .INP(n19), .ZN(n40) );
  INVX0 U11 ( .INP(n29), .ZN(n35) );
  INVX0 U12 ( .INP(n27), .ZN(n33) );
  INVX0 U13 ( .INP(n28), .ZN(n34) );
  INVX0 U14 ( .INP(n26), .ZN(n32) );
  NOR2X0 U15 ( .IN1(n44), .IN2(A[3]), .QN(n22) );
  NOR2X0 U27 ( .IN1(n31), .IN2(A[16]), .QN(n24) );
  NOR2X0 U29 ( .IN1(n37), .IN2(A[10]), .QN(n30) );
  NOR2X0 U31 ( .IN1(n39), .IN2(A[8]), .QN(n17) );
  NOR2X0 U33 ( .IN1(n32), .IN2(A[15]), .QN(n25) );
  NOR2X0 U35 ( .IN1(n43), .IN2(A[4]), .QN(n21) );
  NOR2X0 U37 ( .IN1(n41), .IN2(A[6]), .QN(n19) );
  NOR2X0 U39 ( .IN1(n40), .IN2(A[7]), .QN(n18) );
  NOR2X0 U40 ( .IN1(n36), .IN2(A[11]), .QN(n29) );
  NOR2X0 U41 ( .IN1(n35), .IN2(A[12]), .QN(n28) );
  NOR2X0 U42 ( .IN1(n34), .IN2(A[13]), .QN(n27) );
  NOR2X0 U43 ( .IN1(n33), .IN2(A[14]), .QN(n26) );
  NOR2X0 U44 ( .IN1(n42), .IN2(A[5]), .QN(n20) );
  INVX0 U45 ( .INP(n23), .ZN(n44) );
  NOR2X0 U46 ( .IN1(A[2]), .IN2(A[1]), .QN(n23) );
  INVX0 U47 ( .INP(A[1]), .ZN(SUM[1]) );
endmodule


module eth_txcounters_DW01_inc_1 ( A, SUM );
  input [15:0] A;
  output [15:0] SUM;

  wire   [15:2] carry;

  HADDX1 U1_1_14 ( .A0(A[14]), .B0(carry[14]), .C1(carry[15]), .SO(SUM[14]) );
  HADDX1 U1_1_13 ( .A0(A[13]), .B0(carry[13]), .C1(carry[14]), .SO(SUM[13]) );
  HADDX1 U1_1_12 ( .A0(A[12]), .B0(carry[12]), .C1(carry[13]), .SO(SUM[12]) );
  HADDX1 U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1 U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1 U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1 U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  XOR2X1 U2 ( .IN1(carry[15]), .IN2(A[15]), .Q(SUM[15]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module eth_txcounters_test_1 ( StatePreamble, StateIPG, StateData, StatePAD, 
        StateFCS, StateJam, StateBackOff, StateDefer, StateIdle, StartDefer, 
        StartIPG, StartFCS, StartJam, StartBackoff, TxStartFrm, MTxClk, Reset, 
        MinFL, MaxFL, HugEn, ExDfrEn, PacketFinished_q, DlyCrcEn, StateSFD, 
        ByteCnt, NibCnt, ExcessiveDefer, NibCntEq7, NibCntEq15, MaxFrame, 
        NibbleMinFl, DlyCrcCnt, eth_top_test_point_11887_in, test_si, test_se
 );
  input [1:0] StateData;
  input [15:0] MinFL;
  input [15:0] MaxFL;
  output [15:0] ByteCnt;
  output [15:0] NibCnt;
  output [2:0] DlyCrcCnt;
  input StatePreamble, StateIPG, StatePAD, StateFCS, StateJam, StateBackOff,
         StateDefer, StateIdle, StartDefer, StartIPG, StartFCS, StartJam,
         StartBackoff, TxStartFrm, MTxClk, Reset, HugEn, ExDfrEn,
         PacketFinished_q, DlyCrcEn, StateSFD, eth_top_test_point_11887_in,
         test_si, test_se;
  output ExcessiveDefer, NibCntEq7, NibCntEq15, MaxFrame, NibbleMinFl;
  wire   N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20,
         N21, N41, N42, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54,
         N55, N56, N57, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69,
         N70, N71, N72, N73, N74, N75, N76, N79, N80, N81, N82, N83, N84, N85,
         N86, N87, N88, N89, N90, N91, N92, N93, N94, n52, n53, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n219, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n151;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign N41 = MinFL[0];
  assign N42 = MinFL[1];

  SDFFARX1 \NibCnt_reg[0]  ( .D(n131), .SI(DlyCrcCnt[2]), .SE(test_se), .CLK(
        MTxClk), .RSTB(n3), .Q(NibCnt[0]), .QN(n215) );
  SDFFARX1 \NibCnt_reg[15]  ( .D(n116), .SI(NibCnt[14]), .SE(test_se), .CLK(
        MTxClk), .RSTB(n2), .Q(NibCnt[15]), .QN(n200) );
  SDFFARX1 \NibCnt_reg[1]  ( .D(n129), .SI(NibCnt[0]), .SE(test_se), .CLK(
        MTxClk), .RSTB(n2), .Q(NibCnt[1]), .QN(n201) );
  SDFFARX1 \NibCnt_reg[2]  ( .D(n128), .SI(NibCnt[1]), .SE(test_se), .CLK(
        MTxClk), .RSTB(n3), .Q(NibCnt[2]), .QN(n202) );
  SDFFARX1 \NibCnt_reg[3]  ( .D(n130), .SI(NibCnt[2]), .SE(test_se), .CLK(
        MTxClk), .RSTB(n2), .Q(NibCnt[3]), .QN(n203) );
  SDFFARX1 \NibCnt_reg[4]  ( .D(n127), .SI(NibCnt[3]), .SE(test_se), .CLK(
        MTxClk), .RSTB(n3), .Q(NibCnt[4]), .QN(n204) );
  SDFFARX1 \NibCnt_reg[5]  ( .D(n126), .SI(NibCnt[4]), .SE(test_se), .CLK(
        MTxClk), .RSTB(n2), .Q(NibCnt[5]), .QN(n205) );
  SDFFARX1 \NibCnt_reg[6]  ( .D(n125), .SI(NibCnt[5]), .SE(test_se), .CLK(
        MTxClk), .RSTB(n3), .Q(NibCnt[6]), .QN(n206) );
  SDFFARX1 \NibCnt_reg[7]  ( .D(n124), .SI(NibCnt[6]), .SE(test_se), .CLK(
        MTxClk), .RSTB(n2), .Q(NibCnt[7]), .QN(n207) );
  SDFFARX1 \NibCnt_reg[8]  ( .D(n123), .SI(NibCnt[7]), .SE(test_se), .CLK(
        MTxClk), .RSTB(n3), .Q(NibCnt[8]), .QN(n208) );
  SDFFARX1 \NibCnt_reg[9]  ( .D(n122), .SI(NibCnt[8]), .SE(test_se), .CLK(
        MTxClk), .RSTB(n2), .Q(NibCnt[9]), .QN(n209) );
  SDFFARX1 \NibCnt_reg[10]  ( .D(n121), .SI(NibCnt[9]), .SE(test_se), .CLK(
        MTxClk), .RSTB(n3), .Q(NibCnt[10]), .QN(n210) );
  SDFFARX1 \NibCnt_reg[11]  ( .D(n120), .SI(NibCnt[10]), .SE(test_se), .CLK(
        MTxClk), .RSTB(n2), .Q(NibCnt[11]), .QN(n211) );
  SDFFARX1 \NibCnt_reg[12]  ( .D(n119), .SI(NibCnt[11]), .SE(test_se), .CLK(
        MTxClk), .RSTB(n3), .Q(NibCnt[12]), .QN(n212) );
  SDFFARX1 \NibCnt_reg[13]  ( .D(n118), .SI(NibCnt[12]), .SE(test_se), .CLK(
        MTxClk), .RSTB(n2), .Q(NibCnt[13]), .QN(n213) );
  SDFFARX1 \NibCnt_reg[14]  ( .D(n117), .SI(NibCnt[13]), .SE(test_se), .CLK(
        MTxClk), .RSTB(n3), .Q(NibCnt[14]), .QN(n214) );
  SDFFARX1 \ByteCnt_reg[0]  ( .D(n115), .SI(test_si), .SE(test_se), .CLK(
        MTxClk), .RSTB(n3), .Q(ByteCnt[0]), .QN(n198) );
  SDFFARX1 \ByteCnt_reg[14]  ( .D(n100), .SI(ByteCnt[13]), .SE(test_se), .CLK(
        MTxClk), .RSTB(n3), .Q(ByteCnt[14]), .QN(n188) );
  SDFFARX1 \ByteCnt_reg[1]  ( .D(n113), .SI(ByteCnt[0]), .SE(test_se), .CLK(
        MTxClk), .RSTB(n2), .Q(ByteCnt[1]) );
  SDFFARX1 \ByteCnt_reg[2]  ( .D(n112), .SI(ByteCnt[1]), .SE(test_se), .CLK(
        MTxClk), .RSTB(n3), .Q(ByteCnt[2]), .QN(n199) );
  SDFFARX1 \ByteCnt_reg[3]  ( .D(n111), .SI(ByteCnt[2]), .SE(test_se), .CLK(
        MTxClk), .RSTB(n2), .Q(ByteCnt[3]), .QN(n193) );
  SDFFARX1 \ByteCnt_reg[4]  ( .D(n110), .SI(ByteCnt[3]), .SE(test_se), .CLK(
        MTxClk), .RSTB(n3), .Q(ByteCnt[4]), .QN(n194) );
  SDFFARX1 \ByteCnt_reg[5]  ( .D(n109), .SI(ByteCnt[4]), .SE(test_se), .CLK(
        MTxClk), .RSTB(n2), .Q(ByteCnt[5]), .QN(n195) );
  SDFFARX1 \ByteCnt_reg[6]  ( .D(n108), .SI(ByteCnt[5]), .SE(test_se), .CLK(
        MTxClk), .RSTB(n3), .Q(ByteCnt[6]), .QN(n196) );
  SDFFARX1 \ByteCnt_reg[7]  ( .D(n107), .SI(ByteCnt[6]), .SE(test_se), .CLK(
        MTxClk), .RSTB(n2), .Q(ByteCnt[7]), .QN(n189) );
  SDFFARX1 \ByteCnt_reg[8]  ( .D(n106), .SI(ByteCnt[7]), .SE(test_se), .CLK(
        MTxClk), .RSTB(n3), .Q(ByteCnt[8]), .QN(n190) );
  SDFFARX1 \ByteCnt_reg[9]  ( .D(n105), .SI(ByteCnt[8]), .SE(test_se), .CLK(
        MTxClk), .RSTB(n2), .Q(ByteCnt[9]), .QN(n191) );
  SDFFARX1 \ByteCnt_reg[10]  ( .D(n104), .SI(ByteCnt[9]), .SE(test_se), .CLK(
        MTxClk), .RSTB(n3), .Q(ByteCnt[10]), .QN(n192) );
  SDFFARX1 \ByteCnt_reg[11]  ( .D(n103), .SI(ByteCnt[10]), .SE(test_se), .CLK(
        MTxClk), .RSTB(n2), .Q(ByteCnt[11]), .QN(n185) );
  SDFFARX1 \ByteCnt_reg[12]  ( .D(n102), .SI(ByteCnt[11]), .SE(test_se), .CLK(
        MTxClk), .RSTB(n3), .Q(ByteCnt[12]), .QN(n186) );
  SDFFARX1 \ByteCnt_reg[13]  ( .D(n101), .SI(ByteCnt[12]), .SE(test_se), .CLK(
        MTxClk), .RSTB(n2), .Q(ByteCnt[13]), .QN(n187) );
  SDFFARX1 \ByteCnt_reg[15]  ( .D(n114), .SI(ByteCnt[14]), .SE(test_se), .CLK(
        MTxClk), .RSTB(n2), .Q(ByteCnt[15]), .QN(n219) );
  SDFFARX1 \DlyCrcCnt_reg[0]  ( .D(n99), .SI(ByteCnt[15]), .SE(test_se), .CLK(
        MTxClk), .RSTB(n2), .Q(DlyCrcCnt[0]), .QN(n53) );
  SDFFARX1 \DlyCrcCnt_reg[2]  ( .D(n98), .SI(DlyCrcCnt[1]), .SE(test_se), 
        .CLK(MTxClk), .RSTB(n2), .Q(DlyCrcCnt[2]), .QN(n184) );
  SDFFARX1 \DlyCrcCnt_reg[1]  ( .D(n97), .SI(DlyCrcCnt[0]), .SE(test_se), 
        .CLK(MTxClk), .RSTB(n3), .Q(DlyCrcCnt[1]), .QN(n52) );
  eth_txcounters_DW01_inc_0 add_197 ( .A(ByteCnt), .SUM({N94, N93, N92, N91, 
        N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79}) );
  eth_txcounters_DW01_dec_0 sub_173_2 ( .A({N57, N57, N56, N55, N54, N53, N52, 
        N51, N50, N49, N48, N47, N46, N45, N44, n151, N42, N41, 1'b0}), .SUM({
        N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, 
        N62, N61, N60, N59, SYNOPSYS_UNCONNECTED__0}) );
  eth_txcounters_DW01_inc_1 add_165 ( .A(NibCnt), .SUM({N21, N20, N19, N18, 
        N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6}) );
  INVX0 U4 ( .INP(eth_top_test_point_11887_in), .ZN(n2) );
  INVX0 U5 ( .INP(eth_top_test_point_11887_in), .ZN(n3) );
  INVX0 U6 ( .INP(n4), .ZN(ExcessiveDefer) );
  INVX0 U7 ( .INP(MinFL[2]), .ZN(n151) );
  MUX21X1 U8 ( .IN1(n5), .IN2(n6), .S(n53), .Q(n99) );
  NOR2X0 U9 ( .IN1(n6), .IN2(n7), .QN(n5) );
  MUX21X1 U10 ( .IN1(n8), .IN2(n9), .S(n184), .Q(n98) );
  NOR3X0 U11 ( .IN1(n10), .IN2(n53), .IN3(n52), .QN(n9) );
  AO21X1 U12 ( .IN1(n6), .IN2(n52), .IN3(n11), .Q(n8) );
  INVX0 U13 ( .INP(n10), .ZN(n6) );
  MUX21X1 U14 ( .IN1(n11), .IN2(n12), .S(n52), .Q(n97) );
  NOR2X0 U15 ( .IN1(n53), .IN2(n10), .QN(n12) );
  MUX21X1 U16 ( .IN1(n53), .IN2(n13), .S(n10), .Q(n11) );
  NAND3X0 U17 ( .IN1(n13), .IN2(n14), .IN3(DlyCrcEn), .QN(n10) );
  AO21X1 U18 ( .IN1(StateData[1]), .IN2(n15), .IN3(StateSFD), .Q(n14) );
  NAND2X0 U19 ( .IN1(n53), .IN2(n52), .QN(n15) );
  INVX0 U20 ( .INP(n7), .ZN(n13) );
  NAND3X0 U21 ( .IN1(n16), .IN2(n17), .IN3(n18), .QN(n7) );
  NAND4X0 U22 ( .IN1(n53), .IN2(n52), .IN3(StateData[1]), .IN4(DlyCrcCnt[2]), 
        .QN(n18) );
  INVX0 U23 ( .INP(StartJam), .ZN(n17) );
  AO22X1 U24 ( .IN1(N6), .IN2(n19), .IN3(n20), .IN4(NibCnt[0]), .Q(n131) );
  AO22X1 U25 ( .IN1(N9), .IN2(n19), .IN3(n20), .IN4(NibCnt[3]), .Q(n130) );
  AO22X1 U26 ( .IN1(N7), .IN2(n19), .IN3(n20), .IN4(NibCnt[1]), .Q(n129) );
  AO22X1 U27 ( .IN1(N8), .IN2(n19), .IN3(n20), .IN4(NibCnt[2]), .Q(n128) );
  AO22X1 U28 ( .IN1(N10), .IN2(n19), .IN3(n20), .IN4(NibCnt[4]), .Q(n127) );
  AO22X1 U29 ( .IN1(N11), .IN2(n19), .IN3(n20), .IN4(NibCnt[5]), .Q(n126) );
  AO22X1 U30 ( .IN1(N12), .IN2(n19), .IN3(n20), .IN4(NibCnt[6]), .Q(n125) );
  AO22X1 U31 ( .IN1(N13), .IN2(n19), .IN3(n20), .IN4(NibCnt[7]), .Q(n124) );
  AO22X1 U32 ( .IN1(N14), .IN2(n19), .IN3(n20), .IN4(NibCnt[8]), .Q(n123) );
  AO22X1 U33 ( .IN1(N15), .IN2(n19), .IN3(n20), .IN4(NibCnt[9]), .Q(n122) );
  AO22X1 U34 ( .IN1(N16), .IN2(n19), .IN3(n20), .IN4(NibCnt[10]), .Q(n121) );
  AO22X1 U35 ( .IN1(N17), .IN2(n19), .IN3(n20), .IN4(NibCnt[11]), .Q(n120) );
  AO22X1 U36 ( .IN1(N18), .IN2(n19), .IN3(n20), .IN4(NibCnt[12]), .Q(n119) );
  AO22X1 U37 ( .IN1(N19), .IN2(n19), .IN3(n20), .IN4(NibCnt[13]), .Q(n118) );
  AO22X1 U38 ( .IN1(N20), .IN2(n19), .IN3(n20), .IN4(NibCnt[14]), .Q(n117) );
  AO22X1 U39 ( .IN1(N21), .IN2(n19), .IN3(n20), .IN4(NibCnt[15]), .Q(n116) );
  AND2X1 U40 ( .IN1(n21), .IN2(n22), .Q(n20) );
  INVX0 U41 ( .INP(n22), .ZN(n19) );
  NAND2X0 U42 ( .IN1(n21), .IN2(n23), .QN(n22) );
  NAND4X0 U43 ( .IN1(n24), .IN2(n25), .IN3(n26), .IN4(n27), .QN(n23) );
  NOR4X0 U44 ( .IN1(StatePreamble), .IN2(StateJam), .IN3(StateIPG), .IN4(
        StateData[1]), .QN(n27) );
  NOR2X0 U45 ( .IN1(StateData[0]), .IN2(StateBackOff), .QN(n26) );
  NAND3X0 U46 ( .IN1(StateDefer), .IN2(n4), .IN3(TxStartFrm), .QN(n25) );
  NOR4X0 U47 ( .IN1(StartDefer), .IN2(n28), .IN3(n29), .IN4(n30), .QN(n21) );
  OR4X1 U48 ( .IN1(StartIPG), .IN2(StartFCS), .IN3(StateIdle), .IN4(StartJam), 
        .Q(n30) );
  AO22X1 U49 ( .IN1(StatePreamble), .IN2(NibCntEq15), .IN3(StateJam), .IN4(
        NibCntEq7), .Q(n29) );
  NOR3X0 U50 ( .IN1(n31), .IN2(TxStartFrm), .IN3(n4), .QN(n28) );
  NAND4X0 U51 ( .IN1(n32), .IN2(n203), .IN3(n33), .IN4(n34), .QN(n4) );
  NOR4X0 U52 ( .IN1(n35), .IN2(n204), .IN3(n207), .IN4(n205), .QN(n34) );
  NAND4X0 U53 ( .IN1(NibCnt[8]), .IN2(NibCnt[9]), .IN3(NibCnt[10]), .IN4(
        NibCnt[12]), .QN(n35) );
  AND3X1 U54 ( .IN1(n211), .IN2(n206), .IN3(n213), .Q(n33) );
  NOR2X0 U55 ( .IN1(ExDfrEn), .IN2(n36), .QN(n32) );
  INVX0 U56 ( .INP(StateDefer), .ZN(n31) );
  AO22X1 U57 ( .IN1(N79), .IN2(n37), .IN3(n38), .IN4(ByteCnt[0]), .Q(n115) );
  AO22X1 U58 ( .IN1(N94), .IN2(n37), .IN3(n38), .IN4(ByteCnt[15]), .Q(n114) );
  AO22X1 U59 ( .IN1(N80), .IN2(n37), .IN3(n38), .IN4(ByteCnt[1]), .Q(n113) );
  AO22X1 U60 ( .IN1(N81), .IN2(n37), .IN3(n38), .IN4(ByteCnt[2]), .Q(n112) );
  AO22X1 U61 ( .IN1(N82), .IN2(n37), .IN3(n38), .IN4(ByteCnt[3]), .Q(n111) );
  AO22X1 U62 ( .IN1(N83), .IN2(n37), .IN3(n38), .IN4(ByteCnt[4]), .Q(n110) );
  AO22X1 U63 ( .IN1(N84), .IN2(n37), .IN3(n38), .IN4(ByteCnt[5]), .Q(n109) );
  AO22X1 U64 ( .IN1(N85), .IN2(n37), .IN3(n38), .IN4(ByteCnt[6]), .Q(n108) );
  AO22X1 U65 ( .IN1(N86), .IN2(n37), .IN3(n38), .IN4(ByteCnt[7]), .Q(n107) );
  AO22X1 U66 ( .IN1(N87), .IN2(n37), .IN3(n38), .IN4(ByteCnt[8]), .Q(n106) );
  AO22X1 U67 ( .IN1(N88), .IN2(n37), .IN3(n38), .IN4(ByteCnt[9]), .Q(n105) );
  AO22X1 U68 ( .IN1(N89), .IN2(n37), .IN3(n38), .IN4(ByteCnt[10]), .Q(n104) );
  AO22X1 U69 ( .IN1(N90), .IN2(n37), .IN3(n38), .IN4(ByteCnt[11]), .Q(n103) );
  AO22X1 U70 ( .IN1(N91), .IN2(n37), .IN3(n38), .IN4(ByteCnt[12]), .Q(n102) );
  AO22X1 U71 ( .IN1(N92), .IN2(n37), .IN3(n38), .IN4(ByteCnt[13]), .Q(n101) );
  AO22X1 U72 ( .IN1(N93), .IN2(n37), .IN3(n38), .IN4(ByteCnt[14]), .Q(n100) );
  AND4X1 U73 ( .IN1(n39), .IN2(n40), .IN3(n16), .IN4(n41), .Q(n38) );
  INVX0 U74 ( .INP(n39), .ZN(n37) );
  NAND4X0 U75 ( .IN1(n42), .IN2(n40), .IN3(n41), .IN4(n16), .QN(n39) );
  INVX0 U76 ( .INP(PacketFinished_q), .ZN(n16) );
  INVX0 U77 ( .INP(StartBackoff), .ZN(n41) );
  NAND2X0 U78 ( .IN1(StateIdle), .IN2(TxStartFrm), .QN(n40) );
  OAI21X1 U79 ( .IN1(n43), .IN2(n44), .IN3(n45), .QN(n42) );
  NAND4X0 U80 ( .IN1(StateBackOff), .IN2(NibCntEq15), .IN3(n46), .IN4(
        NibCnt[4]), .QN(n45) );
  NOR2X0 U81 ( .IN1(n206), .IN2(n205), .QN(n46) );
  OA21X1 U82 ( .IN1(n215), .IN2(n24), .IN3(n47), .Q(n44) );
  INVX0 U83 ( .INP(StateData[1]), .ZN(n47) );
  NOR2X0 U84 ( .IN1(StateFCS), .IN2(StatePAD), .QN(n24) );
  NOR4X0 U85 ( .IN1(n48), .IN2(n49), .IN3(n50), .IN4(n51), .QN(n43) );
  NAND4X0 U86 ( .IN1(ByteCnt[11]), .IN2(ByteCnt[12]), .IN3(ByteCnt[13]), .IN4(
        ByteCnt[14]), .QN(n51) );
  NAND4X0 U87 ( .IN1(ByteCnt[7]), .IN2(ByteCnt[8]), .IN3(ByteCnt[9]), .IN4(
        ByteCnt[10]), .QN(n50) );
  NAND4X0 U88 ( .IN1(ByteCnt[3]), .IN2(ByteCnt[4]), .IN3(ByteCnt[5]), .IN4(
        ByteCnt[6]), .QN(n49) );
  NAND4X0 U89 ( .IN1(ByteCnt[1]), .IN2(ByteCnt[0]), .IN3(ByteCnt[2]), .IN4(
        ByteCnt[15]), .QN(n48) );
  NOR4X0 U90 ( .IN1(n54), .IN2(N74), .IN3(N76), .IN4(N75), .QN(NibbleMinFl) );
  AO21X1 U91 ( .IN1(n200), .IN2(N73), .IN3(n55), .Q(n54) );
  OA221X1 U92 ( .IN1(N72), .IN2(n214), .IN3(N73), .IN4(n200), .IN5(n56), .Q(
        n55) );
  AO221X1 U93 ( .IN1(N71), .IN2(n213), .IN3(n214), .IN4(N72), .IN5(n57), .Q(
        n56) );
  OA221X1 U94 ( .IN1(N70), .IN2(n212), .IN3(N71), .IN4(n213), .IN5(n58), .Q(
        n57) );
  AO221X1 U95 ( .IN1(N69), .IN2(n211), .IN3(n212), .IN4(N70), .IN5(n59), .Q(
        n58) );
  OA221X1 U96 ( .IN1(N68), .IN2(n210), .IN3(N69), .IN4(n211), .IN5(n60), .Q(
        n59) );
  AO221X1 U97 ( .IN1(n209), .IN2(N67), .IN3(n210), .IN4(N68), .IN5(n61), .Q(
        n60) );
  OA221X1 U98 ( .IN1(N66), .IN2(n208), .IN3(N67), .IN4(n209), .IN5(n62), .Q(
        n61) );
  AO221X1 U99 ( .IN1(n207), .IN2(N65), .IN3(n208), .IN4(N66), .IN5(n63), .Q(
        n62) );
  OA221X1 U100 ( .IN1(N64), .IN2(n206), .IN3(N65), .IN4(n207), .IN5(n64), .Q(
        n63) );
  AO221X1 U101 ( .IN1(n205), .IN2(N63), .IN3(N64), .IN4(n206), .IN5(n65), .Q(
        n64) );
  OA221X1 U102 ( .IN1(N62), .IN2(n204), .IN3(N63), .IN4(n205), .IN5(n66), .Q(
        n65) );
  AO221X1 U103 ( .IN1(N61), .IN2(n203), .IN3(n204), .IN4(N62), .IN5(n67), .Q(
        n66) );
  OA221X1 U104 ( .IN1(N61), .IN2(n203), .IN3(N60), .IN4(n202), .IN5(n68), .Q(
        n67) );
  AO222X1 U105 ( .IN1(n202), .IN2(N60), .IN3(N59), .IN4(n69), .IN5(n215), 
        .IN6(n201), .Q(n68) );
  NOR2X0 U106 ( .IN1(n36), .IN2(n203), .QN(NibCntEq15) );
  INVX0 U107 ( .INP(NibCntEq7), .ZN(n36) );
  NOR2X0 U108 ( .IN1(n69), .IN2(n202), .QN(NibCntEq7) );
  NAND2X0 U109 ( .IN1(NibCnt[0]), .IN2(NibCnt[1]), .QN(n69) );
  AO21X1 U110 ( .IN1(MinFL[15]), .IN2(n70), .IN3(N57), .Q(N56) );
  NOR2X0 U111 ( .IN1(n70), .IN2(MinFL[15]), .QN(N57) );
  INVX0 U112 ( .INP(n71), .ZN(n70) );
  AO21X1 U113 ( .IN1(MinFL[14]), .IN2(n72), .IN3(n71), .Q(N55) );
  NOR2X0 U114 ( .IN1(n72), .IN2(MinFL[14]), .QN(n71) );
  INVX0 U115 ( .INP(n73), .ZN(n72) );
  AO21X1 U116 ( .IN1(MinFL[13]), .IN2(n74), .IN3(n73), .Q(N54) );
  NOR2X0 U117 ( .IN1(n74), .IN2(MinFL[13]), .QN(n73) );
  INVX0 U118 ( .INP(n75), .ZN(n74) );
  AO21X1 U119 ( .IN1(MinFL[12]), .IN2(n76), .IN3(n75), .Q(N53) );
  NOR2X0 U120 ( .IN1(n76), .IN2(MinFL[12]), .QN(n75) );
  INVX0 U121 ( .INP(n77), .ZN(n76) );
  AO21X1 U122 ( .IN1(MinFL[11]), .IN2(n78), .IN3(n77), .Q(N52) );
  NOR2X0 U123 ( .IN1(n78), .IN2(MinFL[11]), .QN(n77) );
  INVX0 U124 ( .INP(n79), .ZN(n78) );
  AO21X1 U125 ( .IN1(MinFL[10]), .IN2(n80), .IN3(n79), .Q(N51) );
  NOR2X0 U126 ( .IN1(n80), .IN2(MinFL[10]), .QN(n79) );
  INVX0 U127 ( .INP(n81), .ZN(n80) );
  AO21X1 U128 ( .IN1(MinFL[9]), .IN2(n82), .IN3(n81), .Q(N50) );
  NOR2X0 U129 ( .IN1(n82), .IN2(MinFL[9]), .QN(n81) );
  NAND2X0 U130 ( .IN1(n82), .IN2(n83), .QN(N49) );
  AO21X1 U131 ( .IN1(n84), .IN2(n85), .IN3(n86), .Q(n83) );
  NAND3X0 U132 ( .IN1(n85), .IN2(n86), .IN3(n84), .QN(n82) );
  INVX0 U133 ( .INP(MinFL[8]), .ZN(n86) );
  INVX0 U134 ( .INP(MinFL[7]), .ZN(n85) );
  XOR2X1 U135 ( .IN1(MinFL[7]), .IN2(n84), .Q(N48) );
  AO21X1 U136 ( .IN1(MinFL[6]), .IN2(n87), .IN3(n84), .Q(N47) );
  NOR2X0 U137 ( .IN1(n87), .IN2(MinFL[6]), .QN(n84) );
  INVX0 U138 ( .INP(n88), .ZN(n87) );
  AO21X1 U139 ( .IN1(MinFL[5]), .IN2(n89), .IN3(n88), .Q(N46) );
  NOR2X0 U140 ( .IN1(n89), .IN2(MinFL[5]), .QN(n88) );
  INVX0 U141 ( .INP(n90), .ZN(n89) );
  AO21X1 U142 ( .IN1(MinFL[4]), .IN2(n91), .IN3(n90), .Q(N45) );
  NOR2X0 U143 ( .IN1(n91), .IN2(MinFL[4]), .QN(n90) );
  INVX0 U144 ( .INP(n92), .ZN(n91) );
  AO21X1 U145 ( .IN1(MinFL[3]), .IN2(MinFL[2]), .IN3(n92), .Q(N44) );
  NOR2X0 U146 ( .IN1(MinFL[3]), .IN2(MinFL[2]), .QN(n92) );
  NOR4X0 U147 ( .IN1(n93), .IN2(n94), .IN3(n95), .IN4(n96), .QN(MaxFrame) );
  NAND4X0 U148 ( .IN1(n132), .IN2(n133), .IN3(n134), .IN4(n135), .QN(n96) );
  XOR2X1 U149 ( .IN1(n185), .IN2(MaxFL[11]), .Q(n135) );
  XOR2X1 U150 ( .IN1(n186), .IN2(MaxFL[12]), .Q(n134) );
  XOR2X1 U151 ( .IN1(n187), .IN2(MaxFL[13]), .Q(n133) );
  XOR2X1 U152 ( .IN1(n219), .IN2(MaxFL[15]), .Q(n132) );
  NAND4X0 U153 ( .IN1(n136), .IN2(n137), .IN3(n138), .IN4(n139), .QN(n95) );
  XOR2X1 U154 ( .IN1(n192), .IN2(MaxFL[10]), .Q(n139) );
  XOR2X1 U155 ( .IN1(n188), .IN2(MaxFL[14]), .Q(n138) );
  XOR2X1 U156 ( .IN1(n189), .IN2(MaxFL[7]), .Q(n137) );
  XOR2X1 U157 ( .IN1(n190), .IN2(MaxFL[8]), .Q(n136) );
  NAND4X0 U158 ( .IN1(n140), .IN2(n141), .IN3(n142), .IN4(n143), .QN(n94) );
  XOR2X1 U159 ( .IN1(n193), .IN2(MaxFL[3]), .Q(n143) );
  XOR2X1 U160 ( .IN1(n194), .IN2(MaxFL[4]), .Q(n142) );
  XOR2X1 U161 ( .IN1(n195), .IN2(MaxFL[5]), .Q(n141) );
  XOR2X1 U162 ( .IN1(n191), .IN2(MaxFL[9]), .Q(n140) );
  NAND4X0 U163 ( .IN1(n144), .IN2(n145), .IN3(n146), .IN4(n147), .QN(n93) );
  XOR2X1 U164 ( .IN1(n198), .IN2(MaxFL[0]), .Q(n147) );
  NOR2X0 U165 ( .IN1(HugEn), .IN2(n148), .QN(n146) );
  XOR2X1 U166 ( .IN1(ByteCnt[1]), .IN2(MaxFL[1]), .Q(n148) );
  XOR2X1 U167 ( .IN1(n199), .IN2(MaxFL[2]), .Q(n145) );
  XOR2X1 U168 ( .IN1(n196), .IN2(MaxFL[6]), .Q(n144) );
endmodule


module eth_txstatem_test_1 ( MTxClk, Reset, ExcessiveDefer, CarrierSense, 
        NibCnt, IPGT, IPGR1, IPGR2, FullD, TxStartFrm, TxEndFrm, TxUnderRun, 
        Collision, UnderRun, StartTxDone, TooBig, NibCntEq7, NibCntEq15, 
        MaxFrame, Pad, CrcEn, NibbleMinFl, RandomEq0, ColWindow, RetryMax, 
        NoBckof, RandomEqByteCnt, StateIdle, StateIPG, StatePreamble, 
        StateData, StatePAD, StateFCS, StateJam, StateJam_q, StateBackOff, 
        StateDefer, StartFCS, StartJam, StartBackoff, StartDefer, 
        DeferIndication, StartPreamble, StartData, StartIPG, 
        eth_top_test_point_11887_in, test_si, test_se );
  input [6:0] NibCnt;
  input [6:0] IPGT;
  input [6:0] IPGR1;
  input [6:0] IPGR2;
  output [1:0] StateData;
  output [1:0] StartData;
  input MTxClk, Reset, ExcessiveDefer, CarrierSense, FullD, TxStartFrm,
         TxEndFrm, TxUnderRun, Collision, UnderRun, StartTxDone, TooBig,
         NibCntEq7, NibCntEq15, MaxFrame, Pad, CrcEn, NibbleMinFl, RandomEq0,
         ColWindow, RetryMax, NoBckof, RandomEqByteCnt,
         eth_top_test_point_11887_in, test_si, test_se;
  output StateIdle, StateIPG, StatePreamble, StatePAD, StateFCS, StateJam,
         StateJam_q, StateBackOff, StateDefer, StartFCS, StartJam,
         StartBackoff, StartDefer, DeferIndication, StartPreamble, StartIPG;
  wire   n24, n26, n27, n28, n69, n70, n71, n72, n73, n74, n75, n76, n77, n12,
         n100, n101, n102, n103, n108, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n25, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n105;

  SDFFARX1 Rule1_reg ( .D(n77), .SI(test_si), .SE(test_se), .CLK(MTxClk), 
        .RSTB(n105), .Q(n100), .QN(n12) );
  SDFFASX1 StateDefer_reg ( .D(n71), .SI(StateData[1]), .SE(test_se), .CLK(
        MTxClk), .SETB(n105), .Q(StateDefer), .QN(n101) );
  SDFFARX1 StateIPG_reg ( .D(n70), .SI(StateFCS), .SE(test_se), .CLK(MTxClk), 
        .RSTB(n105), .Q(StateIPG), .QN(n108) );
  SDFFARX1 StateIdle_reg ( .D(n76), .SI(StateIPG), .SE(test_se), .CLK(MTxClk), 
        .RSTB(n105), .Q(StateIdle), .QN(n103) );
  SDFFARX1 StateFCS_reg ( .D(n75), .SI(StateDefer), .SE(test_se), .CLK(MTxClk), 
        .RSTB(n105), .Q(StateFCS), .QN(n26) );
  SDFFARX1 StateJam_reg ( .D(n72), .SI(StateJam_q), .SE(test_se), .CLK(MTxClk), 
        .RSTB(n105), .Q(StateJam) );
  SDFFARX1 StateJam_q_reg ( .D(StateJam), .SI(StateIdle), .SE(test_se), .CLK(
        MTxClk), .RSTB(n105), .Q(StateJam_q) );
  SDFFARX1 StateBackOff_reg ( .D(n69), .SI(n100), .SE(test_se), .CLK(MTxClk), 
        .RSTB(n105), .Q(StateBackOff) );
  SDFFARX1 StatePreamble_reg ( .D(n74), .SI(StatePAD), .SE(test_se), .CLK(
        MTxClk), .RSTB(n105), .Q(StatePreamble), .QN(n102) );
  SDFFARX1 \StateData_reg[0]  ( .D(StartData[0]), .SI(StateBackOff), .SE(
        test_se), .CLK(MTxClk), .RSTB(n105), .Q(StateData[0]), .QN(n28) );
  SDFFARX1 \StateData_reg[1]  ( .D(StartData[1]), .SI(StateData[0]), .SE(
        test_se), .CLK(MTxClk), .RSTB(n105), .Q(StateData[1]), .QN(n27) );
  SDFFARX1 StatePAD_reg ( .D(n73), .SI(StateJam), .SE(test_se), .CLK(MTxClk), 
        .RSTB(n105), .Q(StatePAD), .QN(n24) );
  INVX0 U3 ( .INP(eth_top_test_point_11887_in), .ZN(n105) );
  NOR3X0 U4 ( .IN1(StateBackOff), .IN2(n1), .IN3(StateIdle), .QN(n77) );
  AND3X1 U5 ( .IN1(n12), .IN2(n2), .IN3(n102), .Q(n1) );
  INVX0 U6 ( .INP(FullD), .ZN(n2) );
  NOR3X0 U7 ( .IN1(n3), .IN2(StartPreamble), .IN3(StartDefer), .QN(n76) );
  NOR2X0 U8 ( .IN1(n4), .IN2(StateIdle), .QN(n3) );
  NOR3X0 U9 ( .IN1(n5), .IN2(StartJam), .IN3(StartDefer), .QN(n75) );
  AND2X1 U10 ( .IN1(n6), .IN2(n26), .Q(n5) );
  NOR3X0 U11 ( .IN1(n7), .IN2(StartJam), .IN3(StartData[0]), .QN(n74) );
  NOR2X0 U12 ( .IN1(StartPreamble), .IN2(StatePreamble), .QN(n7) );
  NOR3X0 U13 ( .IN1(StartFCS), .IN2(StartJam), .IN3(n8), .QN(n73) );
  AND2X1 U14 ( .IN1(n24), .IN2(n9), .Q(n8) );
  NAND4X0 U15 ( .IN1(Pad), .IN2(TxEndFrm), .IN3(n10), .IN4(StateData[1]), .QN(
        n9) );
  INVX0 U16 ( .INP(n6), .ZN(StartFCS) );
  NAND4X0 U17 ( .IN1(CrcEn), .IN2(n11), .IN3(n13), .IN4(n14), .QN(n6) );
  OAI22X1 U18 ( .IN1(n15), .IN2(n27), .IN3(n10), .IN4(n24), .QN(n13) );
  NAND2X0 U19 ( .IN1(Pad), .IN2(n10), .QN(n11) );
  INVX0 U20 ( .INP(NibbleMinFl), .ZN(n10) );
  NOR3X0 U21 ( .IN1(n16), .IN2(StartDefer), .IN3(StartBackoff), .QN(n72) );
  NOR2X0 U22 ( .IN1(StartJam), .IN2(StateJam), .QN(n16) );
  AOI21X1 U23 ( .IN1(n17), .IN2(n101), .IN3(StartIPG), .QN(n71) );
  NOR3X0 U24 ( .IN1(n18), .IN2(StartDefer), .IN3(n4), .QN(n70) );
  AND2X1 U25 ( .IN1(n19), .IN2(StateIPG), .Q(n4) );
  MUX21X1 U26 ( .IN1(n20), .IN2(n21), .S(n12), .Q(n19) );
  AO21X1 U27 ( .IN1(NibCnt[6]), .IN2(n22), .IN3(n23), .Q(n20) );
  OA221X1 U28 ( .IN1(NibCnt[6]), .IN2(n22), .IN3(NibCnt[5]), .IN4(n25), .IN5(
        n29), .Q(n23) );
  AO221X1 U29 ( .IN1(NibCnt[4]), .IN2(n30), .IN3(NibCnt[5]), .IN4(n25), .IN5(
        n31), .Q(n29) );
  AOI222X1 U30 ( .IN1(n32), .IN2(IPGT[4]), .IN3(n33), .IN4(n34), .IN5(n35), 
        .IN6(IPGT[3]), .QN(n31) );
  OR2X1 U31 ( .IN1(IPGT[3]), .IN2(n35), .Q(n34) );
  AO22X1 U32 ( .IN1(IPGT[2]), .IN2(n36), .IN3(n37), .IN4(n38), .Q(n35) );
  OR2X1 U33 ( .IN1(n36), .IN2(IPGT[2]), .Q(n37) );
  AO22X1 U34 ( .IN1(IPGT[1]), .IN2(n39), .IN3(n40), .IN4(IPGT[0]), .Q(n36) );
  OA21X1 U35 ( .IN1(IPGT[1]), .IN2(n39), .IN3(n41), .Q(n40) );
  INVX0 U36 ( .INP(IPGT[4]), .ZN(n30) );
  INVX0 U37 ( .INP(IPGT[5]), .ZN(n25) );
  INVX0 U38 ( .INP(IPGT[6]), .ZN(n22) );
  NOR2X0 U39 ( .IN1(StartIPG), .IN2(StateIPG), .QN(n18) );
  OA21X1 U40 ( .IN1(StartBackoff), .IN2(StateBackOff), .IN3(n17), .Q(n69) );
  INVX0 U41 ( .INP(StartDefer), .ZN(n17) );
  AND3X1 U42 ( .IN1(n42), .IN2(StateIdle), .IN3(TxStartFrm), .Q(StartPreamble)
         );
  OA21X1 U43 ( .IN1(Collision), .IN2(UnderRun), .IN3(n43), .Q(StartJam) );
  NAND4X0 U44 ( .IN1(n28), .IN2(n27), .IN3(n44), .IN4(n26), .QN(n43) );
  OA21X1 U45 ( .IN1(n102), .IN2(n45), .IN3(n24), .Q(n44) );
  INVX0 U46 ( .INP(NibCntEq15), .ZN(n45) );
  NOR3X0 U47 ( .IN1(n101), .IN2(ExcessiveDefer), .IN3(CarrierSense), .QN(
        StartIPG) );
  NAND4X0 U48 ( .IN1(n46), .IN2(n47), .IN3(n48), .IN4(n49), .QN(StartDefer) );
  NOR3X0 U49 ( .IN1(DeferIndication), .IN2(TooBig), .IN3(StartTxDone), .QN(n49) );
  OAI21X1 U50 ( .IN1(RandomEqByteCnt), .IN2(TxUnderRun), .IN3(StateBackOff), 
        .QN(n48) );
  NAND4X0 U51 ( .IN1(n50), .IN2(CarrierSense), .IN3(n51), .IN4(n52), .QN(n47)
         );
  NAND4X0 U52 ( .IN1(n53), .IN2(n54), .IN3(n55), .IN4(n56), .QN(n52) );
  OA221X1 U53 ( .IN1(IPGR2[5]), .IN2(n57), .IN3(IPGR2[0]), .IN4(n41), .IN5(n58), .Q(n56) );
  OA21X1 U54 ( .IN1(IPGR2[6]), .IN2(n59), .IN3(n21), .Q(n58) );
  AOI22X1 U55 ( .IN1(IPGR2[6]), .IN2(n60), .IN3(n61), .IN4(n59), .QN(n21) );
  OR2X1 U56 ( .IN1(n60), .IN2(IPGR2[6]), .Q(n61) );
  AO22X1 U57 ( .IN1(IPGR2[5]), .IN2(n62), .IN3(n63), .IN4(n57), .Q(n60) );
  OR2X1 U58 ( .IN1(n62), .IN2(IPGR2[5]), .Q(n63) );
  AO22X1 U59 ( .IN1(IPGR2[4]), .IN2(n32), .IN3(n64), .IN4(n65), .Q(n62) );
  NAND2X0 U60 ( .IN1(NibCnt[3]), .IN2(n66), .QN(n65) );
  NOR2X0 U61 ( .IN1(n67), .IN2(n68), .QN(n64) );
  OA222X1 U62 ( .IN1(NibCnt[3]), .IN2(n66), .IN3(n78), .IN4(n79), .IN5(
        NibCnt[2]), .IN6(n80), .Q(n68) );
  OA22X1 U63 ( .IN1(NibCnt[1]), .IN2(n81), .IN3(n82), .IN4(n83), .Q(n79) );
  AO21X1 U64 ( .IN1(NibCnt[1]), .IN2(n81), .IN3(NibCnt[0]), .Q(n83) );
  INVX0 U65 ( .INP(IPGR2[0]), .ZN(n82) );
  INVX0 U66 ( .INP(IPGR2[1]), .ZN(n81) );
  INVX0 U67 ( .INP(n53), .ZN(n78) );
  INVX0 U68 ( .INP(IPGR2[3]), .ZN(n66) );
  OA22X1 U69 ( .IN1(IPGR2[1]), .IN2(n39), .IN3(IPGR2[3]), .IN4(n33), .Q(n55)
         );
  INVX0 U70 ( .INP(n67), .ZN(n54) );
  NOR2X0 U71 ( .IN1(n32), .IN2(IPGR2[4]), .QN(n67) );
  NAND2X0 U72 ( .IN1(NibCnt[2]), .IN2(n80), .QN(n53) );
  INVX0 U73 ( .INP(IPGR2[2]), .ZN(n80) );
  NOR2X0 U74 ( .IN1(n108), .IN2(n84), .QN(n51) );
  OA22X1 U75 ( .IN1(NibCnt[6]), .IN2(n85), .IN3(n86), .IN4(n87), .Q(n84) );
  AOI222X1 U76 ( .IN1(n57), .IN2(IPGR1[5]), .IN3(n32), .IN4(n88), .IN5(n89), 
        .IN6(IPGR1[4]), .QN(n87) );
  OR2X1 U77 ( .IN1(IPGR1[4]), .IN2(n89), .Q(n88) );
  AO22X1 U78 ( .IN1(IPGR1[3]), .IN2(n90), .IN3(n91), .IN4(n33), .Q(n89) );
  INVX0 U79 ( .INP(NibCnt[3]), .ZN(n33) );
  OR2X1 U80 ( .IN1(n90), .IN2(IPGR1[3]), .Q(n91) );
  AO22X1 U81 ( .IN1(IPGR1[2]), .IN2(n92), .IN3(n93), .IN4(n38), .Q(n90) );
  INVX0 U82 ( .INP(NibCnt[2]), .ZN(n38) );
  OR2X1 U83 ( .IN1(n92), .IN2(IPGR1[2]), .Q(n93) );
  AO22X1 U84 ( .IN1(IPGR1[1]), .IN2(n94), .IN3(n95), .IN4(n39), .Q(n92) );
  INVX0 U85 ( .INP(NibCnt[1]), .ZN(n39) );
  OR2X1 U86 ( .IN1(n94), .IN2(IPGR1[1]), .Q(n95) );
  OR2X1 U87 ( .IN1(IPGR1[0]), .IN2(n41), .Q(n94) );
  INVX0 U88 ( .INP(NibCnt[0]), .ZN(n41) );
  INVX0 U89 ( .INP(NibCnt[4]), .ZN(n32) );
  NOR2X0 U90 ( .IN1(IPGR1[5]), .IN2(n57), .QN(n86) );
  INVX0 U91 ( .INP(NibCnt[5]), .ZN(n57) );
  INVX0 U92 ( .INP(IPGR1[6]), .ZN(n85) );
  OA21X1 U93 ( .IN1(IPGR1[6]), .IN2(n59), .IN3(n12), .Q(n50) );
  INVX0 U94 ( .INP(NibCnt[6]), .ZN(n59) );
  NAND3X0 U95 ( .IN1(n96), .IN2(StateJam), .IN3(NibCntEq7), .QN(n46) );
  INVX0 U96 ( .INP(n97), .ZN(n96) );
  NOR4X0 U97 ( .IN1(n28), .IN2(TxUnderRun), .IN3(MaxFrame), .IN4(Collision), 
        .QN(StartData[1]) );
  AND2X1 U98 ( .IN1(n98), .IN2(n14), .Q(StartData[0]) );
  INVX0 U99 ( .INP(Collision), .ZN(n14) );
  AO22X1 U100 ( .IN1(n15), .IN2(StateData[1]), .IN3(NibCntEq15), .IN4(
        StatePreamble), .Q(n98) );
  INVX0 U101 ( .INP(TxEndFrm), .ZN(n15) );
  AND3X1 U102 ( .IN1(NibCntEq7), .IN2(StateJam), .IN3(n97), .Q(StartBackoff)
         );
  NOR4X0 U103 ( .IN1(NoBckof), .IN2(n99), .IN3(RetryMax), .IN4(RandomEq0), 
        .QN(n97) );
  INVX0 U104 ( .INP(ColWindow), .ZN(n99) );
  NOR2X0 U105 ( .IN1(n42), .IN2(n103), .QN(DeferIndication) );
  INVX0 U106 ( .INP(CarrierSense), .ZN(n42) );
endmodule


module eth_crc_test_0 ( Clk, Reset, Data, Enable, Initialize, Crc, CrcError, 
        eth_top_test_point_11887_in, test_si, test_se );
  input [3:0] Data;
  output [31:0] Crc;
  input Clk, Reset, Enable, Initialize, eth_top_test_point_11887_in, test_si,
         test_se;
  output CrcError;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N83, n35, n36, n97, n98, n99, n100, n101, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n68, n69, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59;
  assign CrcError = N83;

  SDFFASX1 \Crc_reg[0]  ( .D(N3), .SI(test_si), .SE(test_se), .CLK(Clk), 
        .SETB(n59), .Q(Crc[0]), .QN(n99) );
  SDFFASX1 \Crc_reg[4]  ( .D(N7), .SI(Crc[3]), .SE(test_se), .CLK(Clk), .SETB(
        n59), .Q(Crc[4]), .QN(n121) );
  SDFFASX1 \Crc_reg[8]  ( .D(N11), .SI(Crc[7]), .SE(test_se), .CLK(Clk), 
        .SETB(n59), .Q(Crc[8]), .QN(n117) );
  SDFFASX1 \Crc_reg[12]  ( .D(N15), .SI(Crc[11]), .SE(test_se), .CLK(Clk), 
        .SETB(n59), .Q(Crc[12]), .QN(n113) );
  SDFFASX1 \Crc_reg[16]  ( .D(N19), .SI(Crc[15]), .SE(test_se), .CLK(Clk), 
        .SETB(n59), .Q(Crc[16]), .QN(n35) );
  SDFFASX1 \Crc_reg[20]  ( .D(N23), .SI(Crc[19]), .SE(test_se), .CLK(Clk), 
        .SETB(n59), .Q(Crc[20]), .QN(n107) );
  SDFFASX1 \Crc_reg[24]  ( .D(N27), .SI(Crc[23]), .SE(test_se), .CLK(Clk), 
        .SETB(n59), .Q(Crc[24]), .QN(n103) );
  SDFFASX1 \Crc_reg[28]  ( .D(N31), .SI(Crc[27]), .SE(test_se), .CLK(Clk), 
        .SETB(n59), .Q(Crc[28]), .QN(n124) );
  SDFFASX1 \Crc_reg[22]  ( .D(N25), .SI(Crc[21]), .SE(test_se), .CLK(Clk), 
        .SETB(n59), .Q(Crc[22]), .QN(n105) );
  SDFFASX1 \Crc_reg[26]  ( .D(N29), .SI(Crc[25]), .SE(test_se), .CLK(Clk), 
        .SETB(n59), .Q(Crc[26]), .QN(n101) );
  SDFFASX1 \Crc_reg[30]  ( .D(N33), .SI(Crc[29]), .SE(test_se), .CLK(Clk), 
        .SETB(n59), .Q(Crc[30]), .QN(n68) );
  SDFFASX1 \Crc_reg[25]  ( .D(N28), .SI(Crc[24]), .SE(test_se), .CLK(Clk), 
        .SETB(n59), .Q(Crc[25]) );
  SDFFASX1 \Crc_reg[29]  ( .D(N32), .SI(Crc[28]), .SE(test_se), .CLK(Clk), 
        .SETB(n59), .Q(Crc[29]), .QN(n122) );
  SDFFASX1 \Crc_reg[1]  ( .D(N4), .SI(Crc[0]), .SE(test_se), .CLK(Clk), .SETB(
        n59), .Q(Crc[1]), .QN(n98) );
  SDFFASX1 \Crc_reg[2]  ( .D(N5), .SI(Crc[1]), .SE(test_se), .CLK(Clk), .SETB(
        n59), .Q(Crc[2]), .QN(n97) );
  SDFFASX1 \Crc_reg[6]  ( .D(N9), .SI(Crc[5]), .SE(test_se), .CLK(Clk), .SETB(
        n59), .Q(Crc[6]), .QN(n119) );
  SDFFASX1 \Crc_reg[10]  ( .D(N13), .SI(Crc[9]), .SE(test_se), .CLK(Clk), 
        .SETB(n59), .Q(Crc[10]), .QN(n115) );
  SDFFASX1 \Crc_reg[3]  ( .D(N6), .SI(Crc[2]), .SE(test_se), .CLK(Clk), .SETB(
        n59), .Q(Crc[3]), .QN(n123) );
  SDFFASX1 \Crc_reg[7]  ( .D(N10), .SI(Crc[6]), .SE(test_se), .CLK(Clk), 
        .SETB(n59), .Q(Crc[7]), .QN(n118) );
  SDFFASX1 \Crc_reg[27]  ( .D(N30), .SI(Crc[26]), .SE(test_se), .CLK(Clk), 
        .SETB(n59), .Q(Crc[27]), .QN(n100) );
  SDFFASX1 \Crc_reg[31]  ( .D(N34), .SI(Crc[30]), .SE(test_se), .CLK(Clk), 
        .SETB(n59), .Q(Crc[31]), .QN(n69) );
  SDFFASX1 \Crc_reg[5]  ( .D(N8), .SI(Crc[4]), .SE(test_se), .CLK(Clk), .SETB(
        n59), .Q(Crc[5]), .QN(n120) );
  SDFFASX1 \Crc_reg[9]  ( .D(N12), .SI(Crc[8]), .SE(test_se), .CLK(Clk), 
        .SETB(n59), .Q(Crc[9]), .QN(n116) );
  SDFFASX1 \Crc_reg[13]  ( .D(N16), .SI(Crc[12]), .SE(test_se), .CLK(Clk), 
        .SETB(n59), .Q(Crc[13]), .QN(n36) );
  SDFFASX1 \Crc_reg[11]  ( .D(N14), .SI(Crc[10]), .SE(test_se), .CLK(Clk), 
        .SETB(n59), .Q(Crc[11]), .QN(n114) );
  SDFFASX1 \Crc_reg[15]  ( .D(N18), .SI(Crc[14]), .SE(test_se), .CLK(Clk), 
        .SETB(n59), .Q(Crc[15]), .QN(n111) );
  SDFFASX1 \Crc_reg[19]  ( .D(N22), .SI(Crc[18]), .SE(test_se), .CLK(Clk), 
        .SETB(n59), .Q(Crc[19]), .QN(n108) );
  SDFFASX1 \Crc_reg[23]  ( .D(N26), .SI(Crc[22]), .SE(test_se), .CLK(Clk), 
        .SETB(n59), .Q(Crc[23]), .QN(n104) );
  SDFFASX1 \Crc_reg[17]  ( .D(N20), .SI(Crc[16]), .SE(test_se), .CLK(Clk), 
        .SETB(n59), .Q(Crc[17]), .QN(n110) );
  SDFFASX1 \Crc_reg[21]  ( .D(N24), .SI(Crc[20]), .SE(test_se), .CLK(Clk), 
        .SETB(n59), .Q(Crc[21]), .QN(n106) );
  SDFFASX1 \Crc_reg[14]  ( .D(N17), .SI(Crc[13]), .SE(test_se), .CLK(Clk), 
        .SETB(n59), .Q(Crc[14]), .QN(n112) );
  SDFFASX1 \Crc_reg[18]  ( .D(N21), .SI(Crc[17]), .SE(test_se), .CLK(Clk), 
        .SETB(n59), .Q(Crc[18]), .QN(n109) );
  INVX0 U3 ( .INP(eth_top_test_point_11887_in), .ZN(n59) );
  NAND2X0 U4 ( .IN1(n1), .IN2(n2), .QN(N9) );
  XNOR2X1 U5 ( .IN1(n97), .IN2(n3), .Q(n1) );
  NAND2X0 U6 ( .IN1(n4), .IN2(n5), .QN(N83) );
  NOR4X0 U7 ( .IN1(n6), .IN2(n7), .IN3(n8), .IN4(n9), .QN(n5) );
  OR4X1 U8 ( .IN1(n103), .IN2(n109), .IN3(n111), .IN4(n112), .Q(n9) );
  OR4X1 U9 ( .IN1(n113), .IN2(n114), .IN3(n115), .IN4(n117), .Q(n8) );
  OR4X1 U10 ( .IN1(n119), .IN2(n120), .IN3(n121), .IN4(n123), .Q(n7) );
  OR4X1 U11 ( .IN1(n68), .IN2(n69), .IN3(n98), .IN4(n99), .Q(n6) );
  NOR4X0 U12 ( .IN1(n10), .IN2(n11), .IN3(n12), .IN4(n13), .QN(n4) );
  NAND4X0 U13 ( .IN1(n36), .IN2(n35), .IN3(n124), .IN4(n118), .QN(n13) );
  NAND4X0 U14 ( .IN1(n116), .IN2(n110), .IN3(n108), .IN4(n107), .QN(n12) );
  NAND4X0 U15 ( .IN1(n106), .IN2(n105), .IN3(n104), .IN4(n100), .QN(n11) );
  NAND4X0 U16 ( .IN1(n97), .IN2(n122), .IN3(Crc[26]), .IN4(Crc[25]), .QN(n10)
         );
  NAND2X0 U17 ( .IN1(n14), .IN2(n2), .QN(N8) );
  XNOR2X1 U18 ( .IN1(n98), .IN2(n15), .Q(n14) );
  NAND2X0 U19 ( .IN1(n16), .IN2(n2), .QN(N7) );
  XNOR2X1 U20 ( .IN1(n99), .IN2(n17), .Q(n16) );
  NAND2X0 U21 ( .IN1(n18), .IN2(n2), .QN(N6) );
  NAND2X0 U22 ( .IN1(n19), .IN2(n2), .QN(N5) );
  OR2X1 U23 ( .IN1(Initialize), .IN2(n20), .Q(N4) );
  NAND2X0 U24 ( .IN1(n100), .IN2(n2), .QN(N34) );
  NAND2X0 U25 ( .IN1(n101), .IN2(n2), .QN(N33) );
  NAND2X0 U26 ( .IN1(n21), .IN2(n2), .QN(N32) );
  XNOR2X1 U27 ( .IN1(Crc[25]), .IN2(n22), .Q(n21) );
  NAND2X0 U28 ( .IN1(n23), .IN2(n2), .QN(N31) );
  XOR2X1 U29 ( .IN1(n103), .IN2(n24), .Q(n23) );
  NAND2X0 U30 ( .IN1(n25), .IN2(n2), .QN(N30) );
  XOR2X1 U31 ( .IN1(n104), .IN2(n26), .Q(n25) );
  OR2X1 U32 ( .IN1(Initialize), .IN2(n27), .Q(N3) );
  NAND2X0 U33 ( .IN1(n28), .IN2(n2), .QN(N29) );
  XNOR2X1 U34 ( .IN1(n105), .IN2(n29), .Q(n28) );
  NAND2X0 U35 ( .IN1(Enable), .IN2(n30), .QN(n29) );
  XOR2X1 U36 ( .IN1(n31), .IN2(n32), .Q(n30) );
  NAND2X0 U37 ( .IN1(n33), .IN2(n2), .QN(N28) );
  XOR2X1 U38 ( .IN1(n106), .IN2(n34), .Q(n33) );
  NAND2X0 U39 ( .IN1(n37), .IN2(n2), .QN(N27) );
  XNOR2X1 U40 ( .IN1(n107), .IN2(n3), .Q(n37) );
  NAND2X0 U41 ( .IN1(n38), .IN2(n2), .QN(N26) );
  XOR2X1 U42 ( .IN1(n108), .IN2(n20), .Q(n38) );
  NAND2X0 U43 ( .IN1(n39), .IN2(n2), .QN(N25) );
  XOR2X1 U44 ( .IN1(n109), .IN2(n27), .Q(n39) );
  NAND2X0 U45 ( .IN1(n110), .IN2(n2), .QN(N24) );
  NAND2X0 U46 ( .IN1(n35), .IN2(n2), .QN(N23) );
  NAND2X0 U47 ( .IN1(n40), .IN2(n2), .QN(N22) );
  XOR2X1 U48 ( .IN1(n111), .IN2(n22), .Q(n40) );
  NAND2X0 U49 ( .IN1(n41), .IN2(n2), .QN(N21) );
  XOR2X1 U50 ( .IN1(n112), .IN2(n24), .Q(n41) );
  NAND2X0 U51 ( .IN1(n42), .IN2(n2), .QN(N20) );
  XOR2X1 U52 ( .IN1(n36), .IN2(n26), .Q(n42) );
  NAND2X0 U53 ( .IN1(n43), .IN2(n2), .QN(N19) );
  XOR2X1 U54 ( .IN1(n113), .IN2(n27), .Q(n43) );
  NAND2X0 U55 ( .IN1(n44), .IN2(n2), .QN(N18) );
  XOR2X1 U56 ( .IN1(n114), .IN2(n22), .Q(n44) );
  NAND2X0 U57 ( .IN1(n45), .IN2(n2), .QN(N17) );
  XOR2X1 U58 ( .IN1(n115), .IN2(n34), .Q(n45) );
  NAND2X0 U59 ( .IN1(n46), .IN2(n2), .QN(N16) );
  XNOR2X1 U60 ( .IN1(n116), .IN2(n18), .Q(n46) );
  AOI22X1 U61 ( .IN1(n34), .IN2(n47), .IN3(n26), .IN4(n48), .QN(n18) );
  NOR2X0 U62 ( .IN1(n49), .IN2(n47), .QN(n26) );
  NAND2X0 U63 ( .IN1(n50), .IN2(n2), .QN(N15) );
  XNOR2X1 U64 ( .IN1(n117), .IN2(n19), .Q(n50) );
  AOI22X1 U65 ( .IN1(n24), .IN2(n51), .IN3(n20), .IN4(n52), .QN(n19) );
  NOR2X0 U66 ( .IN1(n49), .IN2(n52), .QN(n24) );
  NAND2X0 U67 ( .IN1(n53), .IN2(n2), .QN(N14) );
  XNOR2X1 U68 ( .IN1(n118), .IN2(n15), .Q(n53) );
  NAND2X0 U69 ( .IN1(n54), .IN2(n2), .QN(N13) );
  XNOR2X1 U70 ( .IN1(n119), .IN2(n17), .Q(n54) );
  NAND2X0 U71 ( .IN1(n55), .IN2(n2), .QN(N12) );
  XNOR2X1 U72 ( .IN1(n120), .IN2(n3), .Q(n55) );
  NAND2X0 U73 ( .IN1(Enable), .IN2(n56), .QN(n3) );
  XOR2X1 U74 ( .IN1(n47), .IN2(n52), .Q(n56) );
  NAND2X0 U75 ( .IN1(n57), .IN2(n2), .QN(N11) );
  XNOR2X1 U76 ( .IN1(n121), .IN2(n15), .Q(n57) );
  AOI22X1 U77 ( .IN1(n22), .IN2(n51), .IN3(n20), .IN4(n31), .QN(n15) );
  NOR2X0 U78 ( .IN1(n49), .IN2(n51), .QN(n20) );
  XNOR2X1 U79 ( .IN1(n32), .IN2(n47), .Q(n51) );
  XOR2X1 U80 ( .IN1(n122), .IN2(Data[1]), .Q(n47) );
  NOR2X0 U81 ( .IN1(n31), .IN2(n49), .QN(n22) );
  NAND2X0 U82 ( .IN1(n58), .IN2(n2), .QN(N10) );
  INVX0 U83 ( .INP(Initialize), .ZN(n2) );
  XNOR2X1 U84 ( .IN1(n123), .IN2(n17), .Q(n58) );
  AOI22X1 U85 ( .IN1(n34), .IN2(n32), .IN3(n27), .IN4(n48), .QN(n17) );
  NOR2X0 U86 ( .IN1(n32), .IN2(n49), .QN(n27) );
  XOR2X1 U87 ( .IN1(n124), .IN2(Data[0]), .Q(n32) );
  NOR2X0 U88 ( .IN1(n49), .IN2(n48), .QN(n34) );
  XNOR2X1 U89 ( .IN1(n31), .IN2(n52), .Q(n48) );
  XOR2X1 U90 ( .IN1(n68), .IN2(Data[2]), .Q(n52) );
  XOR2X1 U91 ( .IN1(n69), .IN2(Data[3]), .Q(n31) );
  INVX0 U92 ( .INP(Enable), .ZN(n49) );
endmodule


module eth_random_test_1 ( MTxClk, Reset, StateJam, StateJam_q, RetryCnt, 
        NibCnt, ByteCnt, RandomEq0, RandomEqByteCnt, 
        eth_top_test_point_11887_in, test_si, test_so, test_se );
  input [3:0] RetryCnt;
  input [15:0] NibCnt;
  input [9:0] ByteCnt;
  input MTxClk, Reset, StateJam, StateJam_q, eth_top_test_point_11887_in,
         test_si, test_se;
  output RandomEq0, RandomEqByteCnt, test_so;
  wire   N21, n55, n59, n60, n61, n64, n66, n68, n70, n72, n74, n76, n78, n80,
         n82, n94, n1, n2, n3, n4, n5, n6, n7, n8, n9, n46, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n47, n48, n49, n50;
  wire   [9:0] x;
  assign test_so = x[9];
  assign N21 = RetryCnt[3];

  SDFFARX1 \x_reg[0]  ( .D(n94), .SI(n4), .SE(test_se), .CLK(MTxClk), .RSTB(
        n50), .Q(x[0]) );
  SDFFARX1 \x_reg[1]  ( .D(x[0]), .SI(x[0]), .SE(test_se), .CLK(MTxClk), 
        .RSTB(n50), .Q(x[1]) );
  SDFFARX1 \x_reg[2]  ( .D(x[1]), .SI(x[1]), .SE(test_se), .CLK(MTxClk), 
        .RSTB(n50), .Q(x[2]) );
  SDFFARX1 \x_reg[3]  ( .D(x[2]), .SI(x[2]), .SE(test_se), .CLK(MTxClk), 
        .RSTB(n50), .Q(x[3]), .QN(n10) );
  SDFFARX1 \x_reg[4]  ( .D(x[3]), .SI(x[3]), .SE(test_se), .CLK(MTxClk), 
        .RSTB(n50), .Q(x[4]) );
  SDFFARX1 \x_reg[5]  ( .D(x[4]), .SI(x[4]), .SE(test_se), .CLK(MTxClk), 
        .RSTB(n50), .Q(x[5]) );
  SDFFARX1 \x_reg[6]  ( .D(x[5]), .SI(x[5]), .SE(test_se), .CLK(MTxClk), 
        .RSTB(n50), .Q(x[6]) );
  SDFFARX1 \x_reg[7]  ( .D(x[6]), .SI(x[6]), .SE(test_se), .CLK(MTxClk), 
        .RSTB(n50), .Q(x[7]) );
  SDFFARX1 \x_reg[8]  ( .D(x[7]), .SI(x[7]), .SE(test_se), .CLK(MTxClk), 
        .RSTB(n50), .Q(x[8]) );
  SDFFARX1 \x_reg[9]  ( .D(x[8]), .SI(x[8]), .SE(test_se), .CLK(MTxClk), 
        .RSTB(n50), .Q(x[9]) );
  SDFFARX1 \RandomLatched_reg[9]  ( .D(n82), .SI(n2), .SE(test_se), .CLK(
        MTxClk), .RSTB(n50), .Q(n4), .QN(n61) );
  SDFFARX1 \RandomLatched_reg[8]  ( .D(n80), .SI(n5), .SE(test_se), .CLK(
        MTxClk), .RSTB(n50), .Q(n2), .QN(n60) );
  SDFFARX1 \RandomLatched_reg[7]  ( .D(n78), .SI(n7), .SE(test_se), .CLK(
        MTxClk), .RSTB(n50), .Q(n5), .QN(n59) );
  SDFFARX1 \RandomLatched_reg[6]  ( .D(n76), .SI(n6), .SE(test_se), .CLK(
        MTxClk), .RSTB(n50), .Q(n7), .QN(n45) );
  SDFFARX1 \RandomLatched_reg[5]  ( .D(n74), .SI(n9), .SE(test_se), .CLK(
        MTxClk), .RSTB(n50), .Q(n6), .QN(n47) );
  SDFFARX1 \RandomLatched_reg[4]  ( .D(n72), .SI(n46), .SE(test_se), .CLK(
        MTxClk), .RSTB(n50), .Q(n9), .QN(n49) );
  SDFFARX1 \RandomLatched_reg[3]  ( .D(n70), .SI(n8), .SE(test_se), .CLK(
        MTxClk), .RSTB(n50), .Q(n46), .QN(n55) );
  SDFFARX1 \RandomLatched_reg[2]  ( .D(n68), .SI(n3), .SE(test_se), .CLK(
        MTxClk), .RSTB(n50), .Q(n8), .QN(n48) );
  SDFFARX1 \RandomLatched_reg[1]  ( .D(n66), .SI(n1), .SE(test_se), .CLK(
        MTxClk), .RSTB(n50), .Q(n3) );
  SDFFARX1 \RandomLatched_reg[0]  ( .D(n64), .SI(test_si), .SE(test_se), .CLK(
        MTxClk), .RSTB(n50), .Q(n1) );
  INVX0 U3 ( .INP(eth_top_test_point_11887_in), .ZN(n50) );
  XNOR2X1 U4 ( .IN1(x[2]), .IN2(x[9]), .Q(n94) );
  AO22X1 U5 ( .IN1(n11), .IN2(n4), .IN3(n12), .IN4(n13), .Q(n82) );
  AND2X1 U6 ( .IN1(n14), .IN2(x[9]), .Q(n12) );
  AO22X1 U7 ( .IN1(n11), .IN2(n2), .IN3(n15), .IN4(x[8]), .Q(n80) );
  OA21X1 U8 ( .IN1(RetryCnt[0]), .IN2(n14), .IN3(n13), .Q(n15) );
  AO22X1 U9 ( .IN1(n11), .IN2(n5), .IN3(x[7]), .IN4(n13), .Q(n78) );
  AO22X1 U10 ( .IN1(n11), .IN2(n7), .IN3(x[6]), .IN4(n16), .Q(n76) );
  NAND2X0 U11 ( .IN1(n17), .IN2(n18), .QN(n16) );
  NAND3X0 U12 ( .IN1(RetryCnt[0]), .IN2(n19), .IN3(RetryCnt[1]), .QN(n18) );
  AO22X1 U13 ( .IN1(n11), .IN2(n6), .IN3(x[5]), .IN4(n20), .Q(n74) );
  AO22X1 U14 ( .IN1(n11), .IN2(n9), .IN3(x[4]), .IN4(n21), .Q(n72) );
  AO21X1 U15 ( .IN1(RetryCnt[0]), .IN2(n19), .IN3(n20), .Q(n21) );
  AO21X1 U16 ( .IN1(RetryCnt[1]), .IN2(n19), .IN3(n13), .Q(n20) );
  OAI22X1 U17 ( .IN1(n22), .IN2(n55), .IN3(n10), .IN4(n23), .QN(n70) );
  AO22X1 U18 ( .IN1(n11), .IN2(n8), .IN3(x[2]), .IN4(n24), .Q(n68) );
  NAND2X0 U19 ( .IN1(n23), .IN2(n25), .QN(n24) );
  NAND3X0 U20 ( .IN1(RetryCnt[0]), .IN2(n22), .IN3(RetryCnt[1]), .QN(n25) );
  NOR2X0 U21 ( .IN1(n13), .IN2(n19), .QN(n23) );
  AND2X1 U22 ( .IN1(RetryCnt[2]), .IN2(n22), .Q(n19) );
  AO22X1 U23 ( .IN1(n11), .IN2(n3), .IN3(x[1]), .IN4(n26), .Q(n66) );
  AO21X1 U24 ( .IN1(n22), .IN2(n14), .IN3(n13), .Q(n26) );
  INVX0 U25 ( .INP(n17), .ZN(n13) );
  NAND2X0 U26 ( .IN1(N21), .IN2(n22), .QN(n17) );
  OR2X1 U27 ( .IN1(RetryCnt[2]), .IN2(RetryCnt[1]), .Q(n14) );
  MUX21X1 U28 ( .IN1(n1), .IN2(x[0]), .S(n22), .Q(n64) );
  INVX0 U29 ( .INP(n11), .ZN(n22) );
  NAND2X0 U30 ( .IN1(StateJam_q), .IN2(StateJam), .QN(n11) );
  NOR4X0 U31 ( .IN1(n27), .IN2(n28), .IN3(n29), .IN4(n30), .QN(RandomEqByteCnt) );
  NAND4X0 U32 ( .IN1(NibCnt[6]), .IN2(NibCnt[5]), .IN3(NibCnt[4]), .IN4(
        NibCnt[3]), .QN(n30) );
  NAND4X0 U33 ( .IN1(NibCnt[2]), .IN2(NibCnt[1]), .IN3(NibCnt[0]), .IN4(n31), 
        .QN(n29) );
  XOR2X1 U34 ( .IN1(n45), .IN2(ByteCnt[6]), .Q(n31) );
  NAND4X0 U35 ( .IN1(n32), .IN2(n33), .IN3(n34), .IN4(n35), .QN(n28) );
  XOR2X1 U36 ( .IN1(n61), .IN2(ByteCnt[9]), .Q(n35) );
  XOR2X1 U37 ( .IN1(n48), .IN2(ByteCnt[2]), .Q(n34) );
  XOR2X1 U38 ( .IN1(n49), .IN2(ByteCnt[4]), .Q(n33) );
  XOR2X1 U39 ( .IN1(n47), .IN2(ByteCnt[5]), .Q(n32) );
  NAND4X0 U40 ( .IN1(n36), .IN2(n37), .IN3(n38), .IN4(n39), .QN(n27) );
  XOR2X1 U41 ( .IN1(n55), .IN2(ByteCnt[3]), .Q(n39) );
  NOR2X0 U42 ( .IN1(n40), .IN2(n41), .QN(n38) );
  XOR2X1 U43 ( .IN1(n1), .IN2(ByteCnt[0]), .Q(n41) );
  XOR2X1 U44 ( .IN1(n3), .IN2(ByteCnt[1]), .Q(n40) );
  XOR2X1 U45 ( .IN1(n59), .IN2(ByteCnt[7]), .Q(n37) );
  XOR2X1 U46 ( .IN1(n60), .IN2(ByteCnt[8]), .Q(n36) );
  NOR4X0 U47 ( .IN1(n42), .IN2(n43), .IN3(n6), .IN4(n7), .QN(RandomEq0) );
  NAND3X0 U48 ( .IN1(n48), .IN2(n61), .IN3(n49), .QN(n43) );
  NAND4X0 U49 ( .IN1(n60), .IN2(n59), .IN3(n44), .IN4(n55), .QN(n42) );
  NOR2X0 U50 ( .IN1(n3), .IN2(n1), .QN(n44) );
endmodule


module eth_txethmac_test_1 ( MTxClk, Reset, TxStartFrm, TxEndFrm, TxUnderRun, 
        TxData, CarrierSense, Collision, Pad, CrcEn, FullD, HugEn, DlyCrcEn, 
        MinFL, MaxFL, IPGT, IPGR1, IPGR2, CollValid, MaxRet, NoBckof, ExDfrEn, 
        MTxD, MTxEn, MTxErr, TxDone, TxRetry, TxAbort, TxUsedData, 
        WillTransmit, ResetCollision, RetryCnt, StartTxDone, StartTxAbort, 
        MaxCollisionOccured, LateCollision, DeferIndication, StatePreamble, 
        StateData, eth_top_test_point_11887_in, test_si2, test_si1, test_se );
  input [7:0] TxData;
  input [15:0] MinFL;
  input [15:0] MaxFL;
  input [6:0] IPGT;
  input [6:0] IPGR1;
  input [6:0] IPGR2;
  input [5:0] CollValid;
  input [3:0] MaxRet;
  output [3:0] MTxD;
  output [3:0] RetryCnt;
  output [1:0] StateData;
  input MTxClk, Reset, TxStartFrm, TxEndFrm, TxUnderRun, CarrierSense,
         Collision, Pad, CrcEn, FullD, HugEn, DlyCrcEn, NoBckof, ExDfrEn,
         eth_top_test_point_11887_in, test_si2, test_si1, test_se;
  output MTxEn, MTxErr, TxDone, TxRetry, TxAbort, TxUsedData, WillTransmit,
         ResetCollision, StartTxDone, StartTxAbort, MaxCollisionOccured,
         LateCollision, DeferIndication, StatePreamble;
  wire   StatePAD, StateFCS, StateDefer, ExcessiveDefer, NibCntEq7,
         NibbleMinFl, UnderRun, MaxFrame, TooBig, StartJam, ColWindow,
         NibCntEq15, StateSFD, StateIdle, StateIPG, N29, StateJam, RandomEq0,
         StateBackOff, RandomEqByteCnt, N86, StartPreamble, N88,
         PacketFinished_d, PacketFinished_q, PacketFinished, StartDefer,
         StartIPG, StartFCS, StartBackoff, StateJam_q, Initialize_Crc, n33,
         n34, n35, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n94, n95, n111, n112, n113, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;
  wire   [15:0] NibCnt;
  wire   [15:0] ByteCnt;
  wire   [1:0] StartData;
  wire   [31:0] Crc;
  wire   [3:0] MTxD_d;
  wire   [2:0] DlyCrcCnt;
  wire   [3:0] Data_Crc;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33;

  SDFFARX1 PacketFinished_q_reg ( .D(PacketFinished), .SI(MTxEn), .SE(test_se), 
        .CLK(n2), .RSTB(n81), .Q(PacketFinished_q) );
  SDFFARX1 \RetryCnt_reg[1]  ( .D(n106), .SI(RetryCnt[0]), .SE(test_se), .CLK(
        n1), .RSTB(n81), .Q(RetryCnt[1]), .QN(n34) );
  SDFFARX1 \RetryCnt_reg[2]  ( .D(n105), .SI(RetryCnt[1]), .SE(test_se), .CLK(
        n2), .RSTB(n81), .Q(RetryCnt[2]), .QN(n95) );
  SDFFARX1 \RetryCnt_reg[3]  ( .D(n104), .SI(RetryCnt[2]), .SE(test_se), .CLK(
        n2), .RSTB(n81), .Q(RetryCnt[3]), .QN(n33) );
  SDFFARX1 TxUsedData_reg ( .D(N29), .SI(TxRetry), .SE(test_se), .CLK(n2), 
        .RSTB(n81), .Q(TxUsedData) );
  SDFFARX1 StopExcessiveDeferOccured_reg ( .D(n109), .SI(n113), .SE(test_se), 
        .CLK(n2), .RSTB(n81), .Q(n112), .QN(n77) );
  SDFFARX1 MTxErr_reg ( .D(n78), .SI(test_si2), .SE(test_se), .CLK(n1), .RSTB(
        n81), .Q(MTxErr) );
  SDFFARX1 MTxEn_reg ( .D(N86), .SI(MTxD[3]), .SE(test_se), .CLK(n2), .RSTB(
        n81), .Q(MTxEn) );
  SDFFARX1 WillTransmit_reg ( .D(N88), .SI(TxUsedData), .SE(test_se), .CLK(n2), 
        .RSTB(n81), .Q(WillTransmit) );
  SDFFASX1 ColWindow_reg ( .D(n108), .SI(test_si1), .SE(test_se), .CLK(n1), 
        .SETB(n81), .Q(ColWindow) );
  SDFFARX1 StatusLatch_reg ( .D(n103), .SI(RetryCnt[3]), .SE(test_se), .CLK(n2), .RSTB(n81), .Q(n113), .QN(n94) );
  SDFFARX1 TxDone_reg ( .D(n100), .SI(TxAbort), .SE(test_se), .CLK(n2), .RSTB(
        n81), .Q(TxDone) );
  SDFFARX1 \MTxD_reg[3]  ( .D(MTxD_d[3]), .SI(MTxD[2]), .SE(test_se), .CLK(n2), 
        .RSTB(n81), .Q(MTxD[3]) );
  SDFFARX1 \MTxD_reg[2]  ( .D(MTxD_d[2]), .SI(MTxD[1]), .SE(test_se), .CLK(n2), 
        .RSTB(n81), .Q(MTxD[2]) );
  SDFFARX1 \MTxD_reg[1]  ( .D(MTxD_d[1]), .SI(MTxD[0]), .SE(test_se), .CLK(n2), 
        .RSTB(n81), .Q(MTxD[1]) );
  SDFFARX1 \MTxD_reg[0]  ( .D(MTxD_d[0]), .SI(ColWindow), .SE(test_se), .CLK(
        n2), .RSTB(n81), .Q(MTxD[0]) );
  SDFFARX1 TxRetry_reg ( .D(n101), .SI(TxDone), .SE(test_se), .CLK(n2), .RSTB(
        n81), .Q(TxRetry) );
  SDFFARX1 \RetryCnt_reg[0]  ( .D(n107), .SI(PacketFinished), .SE(test_se), 
        .CLK(n1), .RSTB(n81), .Q(RetryCnt[0]), .QN(n35) );
  SDFFARX1 PacketFinished_reg ( .D(PacketFinished_d), .SI(PacketFinished_q), 
        .SE(test_se), .CLK(n2), .RSTB(n81), .Q(PacketFinished) );
  SDFFARX1 TxAbort_reg ( .D(n102), .SI(n112), .SE(test_se), .CLK(n2), .RSTB(
        n81), .Q(TxAbort) );
  eth_txcounters_test_1 txcounters1 ( .StatePreamble(StatePreamble), 
        .StateIPG(StateIPG), .StateData(StateData), .StatePAD(StatePAD), 
        .StateFCS(StateFCS), .StateJam(StateJam), .StateBackOff(StateBackOff), 
        .StateDefer(StateDefer), .StateIdle(StateIdle), .StartDefer(StartDefer), .StartIPG(StartIPG), .StartFCS(StartFCS), .StartJam(StartJam), 
        .StartBackoff(StartBackoff), .TxStartFrm(TxStartFrm), .MTxClk(n1), 
        .Reset(Reset), .MinFL(MinFL), .MaxFL(MaxFL), .HugEn(HugEn), .ExDfrEn(
        ExDfrEn), .PacketFinished_q(PacketFinished_q), .DlyCrcEn(DlyCrcEn), 
        .StateSFD(StateSFD), .ByteCnt({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, ByteCnt[9:0]}), .NibCnt(NibCnt), 
        .ExcessiveDefer(ExcessiveDefer), .NibCntEq7(NibCntEq7), .NibCntEq15(
        NibCntEq15), .MaxFrame(MaxFrame), .NibbleMinFl(NibbleMinFl), 
        .DlyCrcCnt(DlyCrcCnt), .eth_top_test_point_11887_in(
        eth_top_test_point_11887_in), .test_si(n111), .test_se(test_se) );
  eth_txstatem_test_1 txstatem1 ( .MTxClk(n2), .Reset(Reset), .ExcessiveDefer(
        ExcessiveDefer), .CarrierSense(CarrierSense), .NibCnt(NibCnt[6:0]), 
        .IPGT(IPGT), .IPGR1(IPGR1), .IPGR2(IPGR2), .FullD(FullD), .TxStartFrm(
        TxStartFrm), .TxEndFrm(TxEndFrm), .TxUnderRun(TxUnderRun), .Collision(
        Collision), .UnderRun(UnderRun), .StartTxDone(StartTxDone), .TooBig(
        TooBig), .NibCntEq7(NibCntEq7), .NibCntEq15(NibCntEq15), .MaxFrame(
        MaxFrame), .Pad(Pad), .CrcEn(CrcEn), .NibbleMinFl(NibbleMinFl), 
        .RandomEq0(RandomEq0), .ColWindow(ColWindow), .RetryMax(n80), 
        .NoBckof(NoBckof), .RandomEqByteCnt(RandomEqByteCnt), .StateIdle(
        StateIdle), .StateIPG(StateIPG), .StatePreamble(StatePreamble), 
        .StateData(StateData), .StatePAD(StatePAD), .StateFCS(StateFCS), 
        .StateJam(StateJam), .StateJam_q(StateJam_q), .StateBackOff(
        StateBackOff), .StateDefer(StateDefer), .StartFCS(StartFCS), 
        .StartJam(StartJam), .StartBackoff(StartBackoff), .StartDefer(
        StartDefer), .DeferIndication(DeferIndication), .StartPreamble(
        StartPreamble), .StartData(StartData), .StartIPG(StartIPG), 
        .eth_top_test_point_11887_in(eth_top_test_point_11887_in), .test_si(
        Crc[31]), .test_se(test_se) );
  eth_crc_test_0 txcrc ( .Clk(n1), .Reset(Reset), .Data(Data_Crc), .Enable(n79), .Initialize(Initialize_Crc), .Crc({Crc[31:28], SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, SYNOPSYS_UNCONNECTED__16, 
        SYNOPSYS_UNCONNECTED__17, SYNOPSYS_UNCONNECTED__18, 
        SYNOPSYS_UNCONNECTED__19, SYNOPSYS_UNCONNECTED__20, 
        SYNOPSYS_UNCONNECTED__21, SYNOPSYS_UNCONNECTED__22, 
        SYNOPSYS_UNCONNECTED__23, SYNOPSYS_UNCONNECTED__24, 
        SYNOPSYS_UNCONNECTED__25, SYNOPSYS_UNCONNECTED__26, 
        SYNOPSYS_UNCONNECTED__27, SYNOPSYS_UNCONNECTED__28, 
        SYNOPSYS_UNCONNECTED__29, SYNOPSYS_UNCONNECTED__30, 
        SYNOPSYS_UNCONNECTED__31, SYNOPSYS_UNCONNECTED__32, 
        SYNOPSYS_UNCONNECTED__33}), .eth_top_test_point_11887_in(
        eth_top_test_point_11887_in), .test_si(NibCnt[15]), .test_se(test_se)
         );
  eth_random_test_1 random1 ( .MTxClk(n2), .Reset(Reset), .StateJam(StateJam), 
        .StateJam_q(StateJam_q), .RetryCnt(RetryCnt), .NibCnt(NibCnt), 
        .ByteCnt(ByteCnt[9:0]), .RandomEq0(RandomEq0), .RandomEqByteCnt(
        RandomEqByteCnt), .eth_top_test_point_11887_in(
        eth_top_test_point_11887_in), .test_si(WillTransmit), .test_so(n111), 
        .test_se(test_se) );
  NBUFFX4 U3 ( .INP(MTxClk), .Z(n2) );
  DELLN1X2 U4 ( .INP(MTxClk), .Z(n1) );
  INVX0 U5 ( .INP(eth_top_test_point_11887_in), .ZN(n81) );
  AOI21X1 U6 ( .IN1(n3), .IN2(n77), .IN3(n4), .QN(n109) );
  NOR2X0 U7 ( .IN1(n5), .IN2(n6), .QN(n108) );
  NOR3X0 U8 ( .IN1(ColWindow), .IN2(StateIdle), .IN3(StateIPG), .QN(n6) );
  NOR4X0 U9 ( .IN1(n7), .IN2(n8), .IN3(n9), .IN4(n10), .QN(n5) );
  XOR2X1 U10 ( .IN1(CollValid[2]), .IN2(ByteCnt[2]), .Q(n10) );
  XOR2X1 U11 ( .IN1(CollValid[0]), .IN2(ByteCnt[0]), .Q(n9) );
  NAND3X0 U12 ( .IN1(n11), .IN2(n12), .IN3(n13), .QN(n8) );
  OR2X1 U13 ( .IN1(NibCnt[0]), .IN2(StateData[1]), .Q(n13) );
  NAND4X0 U14 ( .IN1(n14), .IN2(n15), .IN3(n16), .IN4(n17), .QN(n7) );
  XNOR2X1 U15 ( .IN1(CollValid[1]), .IN2(ByteCnt[1]), .Q(n17) );
  XNOR2X1 U16 ( .IN1(CollValid[3]), .IN2(ByteCnt[3]), .Q(n16) );
  XNOR2X1 U17 ( .IN1(CollValid[4]), .IN2(ByteCnt[4]), .Q(n15) );
  XNOR2X1 U18 ( .IN1(CollValid[5]), .IN2(ByteCnt[5]), .Q(n14) );
  MUX21X1 U19 ( .IN1(n18), .IN2(n19), .S(RetryCnt[0]), .Q(n107) );
  NOR2X0 U20 ( .IN1(n18), .IN2(n20), .QN(n19) );
  MUX21X1 U21 ( .IN1(n21), .IN2(n22), .S(RetryCnt[1]), .Q(n106) );
  AND2X1 U22 ( .IN1(RetryCnt[0]), .IN2(n18), .Q(n21) );
  MUX21X1 U23 ( .IN1(n23), .IN2(n24), .S(n95), .Q(n105) );
  INVX0 U24 ( .INP(n25), .ZN(n24) );
  MUX21X1 U25 ( .IN1(n26), .IN2(n27), .S(n33), .Q(n104) );
  NOR2X0 U26 ( .IN1(n95), .IN2(n25), .QN(n27) );
  NAND3X0 U27 ( .IN1(RetryCnt[1]), .IN2(RetryCnt[0]), .IN3(n18), .QN(n25) );
  AO21X1 U28 ( .IN1(n18), .IN2(n95), .IN3(n23), .Q(n26) );
  AO21X1 U29 ( .IN1(n18), .IN2(n34), .IN3(n22), .Q(n23) );
  MUX21X1 U30 ( .IN1(n28), .IN2(n35), .S(n18), .Q(n22) );
  INVX0 U31 ( .INP(n20), .ZN(n28) );
  NOR2X0 U32 ( .IN1(n20), .IN2(n29), .QN(n18) );
  AOI22X1 U33 ( .IN1(StateBackOff), .IN2(RandomEqByteCnt), .IN3(n30), .IN4(
        StateJam), .QN(n29) );
  OA21X1 U34 ( .IN1(RandomEq0), .IN2(NoBckof), .IN3(NibCntEq7), .Q(n30) );
  NAND4X0 U35 ( .IN1(n31), .IN2(n3), .IN3(n32), .IN4(n36), .QN(n20) );
  INVX0 U36 ( .INP(StartTxDone), .ZN(n36) );
  NOR2X0 U37 ( .IN1(TxUnderRun), .IN2(n78), .QN(n32) );
  INVX0 U38 ( .INP(n37), .ZN(n78) );
  NAND3X0 U39 ( .IN1(NibCntEq7), .IN2(n38), .IN3(StateJam), .QN(n31) );
  NOR2X0 U40 ( .IN1(n39), .IN2(n4), .QN(n103) );
  INVX0 U41 ( .INP(TxStartFrm), .ZN(n4) );
  AND3X1 U42 ( .IN1(n3), .IN2(n40), .IN3(n94), .Q(n39) );
  AO22X1 U43 ( .IN1(n41), .IN2(TxAbort), .IN3(n42), .IN4(StartTxAbort), .Q(
        n102) );
  NAND2X0 U44 ( .IN1(n43), .IN2(n3), .QN(n42) );
  INVX0 U45 ( .INP(n41), .ZN(n43) );
  OA21X1 U46 ( .IN1(n44), .IN2(TxRetry), .IN3(n41), .Q(n101) );
  NOR3X0 U47 ( .IN1(n38), .IN2(UnderRun), .IN3(n45), .QN(n44) );
  OA21X1 U48 ( .IN1(StartTxDone), .IN2(TxDone), .IN3(n41), .Q(n100) );
  NAND2X0 U49 ( .IN1(n94), .IN2(TxStartFrm), .QN(n41) );
  NOR2X0 U50 ( .IN1(n46), .IN2(n47), .QN(StateSFD) );
  OR2X1 U51 ( .IN1(StartTxAbort), .IN2(StartTxDone), .Q(PacketFinished_d) );
  NOR2X0 U52 ( .IN1(Collision), .IN2(n48), .QN(StartTxDone) );
  OA22X1 U53 ( .IN1(n49), .IN2(n50), .IN3(n79), .IN4(n51), .Q(n48) );
  INVX0 U54 ( .INP(NibCntEq7), .ZN(n51) );
  NAND2X0 U55 ( .IN1(TxEndFrm), .IN2(StateData[1]), .QN(n50) );
  AO21X1 U56 ( .IN1(Pad), .IN2(n52), .IN3(CrcEn), .Q(n49) );
  INVX0 U57 ( .INP(NibbleMinFl), .ZN(n52) );
  NAND3X0 U58 ( .IN1(n3), .IN2(n37), .IN3(n53), .QN(StartTxAbort) );
  NAND2X0 U59 ( .IN1(StartJam), .IN2(n38), .QN(n53) );
  NAND2X0 U60 ( .IN1(ColWindow), .IN2(n54), .QN(n38) );
  NOR2X0 U61 ( .IN1(UnderRun), .IN2(TooBig), .QN(n37) );
  AND3X1 U62 ( .IN1(n55), .IN2(n12), .IN3(MaxFrame), .Q(TooBig) );
  OAI21X1 U63 ( .IN1(n56), .IN2(TxUnderRun), .IN3(n79), .QN(n55) );
  INVX0 U64 ( .INP(StateFCS), .ZN(n79) );
  NAND4X0 U65 ( .IN1(n77), .IN2(TxStartFrm), .IN3(StateDefer), .IN4(
        ExcessiveDefer), .QN(n3) );
  OR2X1 U66 ( .IN1(StartPreamble), .IN2(N86), .Q(N88) );
  NAND2X0 U67 ( .IN1(ResetCollision), .IN2(n57), .QN(N86) );
  NOR3X0 U68 ( .IN1(StateData[0]), .IN2(StatePreamble), .IN3(n11), .QN(
        ResetCollision) );
  NAND2X0 U69 ( .IN1(n58), .IN2(n59), .QN(n11) );
  INVX0 U70 ( .INP(StatePAD), .ZN(n58) );
  OR2X1 U71 ( .IN1(StartData[0]), .IN2(StartData[1]), .Q(N29) );
  AND3X1 U72 ( .IN1(n80), .IN2(ColWindow), .IN3(StartJam), .Q(
        MaxCollisionOccured) );
  INVX0 U73 ( .INP(n54), .ZN(n80) );
  NAND4X0 U74 ( .IN1(n60), .IN2(n61), .IN3(n62), .IN4(n63), .QN(n54) );
  XNOR2X1 U75 ( .IN1(RetryCnt[0]), .IN2(MaxRet[0]), .Q(n63) );
  XNOR2X1 U76 ( .IN1(RetryCnt[1]), .IN2(MaxRet[1]), .Q(n62) );
  XOR2X1 U77 ( .IN1(n95), .IN2(MaxRet[2]), .Q(n61) );
  XOR2X1 U78 ( .IN1(n33), .IN2(MaxRet[3]), .Q(n60) );
  NAND3X0 U79 ( .IN1(n64), .IN2(n65), .IN3(n66), .QN(MTxD_d[3]) );
  OA22X1 U80 ( .IN1(n46), .IN2(n67), .IN3(Crc[28]), .IN4(n68), .Q(n66) );
  INVX0 U81 ( .INP(NibCntEq15), .ZN(n46) );
  INVX0 U82 ( .INP(Data_Crc[0]), .ZN(n65) );
  NAND3X0 U83 ( .IN1(n67), .IN2(n69), .IN3(n70), .QN(MTxD_d[2]) );
  OR2X1 U84 ( .IN1(Crc[29]), .IN2(n68), .Q(n70) );
  INVX0 U85 ( .INP(Data_Crc[1]), .ZN(n69) );
  OAI21X1 U86 ( .IN1(Crc[30]), .IN2(n68), .IN3(n71), .QN(MTxD_d[1]) );
  INVX0 U87 ( .INP(Data_Crc[2]), .ZN(n71) );
  NAND4X0 U88 ( .IN1(n72), .IN2(n67), .IN3(n64), .IN4(n73), .QN(MTxD_d[0]) );
  INVX0 U89 ( .INP(Data_Crc[3]), .ZN(n73) );
  NAND3X0 U90 ( .IN1(n59), .IN2(n56), .IN3(StateJam), .QN(n64) );
  NAND4X0 U91 ( .IN1(StatePreamble), .IN2(n59), .IN3(n56), .IN4(n57), .QN(n67)
         );
  INVX0 U92 ( .INP(StateJam), .ZN(n57) );
  NOR2X0 U93 ( .IN1(StateFCS), .IN2(StateData[1]), .QN(n59) );
  OR2X1 U94 ( .IN1(Crc[31]), .IN2(n68), .Q(n72) );
  NAND3X0 U95 ( .IN1(n56), .IN2(n74), .IN3(StateFCS), .QN(n68) );
  INVX0 U96 ( .INP(StateData[0]), .ZN(n56) );
  NOR3X0 U97 ( .IN1(ColWindow), .IN2(UnderRun), .IN3(n45), .QN(LateCollision)
         );
  INVX0 U98 ( .INP(StartJam), .ZN(n45) );
  AND3X1 U99 ( .IN1(StateData[0]), .IN2(n12), .IN3(TxUnderRun), .Q(UnderRun)
         );
  INVX0 U100 ( .INP(Collision), .ZN(n12) );
  OR4X1 U101 ( .IN1(DlyCrcCnt[1]), .IN2(DlyCrcCnt[0]), .IN3(DlyCrcCnt[2]), 
        .IN4(n75), .Q(Initialize_Crc) );
  NAND2X0 U102 ( .IN1(n40), .IN2(n47), .QN(n75) );
  INVX0 U103 ( .INP(StatePreamble), .ZN(n47) );
  INVX0 U104 ( .INP(StateIdle), .ZN(n40) );
  AO22X1 U105 ( .IN1(TxData[0]), .IN2(StateData[0]), .IN3(TxData[4]), .IN4(n76), .Q(Data_Crc[3]) );
  AO22X1 U106 ( .IN1(TxData[1]), .IN2(StateData[0]), .IN3(TxData[5]), .IN4(n76), .Q(Data_Crc[2]) );
  AO22X1 U107 ( .IN1(TxData[2]), .IN2(StateData[0]), .IN3(TxData[6]), .IN4(n76), .Q(Data_Crc[1]) );
  AO22X1 U108 ( .IN1(TxData[3]), .IN2(StateData[0]), .IN3(TxData[7]), .IN4(n76), .Q(Data_Crc[0]) );
  NOR2X0 U109 ( .IN1(n74), .IN2(StateData[0]), .QN(n76) );
  INVX0 U110 ( .INP(StateData[1]), .ZN(n74) );
endmodule


module eth_rxstatem_test_1 ( MRxClk, Reset, MRxDV, ByteCntEq0, ByteCntGreat2, 
        Transmitting, MRxDEq5, MRxDEqD, IFGCounterEq24, ByteCntMaxFrame, 
        StateData, StateIdle, StatePreamble, StateSFD, StateDrop, 
        eth_top_test_point_11887_in, test_si, test_se );
  output [1:0] StateData;
  input MRxClk, Reset, MRxDV, ByteCntEq0, ByteCntGreat2, Transmitting, MRxDEq5,
         MRxDEqD, IFGCounterEq24, ByteCntMaxFrame, eth_top_test_point_11887_in,
         test_si, test_se;
  output StateIdle, StatePreamble, StateSFD, StateDrop;
  wire   n29, n30, n31, n32, n33, n34, n25, n26, n27, n28, n35, n36, n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19;

  SDFFASX1 StateDrop_reg ( .D(n34), .SI(StateData[1]), .SE(test_se), .CLK(
        MRxClk), .SETB(n19), .Q(StateDrop), .QN(n25) );
  SDFFARX1 StateIdle_reg ( .D(n33), .SI(StateDrop), .SE(test_se), .CLK(MRxClk), 
        .RSTB(n19), .Q(StateIdle), .QN(n28) );
  SDFFARX1 StatePreamble_reg ( .D(n32), .SI(StateIdle), .SE(test_se), .CLK(
        MRxClk), .RSTB(n19), .Q(StatePreamble), .QN(n27) );
  SDFFARX1 StateData1_reg ( .D(n31), .SI(StateData[0]), .SE(test_se), .CLK(
        MRxClk), .RSTB(n19), .Q(StateData[1]), .QN(n26) );
  SDFFARX1 StateData0_reg ( .D(n29), .SI(test_si), .SE(test_se), .CLK(MRxClk), 
        .RSTB(n19), .Q(StateData[0]), .QN(n36) );
  SDFFARX1 StateSFD_reg ( .D(n30), .SI(StatePreamble), .SE(test_se), .CLK(
        MRxClk), .RSTB(n19), .Q(StateSFD), .QN(n35) );
  INVX0 U2 ( .INP(eth_top_test_point_11887_in), .ZN(n19) );
  AOI21X1 U3 ( .IN1(n1), .IN2(n25), .IN3(n2), .QN(n34) );
  NAND2X0 U4 ( .IN1(n3), .IN2(MRxDV), .QN(n1) );
  AO21X1 U5 ( .IN1(n4), .IN2(StateIdle), .IN3(n2), .Q(n33) );
  INVX0 U6 ( .INP(n5), .ZN(n4) );
  MUX21X1 U7 ( .IN1(StatePreamble), .IN2(n6), .S(n5), .Q(n32) );
  AND2X1 U8 ( .IN1(n7), .IN2(n8), .Q(n6) );
  AND3X1 U9 ( .IN1(n9), .IN2(StateData[0]), .IN3(n8), .Q(n31) );
  NOR2X0 U10 ( .IN1(n10), .IN2(n11), .QN(n30) );
  OA22X1 U11 ( .IN1(n35), .IN2(n5), .IN3(n12), .IN4(n7), .Q(n10) );
  NAND3X0 U12 ( .IN1(n13), .IN2(n7), .IN3(n8), .QN(n5) );
  NAND3X0 U13 ( .IN1(MRxDV), .IN2(n14), .IN3(MRxDEq5), .QN(n7) );
  NAND2X0 U14 ( .IN1(n28), .IN2(n27), .QN(n14) );
  NAND2X0 U15 ( .IN1(MRxDV), .IN2(StateIdle), .QN(n13) );
  AND3X1 U16 ( .IN1(n8), .IN2(n11), .IN3(n36), .Q(n29) );
  INVX0 U17 ( .INP(n9), .ZN(n11) );
  OA21X1 U18 ( .IN1(n15), .IN2(n35), .IN3(n26), .Q(n9) );
  INVX0 U19 ( .INP(MRxDEqD), .ZN(n15) );
  INVX0 U20 ( .INP(n12), .ZN(n8) );
  AO21X1 U21 ( .IN1(MRxDV), .IN2(n3), .IN3(n2), .Q(n12) );
  NOR2X0 U22 ( .IN1(n16), .IN2(MRxDV), .QN(n2) );
  AND4X1 U23 ( .IN1(n36), .IN2(n35), .IN3(n17), .IN4(n27), .Q(n16) );
  AND2X1 U24 ( .IN1(n25), .IN2(n26), .Q(n17) );
  AO222X1 U25 ( .IN1(ByteCntMaxFrame), .IN2(StateData[0]), .IN3(n18), .IN4(
        MRxDEqD), .IN5(Transmitting), .IN6(StateIdle), .Q(n3) );
  NOR2X0 U26 ( .IN1(n35), .IN2(IFGCounterEq24), .QN(n18) );
endmodule


module eth_rxcounters_DW01_inc_1 ( A, SUM );
  input [15:0] A;
  output [15:0] SUM;

  wire   [15:2] carry;

  HADDX1 U1_1_14 ( .A0(A[14]), .B0(carry[14]), .C1(carry[15]), .SO(SUM[14]) );
  HADDX1 U1_1_13 ( .A0(A[13]), .B0(carry[13]), .C1(carry[14]), .SO(SUM[13]) );
  HADDX1 U1_1_12 ( .A0(A[12]), .B0(carry[12]), .C1(carry[13]), .SO(SUM[12]) );
  HADDX1 U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1 U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1 U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1 U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  XOR2X1 U2 ( .IN1(carry[15]), .IN2(A[15]), .Q(SUM[15]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module eth_rxcounters_test_1 ( MRxClk, Reset, MRxDV, StateIdle, StateSFD, 
        StateData, StateDrop, StatePreamble, MRxDEqD, DlyCrcEn, DlyCrcCnt, 
        Transmitting, MaxFL, r_IFG, HugEn, IFGCounterEq24, ByteCntEq0, 
        ByteCntEq1, ByteCntEq2, ByteCntEq3, ByteCntEq4, ByteCntEq5, ByteCntEq6, 
        ByteCntEq7, ByteCntGreat2, ByteCntSmall7, ByteCntMaxFrame, ByteCntOut, 
        eth_top_test_point_11887_in, test_si, test_so, test_se );
  input [1:0] StateData;
  output [3:0] DlyCrcCnt;
  input [15:0] MaxFL;
  output [15:0] ByteCntOut;
  input MRxClk, Reset, MRxDV, StateIdle, StateSFD, StateDrop, StatePreamble,
         MRxDEqD, DlyCrcEn, Transmitting, r_IFG, HugEn,
         eth_top_test_point_11887_in, test_si, test_se;
  output IFGCounterEq24, ByteCntEq0, ByteCntEq1, ByteCntEq2, ByteCntEq3,
         ByteCntEq4, ByteCntEq5, ByteCntEq6, ByteCntEq7, ByteCntGreat2,
         ByteCntSmall7, ByteCntMaxFrame, test_so;
  wire   N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20,
         N21, N22, n37, n38, n40, n41, n46, n47, n48, n49, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n1, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n175,
         n176, n177, n158, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n39, n42, n43, n44, n45,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n136;
  wire   [15:0] ByteCnt;

  SDFFARX1 \IFGCounter_reg[0]  ( .D(n118), .SI(DlyCrcCnt[3]), .SE(test_se), 
        .CLK(MRxClk), .RSTB(n136), .Q(n1), .QN(n160) );
  SDFFARX1 \IFGCounter_reg[3]  ( .D(n114), .SI(n176), .SE(test_se), .CLK(
        MRxClk), .RSTB(n136), .Q(n175), .QN(n132) );
  SDFFARX1 \IFGCounter_reg[1]  ( .D(n116), .SI(n1), .SE(test_se), .CLK(MRxClk), 
        .RSTB(n136), .Q(n177), .QN(n133) );
  SDFFARX1 \IFGCounter_reg[2]  ( .D(n115), .SI(n177), .SE(test_se), .CLK(
        MRxClk), .RSTB(n136), .Q(n176), .QN(n134) );
  SDFFARX1 \IFGCounter_reg[4]  ( .D(n117), .SI(n175), .SE(test_se), .CLK(
        MRxClk), .RSTB(n136), .Q(test_so) );
  SDFFARX1 \DlyCrcCnt_reg[0]  ( .D(n113), .SI(ByteCnt[15]), .SE(test_se), 
        .CLK(MRxClk), .RSTB(n136), .Q(DlyCrcCnt[0]), .QN(n49) );
  SDFFARX1 \DlyCrcCnt_reg[3]  ( .D(n112), .SI(DlyCrcCnt[2]), .SE(test_se), 
        .CLK(MRxClk), .RSTB(n136), .Q(DlyCrcCnt[3]), .QN(n46) );
  SDFFARX1 \ByteCnt_reg[14]  ( .D(n94), .SI(ByteCnt[13]), .SE(test_se), .CLK(
        MRxClk), .RSTB(n136), .Q(ByteCnt[14]), .QN(n168) );
  SDFFARX1 \ByteCnt_reg[15]  ( .D(n109), .SI(ByteCnt[14]), .SE(test_se), .CLK(
        MRxClk), .RSTB(n136), .Q(ByteCnt[15]), .QN(n169) );
  SDFFARX1 \ByteCnt_reg[13]  ( .D(n95), .SI(ByteCnt[12]), .SE(test_se), .CLK(
        MRxClk), .RSTB(n136), .Q(ByteCnt[13]), .QN(n167) );
  SDFFARX1 \ByteCnt_reg[12]  ( .D(n96), .SI(ByteCnt[11]), .SE(test_se), .CLK(
        MRxClk), .RSTB(n136), .Q(ByteCnt[12]), .QN(n166) );
  SDFFARX1 \ByteCnt_reg[11]  ( .D(n97), .SI(ByteCnt[10]), .SE(test_se), .CLK(
        MRxClk), .RSTB(n136), .Q(ByteCnt[11]), .QN(n171) );
  SDFFARX1 \ByteCnt_reg[10]  ( .D(n98), .SI(ByteCnt[9]), .SE(test_se), .CLK(
        MRxClk), .RSTB(n136), .Q(ByteCnt[10]), .QN(n170) );
  SDFFARX1 \ByteCnt_reg[9]  ( .D(n99), .SI(ByteCnt[8]), .SE(test_se), .CLK(
        MRxClk), .RSTB(n136), .Q(ByteCnt[9]), .QN(n158) );
  SDFFARX1 \ByteCnt_reg[8]  ( .D(n100), .SI(ByteCnt[7]), .SE(test_se), .CLK(
        MRxClk), .RSTB(n136), .Q(ByteCnt[8]), .QN(n163) );
  SDFFARX1 \ByteCnt_reg[7]  ( .D(n101), .SI(ByteCnt[6]), .SE(test_se), .CLK(
        MRxClk), .RSTB(n136), .Q(ByteCnt[7]), .QN(n165) );
  SDFFARX1 \ByteCnt_reg[6]  ( .D(n102), .SI(ByteCnt[5]), .SE(test_se), .CLK(
        MRxClk), .RSTB(n136), .Q(ByteCnt[6]), .QN(n164) );
  SDFFARX1 \ByteCnt_reg[5]  ( .D(n103), .SI(ByteCnt[4]), .SE(test_se), .CLK(
        MRxClk), .RSTB(n136), .Q(ByteCnt[5]), .QN(n162) );
  SDFFARX1 \ByteCnt_reg[4]  ( .D(n104), .SI(ByteCnt[3]), .SE(test_se), .CLK(
        MRxClk), .RSTB(n136), .Q(ByteCnt[4]), .QN(n161) );
  SDFFARX1 \ByteCnt_reg[3]  ( .D(n105), .SI(ByteCnt[2]), .SE(test_se), .CLK(
        MRxClk), .RSTB(n136), .Q(ByteCnt[3]), .QN(n37) );
  SDFFARX1 \ByteCnt_reg[2]  ( .D(n106), .SI(ByteCntOut[1]), .SE(test_se), 
        .CLK(MRxClk), .RSTB(n136), .Q(ByteCnt[2]), .QN(n38) );
  SDFFARX1 \ByteCnt_reg[1]  ( .D(n107), .SI(ByteCntOut[0]), .SE(test_se), 
        .CLK(MRxClk), .RSTB(n136), .Q(ByteCntOut[1]), .QN(n40) );
  SDFFARX1 \ByteCnt_reg[0]  ( .D(n108), .SI(test_si), .SE(test_se), .CLK(
        MRxClk), .RSTB(n136), .Q(ByteCntOut[0]), .QN(n41) );
  SDFFARX1 \DlyCrcCnt_reg[2]  ( .D(n110), .SI(DlyCrcCnt[1]), .SE(test_se), 
        .CLK(MRxClk), .RSTB(n136), .Q(DlyCrcCnt[2]), .QN(n47) );
  SDFFARX1 \DlyCrcCnt_reg[1]  ( .D(n111), .SI(DlyCrcCnt[0]), .SE(test_se), 
        .CLK(MRxClk), .RSTB(n136), .Q(DlyCrcCnt[1]), .QN(n48) );
  eth_rxcounters_DW01_inc_1 add_159 ( .A({ByteCnt[15:2], ByteCntOut[1:0]}), 
        .SUM({N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, 
        N9, N8, N7}) );
  INVX0 U3 ( .INP(n2), .ZN(IFGCounterEq24) );
  INVX0 U4 ( .INP(eth_top_test_point_11887_in), .ZN(n136) );
  AO22X1 U5 ( .IN1(N16), .IN2(n3), .IN3(n4), .IN4(ByteCnt[9]), .Q(n99) );
  AO22X1 U6 ( .IN1(N17), .IN2(n3), .IN3(n4), .IN4(ByteCnt[10]), .Q(n98) );
  AO22X1 U7 ( .IN1(N18), .IN2(n3), .IN3(n4), .IN4(ByteCnt[11]), .Q(n97) );
  AO22X1 U8 ( .IN1(N19), .IN2(n3), .IN3(n4), .IN4(ByteCnt[12]), .Q(n96) );
  AO22X1 U9 ( .IN1(N20), .IN2(n3), .IN3(n4), .IN4(ByteCnt[13]), .Q(n95) );
  AO22X1 U10 ( .IN1(N21), .IN2(n3), .IN3(n4), .IN4(ByteCnt[14]), .Q(n94) );
  MUX21X1 U11 ( .IN1(n5), .IN2(n6), .S(n1), .Q(n118) );
  MUX21X1 U12 ( .IN1(n7), .IN2(n8), .S(test_so), .Q(n117) );
  AO21X1 U13 ( .IN1(n132), .IN2(n5), .IN3(n9), .Q(n8) );
  NOR3X0 U14 ( .IN1(n10), .IN2(n132), .IN3(n11), .QN(n7) );
  MUX21X1 U15 ( .IN1(n12), .IN2(n13), .S(n133), .Q(n116) );
  NOR2X0 U16 ( .IN1(n160), .IN2(n11), .QN(n13) );
  MUX21X1 U17 ( .IN1(n14), .IN2(n15), .S(n176), .Q(n115) );
  AO21X1 U18 ( .IN1(n5), .IN2(n133), .IN3(n12), .Q(n15) );
  AO21X1 U19 ( .IN1(n5), .IN2(n160), .IN3(n6), .Q(n12) );
  NOR3X0 U20 ( .IN1(n11), .IN2(n133), .IN3(n160), .QN(n14) );
  MUX21X1 U21 ( .IN1(n9), .IN2(n16), .S(n132), .Q(n114) );
  NOR2X0 U22 ( .IN1(n11), .IN2(n10), .QN(n16) );
  AO21X1 U23 ( .IN1(n5), .IN2(n10), .IN3(n6), .Q(n9) );
  AND3X1 U24 ( .IN1(n17), .IN2(n18), .IN3(n11), .Q(n6) );
  OR3X1 U25 ( .IN1(n134), .IN2(n133), .IN3(n160), .Q(n10) );
  INVX0 U26 ( .INP(n11), .ZN(n5) );
  NAND4X0 U27 ( .IN1(n19), .IN2(n17), .IN3(n2), .IN4(n18), .QN(n11) );
  INVX0 U28 ( .INP(StateDrop), .ZN(n18) );
  NOR2X0 U29 ( .IN1(n20), .IN2(r_IFG), .QN(n2) );
  NOR4X0 U30 ( .IN1(n21), .IN2(n176), .IN3(n132), .IN4(n1), .QN(n20) );
  NAND2X0 U31 ( .IN1(test_so), .IN2(n133), .QN(n21) );
  NAND3X0 U32 ( .IN1(n22), .IN2(n23), .IN3(n24), .QN(n19) );
  AO21X1 U33 ( .IN1(n25), .IN2(n26), .IN3(n27), .Q(n113) );
  MUX21X1 U34 ( .IN1(n28), .IN2(n29), .S(DlyCrcCnt[0]), .Q(n27) );
  MUX21X1 U35 ( .IN1(n30), .IN2(n31), .S(DlyCrcCnt[3]), .Q(n112) );
  AO21X1 U36 ( .IN1(n28), .IN2(n47), .IN3(n32), .Q(n31) );
  NOR2X0 U37 ( .IN1(n47), .IN2(n33), .QN(n30) );
  INVX0 U38 ( .INP(n34), .ZN(n33) );
  MUX21X1 U39 ( .IN1(n35), .IN2(n36), .S(n48), .Q(n111) );
  NOR2X0 U40 ( .IN1(n49), .IN2(n39), .QN(n36) );
  MUX21X1 U41 ( .IN1(n32), .IN2(n34), .S(n47), .Q(n110) );
  NOR3X0 U42 ( .IN1(n48), .IN2(n49), .IN3(n39), .QN(n34) );
  AO21X1 U43 ( .IN1(n28), .IN2(n48), .IN3(n35), .Q(n32) );
  AO21X1 U44 ( .IN1(n28), .IN2(n49), .IN3(n29), .Q(n35) );
  AND3X1 U45 ( .IN1(n42), .IN2(n26), .IN3(n39), .Q(n29) );
  INVX0 U46 ( .INP(n39), .ZN(n28) );
  NAND3X0 U47 ( .IN1(n42), .IN2(n26), .IN3(n43), .QN(n39) );
  INVX0 U48 ( .INP(n44), .ZN(n43) );
  NAND4X0 U49 ( .IN1(n48), .IN2(n47), .IN3(DlyCrcCnt[3]), .IN4(DlyCrcCnt[0]), 
        .QN(n26) );
  INVX0 U50 ( .INP(n25), .ZN(n42) );
  NOR2X0 U51 ( .IN1(n45), .IN2(n23), .QN(n25) );
  AO22X1 U52 ( .IN1(N22), .IN2(n3), .IN3(n4), .IN4(ByteCnt[15]), .Q(n109) );
  AO22X1 U53 ( .IN1(N7), .IN2(n3), .IN3(n4), .IN4(ByteCntOut[0]), .Q(n108) );
  AO22X1 U54 ( .IN1(N8), .IN2(n3), .IN3(n4), .IN4(ByteCntOut[1]), .Q(n107) );
  AO22X1 U55 ( .IN1(N9), .IN2(n3), .IN3(n4), .IN4(ByteCnt[2]), .Q(n106) );
  AO22X1 U56 ( .IN1(N10), .IN2(n3), .IN3(n4), .IN4(ByteCnt[3]), .Q(n105) );
  AO22X1 U57 ( .IN1(N11), .IN2(n3), .IN3(n4), .IN4(ByteCnt[4]), .Q(n104) );
  AO22X1 U58 ( .IN1(N12), .IN2(n3), .IN3(n4), .IN4(ByteCnt[5]), .Q(n103) );
  AO22X1 U59 ( .IN1(N13), .IN2(n3), .IN3(n4), .IN4(ByteCnt[6]), .Q(n102) );
  AO22X1 U60 ( .IN1(N14), .IN2(n3), .IN3(n4), .IN4(ByteCnt[7]), .Q(n101) );
  AO22X1 U61 ( .IN1(N15), .IN2(n3), .IN3(n4), .IN4(ByteCnt[8]), .Q(n100) );
  AND3X1 U62 ( .IN1(n50), .IN2(n17), .IN3(n51), .Q(n4) );
  NAND3X0 U63 ( .IN1(ByteCntMaxFrame), .IN2(MRxDV), .IN3(StateData[0]), .QN(
        n51) );
  INVX0 U64 ( .INP(n50), .ZN(n3) );
  NAND4X0 U65 ( .IN1(MRxDV), .IN2(n52), .IN3(n53), .IN4(n17), .QN(n50) );
  NAND3X0 U66 ( .IN1(MRxDV), .IN2(MRxDEqD), .IN3(StateSFD), .QN(n17) );
  NAND4X0 U67 ( .IN1(n54), .IN2(n55), .IN3(n22), .IN4(n23), .QN(n53) );
  INVX0 U68 ( .INP(StateSFD), .ZN(n23) );
  INVX0 U69 ( .INP(StatePreamble), .ZN(n22) );
  NAND3X0 U70 ( .IN1(n56), .IN2(n44), .IN3(StateData[1]), .QN(n55) );
  NAND2X0 U71 ( .IN1(DlyCrcEn), .IN2(n57), .QN(n44) );
  NAND4X0 U72 ( .IN1(n49), .IN2(n48), .IN3(n47), .IN4(n46), .QN(n57) );
  NAND4X0 U73 ( .IN1(n58), .IN2(n59), .IN3(n60), .IN4(n61), .QN(n56) );
  NOR4X0 U74 ( .IN1(n62), .IN2(n166), .IN3(n168), .IN4(n167), .QN(n61) );
  NAND4X0 U75 ( .IN1(ByteCnt[15]), .IN2(ByteCnt[10]), .IN3(ByteCnt[11]), .IN4(
        ByteCnt[3]), .QN(n62) );
  NOR4X0 U76 ( .IN1(n165), .IN2(n164), .IN3(n163), .IN4(n162), .QN(n60) );
  NOR2X0 U77 ( .IN1(n161), .IN2(n158), .QN(n58) );
  OR2X1 U78 ( .IN1(Transmitting), .IN2(n24), .Q(n54) );
  INVX0 U79 ( .INP(StateIdle), .ZN(n24) );
  NAND2X0 U80 ( .IN1(StateData[0]), .IN2(ByteCntMaxFrame), .QN(n52) );
  NOR2X0 U81 ( .IN1(n59), .IN2(n63), .QN(ByteCntSmall7) );
  INVX0 U82 ( .INP(n64), .ZN(n59) );
  XNOR2X1 U83 ( .IN1(n158), .IN2(n65), .Q(ByteCntOut[9]) );
  XNOR2X1 U84 ( .IN1(n66), .IN2(ByteCnt[8]), .Q(ByteCntOut[8]) );
  XNOR2X1 U85 ( .IN1(n165), .IN2(n67), .Q(ByteCntOut[7]) );
  XNOR2X1 U86 ( .IN1(n68), .IN2(ByteCnt[6]), .Q(ByteCntOut[6]) );
  XNOR2X1 U87 ( .IN1(n69), .IN2(ByteCnt[5]), .Q(ByteCntOut[5]) );
  NAND2X0 U88 ( .IN1(n70), .IN2(ByteCnt[4]), .QN(n69) );
  XNOR2X1 U89 ( .IN1(n161), .IN2(n70), .Q(ByteCntOut[4]) );
  XNOR2X1 U90 ( .IN1(n37), .IN2(n71), .Q(ByteCntOut[3]) );
  NOR2X0 U91 ( .IN1(n38), .IN2(n45), .QN(n71) );
  INVX0 U92 ( .INP(DlyCrcEn), .ZN(n45) );
  XNOR2X1 U93 ( .IN1(DlyCrcEn), .IN2(n38), .Q(ByteCntOut[2]) );
  XNOR2X1 U94 ( .IN1(n169), .IN2(n72), .Q(ByteCntOut[15]) );
  NOR2X0 U95 ( .IN1(n168), .IN2(n73), .QN(n72) );
  XNOR2X1 U96 ( .IN1(n73), .IN2(ByteCnt[14]), .Q(ByteCntOut[14]) );
  NAND3X0 U97 ( .IN1(ByteCnt[12]), .IN2(ByteCnt[13]), .IN3(n74), .QN(n73) );
  XNOR2X1 U98 ( .IN1(n75), .IN2(ByteCnt[13]), .Q(ByteCntOut[13]) );
  NAND2X0 U99 ( .IN1(n74), .IN2(ByteCnt[12]), .QN(n75) );
  XNOR2X1 U100 ( .IN1(n166), .IN2(n74), .Q(ByteCntOut[12]) );
  NOR3X0 U101 ( .IN1(n170), .IN2(n171), .IN3(n76), .QN(n74) );
  XNOR2X1 U102 ( .IN1(n171), .IN2(n77), .Q(ByteCntOut[11]) );
  NOR2X0 U103 ( .IN1(n170), .IN2(n76), .QN(n77) );
  XNOR2X1 U104 ( .IN1(n76), .IN2(ByteCnt[10]), .Q(ByteCntOut[10]) );
  NAND2X0 U105 ( .IN1(n65), .IN2(ByteCnt[9]), .QN(n76) );
  NOR2X0 U106 ( .IN1(n66), .IN2(n163), .QN(n65) );
  NAND2X0 U107 ( .IN1(n67), .IN2(ByteCnt[7]), .QN(n66) );
  NOR2X0 U108 ( .IN1(n68), .IN2(n164), .QN(n67) );
  NAND3X0 U109 ( .IN1(ByteCnt[4]), .IN2(ByteCnt[5]), .IN3(n70), .QN(n68) );
  AND3X1 U110 ( .IN1(ByteCnt[3]), .IN2(ByteCnt[2]), .IN3(DlyCrcEn), .Q(n70) );
  NOR4X0 U111 ( .IN1(n78), .IN2(n79), .IN3(n80), .IN4(n81), .QN(
        ByteCntMaxFrame) );
  NAND4X0 U112 ( .IN1(n82), .IN2(n83), .IN3(n84), .IN4(n85), .QN(n81) );
  XNOR2X1 U113 ( .IN1(ByteCnt[15]), .IN2(MaxFL[15]), .Q(n85) );
  XNOR2X1 U114 ( .IN1(ByteCnt[3]), .IN2(MaxFL[3]), .Q(n84) );
  XNOR2X1 U115 ( .IN1(ByteCnt[4]), .IN2(MaxFL[4]), .Q(n83) );
  XNOR2X1 U116 ( .IN1(ByteCnt[5]), .IN2(MaxFL[5]), .Q(n82) );
  NAND4X0 U117 ( .IN1(n86), .IN2(n87), .IN3(n88), .IN4(n89), .QN(n80) );
  XNOR2X1 U118 ( .IN1(ByteCntOut[0]), .IN2(MaxFL[0]), .Q(n89) );
  NOR2X0 U119 ( .IN1(HugEn), .IN2(n90), .QN(n88) );
  XNOR2X1 U120 ( .IN1(n40), .IN2(MaxFL[1]), .Q(n90) );
  XNOR2X1 U121 ( .IN1(ByteCnt[2]), .IN2(MaxFL[2]), .Q(n87) );
  XNOR2X1 U122 ( .IN1(ByteCnt[6]), .IN2(MaxFL[6]), .Q(n86) );
  NAND4X0 U123 ( .IN1(n91), .IN2(n92), .IN3(n93), .IN4(n119), .QN(n79) );
  XNOR2X1 U124 ( .IN1(ByteCnt[11]), .IN2(MaxFL[11]), .Q(n119) );
  XNOR2X1 U125 ( .IN1(ByteCnt[12]), .IN2(MaxFL[12]), .Q(n93) );
  XNOR2X1 U126 ( .IN1(ByteCnt[13]), .IN2(MaxFL[13]), .Q(n92) );
  XNOR2X1 U127 ( .IN1(ByteCnt[14]), .IN2(MaxFL[14]), .Q(n91) );
  NAND4X0 U128 ( .IN1(n120), .IN2(n121), .IN3(n122), .IN4(n123), .QN(n78) );
  XNOR2X1 U129 ( .IN1(ByteCnt[10]), .IN2(MaxFL[10]), .Q(n123) );
  XNOR2X1 U130 ( .IN1(ByteCnt[7]), .IN2(MaxFL[7]), .Q(n122) );
  XNOR2X1 U131 ( .IN1(ByteCnt[8]), .IN2(MaxFL[8]), .Q(n121) );
  XNOR2X1 U132 ( .IN1(ByteCnt[9]), .IN2(MaxFL[9]), .Q(n120) );
  NAND3X0 U133 ( .IN1(n38), .IN2(n124), .IN3(n125), .QN(ByteCntGreat2) );
  NAND2X0 U134 ( .IN1(ByteCntOut[1]), .IN2(ByteCntOut[0]), .QN(n124) );
  NOR2X0 U135 ( .IN1(n64), .IN2(n63), .QN(ByteCntEq7) );
  NAND3X0 U136 ( .IN1(ByteCntOut[1]), .IN2(ByteCntOut[0]), .IN3(ByteCnt[2]), 
        .QN(n64) );
  NOR3X0 U137 ( .IN1(n126), .IN2(n40), .IN3(n38), .QN(ByteCntEq6) );
  NOR2X0 U138 ( .IN1(n38), .IN2(n127), .QN(ByteCntEq5) );
  NOR3X0 U139 ( .IN1(n126), .IN2(n38), .IN3(ByteCntOut[1]), .QN(ByteCntEq4) );
  NOR4X0 U140 ( .IN1(n41), .IN2(n40), .IN3(ByteCnt[2]), .IN4(n63), .QN(
        ByteCntEq3) );
  NOR3X0 U141 ( .IN1(n126), .IN2(n40), .IN3(ByteCnt[2]), .QN(ByteCntEq2) );
  NOR2X0 U142 ( .IN1(ByteCnt[2]), .IN2(n127), .QN(ByteCntEq1) );
  NAND3X0 U143 ( .IN1(n40), .IN2(ByteCntOut[0]), .IN3(n125), .QN(n127) );
  NOR3X0 U144 ( .IN1(n126), .IN2(ByteCntOut[1]), .IN3(ByteCnt[2]), .QN(
        ByteCntEq0) );
  NAND2X0 U145 ( .IN1(n125), .IN2(n41), .QN(n126) );
  INVX0 U146 ( .INP(n63), .ZN(n125) );
  NAND4X0 U147 ( .IN1(n128), .IN2(n168), .IN3(n129), .IN4(n130), .QN(n63) );
  NOR4X0 U148 ( .IN1(n131), .IN2(ByteCnt[7]), .IN3(ByteCnt[5]), .IN4(
        ByteCnt[10]), .QN(n130) );
  NAND4X0 U149 ( .IN1(n161), .IN2(n37), .IN3(n169), .IN4(n164), .QN(n131) );
  NOR3X0 U150 ( .IN1(ByteCnt[9]), .IN2(ByteCnt[8]), .IN3(ByteCnt[11]), .QN(
        n129) );
  NOR2X0 U151 ( .IN1(ByteCnt[12]), .IN2(ByteCnt[13]), .QN(n128) );
endmodule


module eth_rxaddrcheck_test_1 ( MRxClk, Reset, RxData, Broadcast, r_Bro, r_Pro, 
        ByteCntEq2, ByteCntEq3, ByteCntEq4, ByteCntEq5, ByteCntEq6, ByteCntEq7, 
        HASH0, HASH1, CrcHash, CrcHashGood, StateData, RxEndFrm, Multicast, 
        MAC, RxAbort, AddressMiss, PassAll, ControlFrmAddressOK, 
        eth_top_test_point_11887_in, test_si, test_so, test_se );
  input [7:0] RxData;
  input [31:0] HASH0;
  input [31:0] HASH1;
  input [5:0] CrcHash;
  input [1:0] StateData;
  input [47:0] MAC;
  input MRxClk, Reset, Broadcast, r_Bro, r_Pro, ByteCntEq2, ByteCntEq3,
         ByteCntEq4, ByteCntEq5, ByteCntEq6, ByteCntEq7, CrcHashGood, RxEndFrm,
         Multicast, PassAll, ControlFrmAddressOK, eth_top_test_point_11887_in,
         test_si, test_se;
  output RxAbort, AddressMiss, test_so;
  wire   N7, N8, N9, N10, n102, n109, n110, n119, n120, n133, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n103,
         n104, n105, n106, n107, n108, n111, n112, n113, n114, n115, n116,
         n117, n118, n121, n122, n123, n124, n125, n126;
  assign N7 = CrcHash[0];
  assign N8 = CrcHash[1];
  assign N9 = CrcHash[2];
  assign test_so = n120;

  SDFFARX1 UnicastOK_reg ( .D(n110), .SI(RxAbort), .SE(test_se), .CLK(MRxClk), 
        .RSTB(n126), .Q(n120), .QN(n133) );
  SDFFARX1 RxAbort_reg ( .D(N10), .SI(n119), .SE(test_se), .CLK(MRxClk), 
        .RSTB(n126), .Q(RxAbort), .QN(n125) );
  SDFFARX1 MulticastOK_reg ( .D(n109), .SI(AddressMiss), .SE(test_se), .CLK(
        MRxClk), .RSTB(n126), .Q(n119) );
  SDFFARX1 AddressMiss_reg ( .D(n102), .SI(test_si), .SE(test_se), .CLK(MRxClk), .RSTB(n126), .Q(AddressMiss) );
  INVX0 U3 ( .INP(eth_top_test_point_11887_in), .ZN(n126) );
  NAND2X0 U4 ( .IN1(n1), .IN2(n2), .QN(n110) );
  NAND4X0 U5 ( .IN1(n125), .IN2(n3), .IN3(n4), .IN4(n5), .QN(n2) );
  NOR2X0 U6 ( .IN1(n133), .IN2(RxEndFrm), .QN(n4) );
  OR4X1 U7 ( .IN1(n6), .IN2(n7), .IN3(n8), .IN4(n9), .Q(n1) );
  NAND4X0 U8 ( .IN1(n10), .IN2(n11), .IN3(n12), .IN4(n13), .QN(n9) );
  XOR2X1 U9 ( .IN1(RxData[0]), .IN2(n14), .Q(n13) );
  NOR2X0 U10 ( .IN1(n15), .IN2(n16), .QN(n14) );
  AO222X1 U11 ( .IN1(MAC[8]), .IN2(n17), .IN3(MAC[24]), .IN4(n18), .IN5(
        MAC[40]), .IN6(n19), .Q(n16) );
  AO222X1 U12 ( .IN1(MAC[0]), .IN2(n3), .IN3(MAC[32]), .IN4(n20), .IN5(MAC[16]), .IN6(n21), .Q(n15) );
  OA21X1 U13 ( .IN1(n19), .IN2(n120), .IN3(n22), .Q(n12) );
  NAND4X0 U14 ( .IN1(n23), .IN2(n24), .IN3(n25), .IN4(n5), .QN(n22) );
  OAI21X1 U15 ( .IN1(ByteCntEq4), .IN2(ByteCntEq6), .IN3(n26), .QN(n24) );
  XOR2X1 U16 ( .IN1(RxData[1]), .IN2(n27), .Q(n11) );
  NOR2X0 U17 ( .IN1(n28), .IN2(n29), .QN(n27) );
  AO222X1 U18 ( .IN1(MAC[9]), .IN2(n17), .IN3(MAC[25]), .IN4(n18), .IN5(
        MAC[41]), .IN6(n19), .Q(n29) );
  AO222X1 U19 ( .IN1(MAC[1]), .IN2(n3), .IN3(MAC[33]), .IN4(n20), .IN5(MAC[17]), .IN6(n21), .Q(n28) );
  XOR2X1 U20 ( .IN1(RxData[2]), .IN2(n30), .Q(n10) );
  NOR2X0 U21 ( .IN1(n31), .IN2(n32), .QN(n30) );
  AO222X1 U22 ( .IN1(MAC[10]), .IN2(n17), .IN3(MAC[26]), .IN4(n18), .IN5(
        MAC[42]), .IN6(n19), .Q(n32) );
  AO222X1 U23 ( .IN1(MAC[2]), .IN2(n3), .IN3(MAC[34]), .IN4(n20), .IN5(MAC[18]), .IN6(n21), .Q(n31) );
  NAND3X0 U24 ( .IN1(n33), .IN2(n34), .IN3(n35), .QN(n8) );
  XOR2X1 U25 ( .IN1(RxData[4]), .IN2(n36), .Q(n35) );
  NOR2X0 U26 ( .IN1(n37), .IN2(n38), .QN(n36) );
  AO222X1 U27 ( .IN1(MAC[12]), .IN2(n17), .IN3(MAC[28]), .IN4(n18), .IN5(
        MAC[44]), .IN6(n19), .Q(n38) );
  AO222X1 U28 ( .IN1(MAC[4]), .IN2(n3), .IN3(MAC[36]), .IN4(n20), .IN5(MAC[20]), .IN6(n21), .Q(n37) );
  XOR2X1 U29 ( .IN1(RxData[5]), .IN2(n39), .Q(n34) );
  NOR2X0 U30 ( .IN1(n40), .IN2(n41), .QN(n39) );
  AO222X1 U31 ( .IN1(MAC[13]), .IN2(n17), .IN3(MAC[29]), .IN4(n18), .IN5(
        MAC[45]), .IN6(n19), .Q(n41) );
  AO222X1 U32 ( .IN1(MAC[5]), .IN2(n3), .IN3(MAC[37]), .IN4(n20), .IN5(MAC[21]), .IN6(n21), .Q(n40) );
  XOR2X1 U33 ( .IN1(RxData[3]), .IN2(n42), .Q(n33) );
  NOR2X0 U34 ( .IN1(n43), .IN2(n44), .QN(n42) );
  AO222X1 U35 ( .IN1(MAC[11]), .IN2(n17), .IN3(MAC[27]), .IN4(n18), .IN5(
        MAC[43]), .IN6(n19), .Q(n44) );
  AO222X1 U36 ( .IN1(MAC[3]), .IN2(n3), .IN3(MAC[35]), .IN4(n20), .IN5(MAC[19]), .IN6(n21), .Q(n43) );
  XNOR2X1 U37 ( .IN1(RxData[7]), .IN2(n45), .Q(n7) );
  NOR2X0 U38 ( .IN1(n46), .IN2(n47), .QN(n45) );
  AO222X1 U39 ( .IN1(MAC[15]), .IN2(n17), .IN3(MAC[31]), .IN4(n18), .IN5(
        MAC[47]), .IN6(n19), .Q(n47) );
  AO222X1 U40 ( .IN1(MAC[7]), .IN2(n3), .IN3(MAC[39]), .IN4(n20), .IN5(MAC[23]), .IN6(n21), .Q(n46) );
  XNOR2X1 U41 ( .IN1(RxData[6]), .IN2(n48), .Q(n6) );
  NOR2X0 U42 ( .IN1(n49), .IN2(n50), .QN(n48) );
  AO222X1 U43 ( .IN1(MAC[14]), .IN2(n17), .IN3(MAC[30]), .IN4(n18), .IN5(
        MAC[46]), .IN6(n19), .Q(n50) );
  NOR2X0 U44 ( .IN1(n51), .IN2(n52), .QN(n18) );
  NOR3X0 U45 ( .IN1(n53), .IN2(n54), .IN3(n55), .QN(n17) );
  INVX0 U46 ( .INP(n25), .ZN(n54) );
  AO222X1 U47 ( .IN1(MAC[6]), .IN2(n3), .IN3(MAC[38]), .IN4(n20), .IN5(MAC[22]), .IN6(n21), .Q(n49) );
  NOR2X0 U48 ( .IN1(n25), .IN2(n53), .QN(n21) );
  INVX0 U49 ( .INP(n56), .ZN(n53) );
  AND2X1 U50 ( .IN1(ByteCntEq3), .IN2(n57), .Q(n20) );
  AND3X1 U51 ( .IN1(n55), .IN2(n25), .IN3(n56), .Q(n3) );
  OA21X1 U52 ( .IN1(n52), .IN2(n58), .IN3(n23), .Q(n56) );
  INVX0 U53 ( .INP(n51), .ZN(n23) );
  AO21X1 U54 ( .IN1(ByteCntEq3), .IN2(n26), .IN3(n19), .Q(n51) );
  INVX0 U55 ( .INP(n57), .ZN(n19) );
  NAND2X0 U56 ( .IN1(ByteCntEq2), .IN2(n26), .QN(n57) );
  INVX0 U57 ( .INP(ByteCntEq4), .ZN(n52) );
  NAND2X0 U58 ( .IN1(ByteCntEq5), .IN2(n26), .QN(n25) );
  NAND2X0 U59 ( .IN1(ByteCntEq6), .IN2(n26), .QN(n55) );
  AND3X1 U60 ( .IN1(n125), .IN2(n59), .IN3(n60), .Q(n109) );
  MUX21X1 U61 ( .IN1(n119), .IN2(n61), .S(n62), .Q(n60) );
  AND2X1 U62 ( .IN1(Multicast), .IN2(CrcHashGood), .Q(n62) );
  MUX41X1 U63 ( .IN1(n63), .IN3(n64), .IN2(n65), .IN4(n66), .S0(N9), .S1(N8), 
        .Q(n61) );
  AO221X1 U64 ( .IN1(n67), .IN2(n68), .IN3(n69), .IN4(n70), .IN5(n71), .Q(n66)
         );
  AO22X1 U65 ( .IN1(n72), .IN2(n73), .IN3(n74), .IN4(n75), .Q(n71) );
  AO221X1 U66 ( .IN1(HASH0[22]), .IN2(n76), .IN3(HASH0[30]), .IN4(n77), .IN5(
        n78), .Q(n75) );
  AO22X1 U67 ( .IN1(HASH0[14]), .IN2(n79), .IN3(HASH0[6]), .IN4(n80), .Q(n78)
         );
  AO221X1 U68 ( .IN1(HASH1[22]), .IN2(n76), .IN3(HASH1[30]), .IN4(n77), .IN5(
        n81), .Q(n73) );
  AO22X1 U69 ( .IN1(HASH1[14]), .IN2(n79), .IN3(HASH1[6]), .IN4(n80), .Q(n81)
         );
  AO221X1 U70 ( .IN1(HASH0[23]), .IN2(n76), .IN3(HASH0[31]), .IN4(n77), .IN5(
        n82), .Q(n70) );
  AO22X1 U71 ( .IN1(HASH0[15]), .IN2(n79), .IN3(HASH0[7]), .IN4(n80), .Q(n82)
         );
  AO221X1 U72 ( .IN1(HASH1[23]), .IN2(n76), .IN3(HASH1[31]), .IN4(n77), .IN5(
        n83), .Q(n68) );
  AO22X1 U73 ( .IN1(HASH1[15]), .IN2(n79), .IN3(HASH1[7]), .IN4(n80), .Q(n83)
         );
  AO221X1 U74 ( .IN1(n67), .IN2(n84), .IN3(n69), .IN4(n85), .IN5(n86), .Q(n65)
         );
  AO22X1 U75 ( .IN1(n72), .IN2(n87), .IN3(n74), .IN4(n88), .Q(n86) );
  AO221X1 U76 ( .IN1(HASH0[18]), .IN2(n76), .IN3(HASH0[26]), .IN4(n77), .IN5(
        n89), .Q(n88) );
  AO22X1 U77 ( .IN1(HASH0[10]), .IN2(n79), .IN3(HASH0[2]), .IN4(n80), .Q(n89)
         );
  AO221X1 U78 ( .IN1(HASH1[18]), .IN2(n76), .IN3(HASH1[26]), .IN4(n77), .IN5(
        n90), .Q(n87) );
  AO22X1 U79 ( .IN1(HASH1[10]), .IN2(n79), .IN3(HASH1[2]), .IN4(n80), .Q(n90)
         );
  AO221X1 U80 ( .IN1(HASH0[19]), .IN2(n76), .IN3(HASH0[27]), .IN4(n77), .IN5(
        n91), .Q(n85) );
  AO22X1 U81 ( .IN1(HASH0[11]), .IN2(n79), .IN3(HASH0[3]), .IN4(n80), .Q(n91)
         );
  AO221X1 U82 ( .IN1(HASH1[19]), .IN2(n76), .IN3(HASH1[27]), .IN4(n77), .IN5(
        n92), .Q(n84) );
  AO22X1 U83 ( .IN1(HASH1[11]), .IN2(n79), .IN3(HASH1[3]), .IN4(n80), .Q(n92)
         );
  AO221X1 U84 ( .IN1(n67), .IN2(n93), .IN3(n69), .IN4(n94), .IN5(n95), .Q(n64)
         );
  AO22X1 U85 ( .IN1(n72), .IN2(n96), .IN3(n74), .IN4(n97), .Q(n95) );
  AO221X1 U86 ( .IN1(HASH0[20]), .IN2(n76), .IN3(HASH0[28]), .IN4(n77), .IN5(
        n98), .Q(n97) );
  AO22X1 U87 ( .IN1(HASH0[12]), .IN2(n79), .IN3(HASH0[4]), .IN4(n80), .Q(n98)
         );
  AO221X1 U88 ( .IN1(HASH1[20]), .IN2(n76), .IN3(HASH1[28]), .IN4(n77), .IN5(
        n99), .Q(n96) );
  AO22X1 U89 ( .IN1(HASH1[12]), .IN2(n79), .IN3(HASH1[4]), .IN4(n80), .Q(n99)
         );
  AO221X1 U90 ( .IN1(HASH0[21]), .IN2(n76), .IN3(HASH0[29]), .IN4(n77), .IN5(
        n100), .Q(n94) );
  AO22X1 U91 ( .IN1(HASH0[13]), .IN2(n79), .IN3(HASH0[5]), .IN4(n80), .Q(n100)
         );
  AO221X1 U92 ( .IN1(HASH1[21]), .IN2(n76), .IN3(HASH1[29]), .IN4(n77), .IN5(
        n101), .Q(n93) );
  AO22X1 U93 ( .IN1(HASH1[13]), .IN2(n79), .IN3(HASH1[5]), .IN4(n80), .Q(n101)
         );
  AO221X1 U94 ( .IN1(n67), .IN2(n103), .IN3(n69), .IN4(n104), .IN5(n105), .Q(
        n63) );
  AO22X1 U95 ( .IN1(n72), .IN2(n106), .IN3(n74), .IN4(n107), .Q(n105) );
  AO221X1 U96 ( .IN1(HASH0[16]), .IN2(n76), .IN3(HASH0[24]), .IN4(n77), .IN5(
        n108), .Q(n107) );
  AO22X1 U97 ( .IN1(HASH0[8]), .IN2(n79), .IN3(HASH0[0]), .IN4(n80), .Q(n108)
         );
  NOR2X0 U98 ( .IN1(CrcHash[5]), .IN2(N7), .QN(n74) );
  AO221X1 U99 ( .IN1(HASH1[16]), .IN2(n76), .IN3(HASH1[24]), .IN4(n77), .IN5(
        n111), .Q(n106) );
  AO22X1 U100 ( .IN1(HASH1[8]), .IN2(n79), .IN3(HASH1[0]), .IN4(n80), .Q(n111)
         );
  NOR2X0 U101 ( .IN1(n112), .IN2(N7), .QN(n72) );
  AO221X1 U102 ( .IN1(HASH0[17]), .IN2(n76), .IN3(HASH0[25]), .IN4(n77), .IN5(
        n113), .Q(n104) );
  AO22X1 U103 ( .IN1(HASH0[9]), .IN2(n79), .IN3(HASH0[1]), .IN4(n80), .Q(n113)
         );
  NOR2X0 U104 ( .IN1(n114), .IN2(CrcHash[5]), .QN(n69) );
  AO221X1 U105 ( .IN1(HASH1[17]), .IN2(n76), .IN3(HASH1[25]), .IN4(n77), .IN5(
        n115), .Q(n103) );
  AO22X1 U106 ( .IN1(HASH1[9]), .IN2(n79), .IN3(HASH1[1]), .IN4(n80), .Q(n115)
         );
  NOR2X0 U107 ( .IN1(CrcHash[3]), .IN2(CrcHash[4]), .QN(n80) );
  NOR2X0 U108 ( .IN1(n116), .IN2(CrcHash[4]), .QN(n79) );
  NOR2X0 U109 ( .IN1(n117), .IN2(n116), .QN(n77) );
  INVX0 U110 ( .INP(CrcHash[3]), .ZN(n116) );
  NOR2X0 U111 ( .IN1(n117), .IN2(CrcHash[3]), .QN(n76) );
  INVX0 U112 ( .INP(CrcHash[4]), .ZN(n117) );
  NOR2X0 U113 ( .IN1(n114), .IN2(n112), .QN(n67) );
  INVX0 U114 ( .INP(CrcHash[5]), .ZN(n112) );
  INVX0 U115 ( .INP(N7), .ZN(n114) );
  INVX0 U116 ( .INP(RxEndFrm), .ZN(n59) );
  MUX21X1 U117 ( .IN1(n118), .IN2(AddressMiss), .S(n5), .Q(n102) );
  NOR4X0 U118 ( .IN1(n119), .IN2(n120), .IN3(n121), .IN4(n122), .QN(n118) );
  AND2X1 U119 ( .IN1(PassAll), .IN2(ControlFrmAddressOK), .Q(n121) );
  NOR4X0 U120 ( .IN1(n123), .IN2(n120), .IN3(r_Pro), .IN4(n122), .QN(N10) );
  NOR2X0 U121 ( .IN1(n124), .IN2(r_Bro), .QN(n122) );
  INVX0 U122 ( .INP(Broadcast), .ZN(n124) );
  OR2X1 U123 ( .IN1(n5), .IN2(n119), .Q(n123) );
  NAND2X0 U124 ( .IN1(ByteCntEq7), .IN2(n26), .QN(n5) );
  INVX0 U125 ( .INP(n58), .ZN(n26) );
  NOR2X0 U126 ( .IN1(StateData[0]), .IN2(StateData[1]), .QN(n58) );
endmodule


module eth_crc_test_1 ( Clk, Reset, Data, Enable, Initialize, Crc, CrcError, 
        eth_top_test_point_11887_in, test_si, test_se );
  input [3:0] Data;
  output [31:0] Crc;
  input Clk, Reset, Enable, Initialize, eth_top_test_point_11887_in, test_si,
         test_se;
  output CrcError;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N83, n97, n98, n99, n100, n101, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n126, n127, n66, n67, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57;
  assign CrcError = N83;

  SDFFASX1 \Crc_reg[0]  ( .D(N3), .SI(test_si), .SE(test_se), .CLK(Clk), 
        .SETB(n57), .Q(Crc[0]), .QN(n99) );
  SDFFASX1 \Crc_reg[4]  ( .D(N7), .SI(Crc[3]), .SE(test_se), .CLK(Clk), .SETB(
        n57), .Q(Crc[4]), .QN(n121) );
  SDFFASX1 \Crc_reg[8]  ( .D(N11), .SI(Crc[7]), .SE(test_se), .CLK(Clk), 
        .SETB(n57), .Q(Crc[8]), .QN(n117) );
  SDFFASX1 \Crc_reg[12]  ( .D(N15), .SI(Crc[11]), .SE(test_se), .CLK(Clk), 
        .SETB(n57), .Q(Crc[12]), .QN(n113) );
  SDFFASX1 \Crc_reg[16]  ( .D(N19), .SI(Crc[15]), .SE(test_se), .CLK(Clk), 
        .SETB(n57), .Q(Crc[16]), .QN(n127) );
  SDFFASX1 \Crc_reg[20]  ( .D(N23), .SI(Crc[19]), .SE(test_se), .CLK(Clk), 
        .SETB(n57), .Q(Crc[20]), .QN(n107) );
  SDFFASX1 \Crc_reg[24]  ( .D(N27), .SI(Crc[23]), .SE(test_se), .CLK(Clk), 
        .SETB(n57), .Q(Crc[24]), .QN(n103) );
  SDFFASX1 \Crc_reg[28]  ( .D(N31), .SI(Crc[27]), .SE(test_se), .CLK(Clk), 
        .SETB(n57), .Q(Crc[28]), .QN(n124) );
  SDFFASX1 \Crc_reg[22]  ( .D(N25), .SI(Crc[21]), .SE(test_se), .CLK(Clk), 
        .SETB(n57), .Q(Crc[22]), .QN(n105) );
  SDFFASX1 \Crc_reg[26]  ( .D(N29), .SI(Crc[25]), .SE(test_se), .CLK(Clk), 
        .SETB(n57), .Q(Crc[26]), .QN(n101) );
  SDFFASX1 \Crc_reg[30]  ( .D(N33), .SI(Crc[29]), .SE(test_se), .CLK(Clk), 
        .SETB(n57), .Q(Crc[30]), .QN(n66) );
  SDFFASX1 \Crc_reg[25]  ( .D(N28), .SI(Crc[24]), .SE(test_se), .CLK(Clk), 
        .SETB(n57), .Q(Crc[25]) );
  SDFFASX1 \Crc_reg[29]  ( .D(N32), .SI(Crc[28]), .SE(test_se), .CLK(Clk), 
        .SETB(n57), .Q(Crc[29]), .QN(n122) );
  SDFFASX1 \Crc_reg[1]  ( .D(N4), .SI(Crc[0]), .SE(test_se), .CLK(Clk), .SETB(
        n57), .Q(Crc[1]), .QN(n98) );
  SDFFASX1 \Crc_reg[2]  ( .D(N5), .SI(Crc[1]), .SE(test_se), .CLK(Clk), .SETB(
        n57), .Q(Crc[2]), .QN(n97) );
  SDFFASX1 \Crc_reg[6]  ( .D(N9), .SI(Crc[5]), .SE(test_se), .CLK(Clk), .SETB(
        n57), .Q(Crc[6]), .QN(n119) );
  SDFFASX1 \Crc_reg[10]  ( .D(N13), .SI(Crc[9]), .SE(test_se), .CLK(Clk), 
        .SETB(n57), .Q(Crc[10]), .QN(n115) );
  SDFFASX1 \Crc_reg[3]  ( .D(N6), .SI(Crc[2]), .SE(test_se), .CLK(Clk), .SETB(
        n57), .Q(Crc[3]), .QN(n123) );
  SDFFASX1 \Crc_reg[7]  ( .D(N10), .SI(Crc[6]), .SE(test_se), .CLK(Clk), 
        .SETB(n57), .Q(Crc[7]), .QN(n118) );
  SDFFASX1 \Crc_reg[27]  ( .D(N30), .SI(Crc[26]), .SE(test_se), .CLK(Clk), 
        .SETB(n57), .Q(Crc[27]), .QN(n100) );
  SDFFASX1 \Crc_reg[31]  ( .D(N34), .SI(Crc[30]), .SE(test_se), .CLK(Clk), 
        .SETB(n57), .Q(Crc[31]), .QN(n67) );
  SDFFASX1 \Crc_reg[5]  ( .D(N8), .SI(Crc[4]), .SE(test_se), .CLK(Clk), .SETB(
        n57), .Q(Crc[5]), .QN(n120) );
  SDFFASX1 \Crc_reg[9]  ( .D(N12), .SI(Crc[8]), .SE(test_se), .CLK(Clk), 
        .SETB(n57), .Q(Crc[9]), .QN(n116) );
  SDFFASX1 \Crc_reg[13]  ( .D(N16), .SI(Crc[12]), .SE(test_se), .CLK(Clk), 
        .SETB(n57), .Q(Crc[13]), .QN(n126) );
  SDFFASX1 \Crc_reg[11]  ( .D(N14), .SI(Crc[10]), .SE(test_se), .CLK(Clk), 
        .SETB(n57), .Q(Crc[11]), .QN(n114) );
  SDFFASX1 \Crc_reg[15]  ( .D(N18), .SI(Crc[14]), .SE(test_se), .CLK(Clk), 
        .SETB(n57), .Q(Crc[15]), .QN(n111) );
  SDFFASX1 \Crc_reg[19]  ( .D(N22), .SI(Crc[18]), .SE(test_se), .CLK(Clk), 
        .SETB(n57), .Q(Crc[19]), .QN(n108) );
  SDFFASX1 \Crc_reg[23]  ( .D(N26), .SI(Crc[22]), .SE(test_se), .CLK(Clk), 
        .SETB(n57), .Q(Crc[23]), .QN(n104) );
  SDFFASX1 \Crc_reg[17]  ( .D(N20), .SI(Crc[16]), .SE(test_se), .CLK(Clk), 
        .SETB(n57), .Q(Crc[17]), .QN(n110) );
  SDFFASX1 \Crc_reg[21]  ( .D(N24), .SI(Crc[20]), .SE(test_se), .CLK(Clk), 
        .SETB(n57), .Q(Crc[21]), .QN(n106) );
  SDFFASX1 \Crc_reg[14]  ( .D(N17), .SI(Crc[13]), .SE(test_se), .CLK(Clk), 
        .SETB(n57), .Q(Crc[14]), .QN(n112) );
  SDFFASX1 \Crc_reg[18]  ( .D(N21), .SI(Crc[17]), .SE(test_se), .CLK(Clk), 
        .SETB(n57), .Q(Crc[18]), .QN(n109) );
  INVX0 U3 ( .INP(eth_top_test_point_11887_in), .ZN(n57) );
  NAND2X0 U4 ( .IN1(n1), .IN2(n2), .QN(N9) );
  XNOR2X1 U5 ( .IN1(n97), .IN2(n3), .Q(n1) );
  NAND2X0 U6 ( .IN1(n4), .IN2(n5), .QN(N83) );
  NOR4X0 U7 ( .IN1(n6), .IN2(n7), .IN3(n8), .IN4(n9), .QN(n5) );
  OR4X1 U8 ( .IN1(n103), .IN2(n109), .IN3(n111), .IN4(n112), .Q(n9) );
  OR4X1 U9 ( .IN1(n113), .IN2(n114), .IN3(n115), .IN4(n117), .Q(n8) );
  OR4X1 U10 ( .IN1(n119), .IN2(n120), .IN3(n121), .IN4(n123), .Q(n7) );
  OR4X1 U11 ( .IN1(n66), .IN2(n67), .IN3(n98), .IN4(n99), .Q(n6) );
  NOR4X0 U12 ( .IN1(n10), .IN2(n11), .IN3(n12), .IN4(n13), .QN(n4) );
  NAND4X0 U13 ( .IN1(n127), .IN2(n126), .IN3(n124), .IN4(n118), .QN(n13) );
  NAND4X0 U14 ( .IN1(n116), .IN2(n110), .IN3(n108), .IN4(n107), .QN(n12) );
  NAND4X0 U15 ( .IN1(n106), .IN2(n105), .IN3(n104), .IN4(n100), .QN(n11) );
  NAND4X0 U16 ( .IN1(n97), .IN2(n122), .IN3(Crc[26]), .IN4(Crc[25]), .QN(n10)
         );
  NAND2X0 U17 ( .IN1(n14), .IN2(n2), .QN(N8) );
  XNOR2X1 U18 ( .IN1(n98), .IN2(n15), .Q(n14) );
  NAND2X0 U19 ( .IN1(n16), .IN2(n2), .QN(N7) );
  XNOR2X1 U20 ( .IN1(n99), .IN2(n17), .Q(n16) );
  NAND2X0 U21 ( .IN1(n18), .IN2(n2), .QN(N6) );
  NAND2X0 U22 ( .IN1(n19), .IN2(n2), .QN(N5) );
  OR2X1 U23 ( .IN1(Initialize), .IN2(n20), .Q(N4) );
  NAND2X0 U24 ( .IN1(n100), .IN2(n2), .QN(N34) );
  NAND2X0 U25 ( .IN1(n101), .IN2(n2), .QN(N33) );
  NAND2X0 U26 ( .IN1(n21), .IN2(n2), .QN(N32) );
  XNOR2X1 U27 ( .IN1(Crc[25]), .IN2(n22), .Q(n21) );
  NAND2X0 U28 ( .IN1(n23), .IN2(n2), .QN(N31) );
  XOR2X1 U29 ( .IN1(n103), .IN2(n24), .Q(n23) );
  NAND2X0 U30 ( .IN1(n25), .IN2(n2), .QN(N30) );
  XOR2X1 U31 ( .IN1(n104), .IN2(n26), .Q(n25) );
  OR2X1 U32 ( .IN1(Initialize), .IN2(n27), .Q(N3) );
  NAND2X0 U33 ( .IN1(n28), .IN2(n2), .QN(N29) );
  XNOR2X1 U34 ( .IN1(n105), .IN2(n29), .Q(n28) );
  NAND2X0 U35 ( .IN1(Enable), .IN2(n30), .QN(n29) );
  XOR2X1 U36 ( .IN1(n31), .IN2(n32), .Q(n30) );
  NAND2X0 U37 ( .IN1(n33), .IN2(n2), .QN(N28) );
  XOR2X1 U38 ( .IN1(n106), .IN2(n34), .Q(n33) );
  NAND2X0 U39 ( .IN1(n35), .IN2(n2), .QN(N27) );
  XNOR2X1 U40 ( .IN1(n107), .IN2(n3), .Q(n35) );
  NAND2X0 U41 ( .IN1(n36), .IN2(n2), .QN(N26) );
  XOR2X1 U42 ( .IN1(n108), .IN2(n20), .Q(n36) );
  NAND2X0 U43 ( .IN1(n37), .IN2(n2), .QN(N25) );
  XOR2X1 U44 ( .IN1(n109), .IN2(n27), .Q(n37) );
  NAND2X0 U45 ( .IN1(n110), .IN2(n2), .QN(N24) );
  NAND2X0 U46 ( .IN1(n127), .IN2(n2), .QN(N23) );
  NAND2X0 U47 ( .IN1(n38), .IN2(n2), .QN(N22) );
  XOR2X1 U48 ( .IN1(n111), .IN2(n22), .Q(n38) );
  NAND2X0 U49 ( .IN1(n39), .IN2(n2), .QN(N21) );
  XOR2X1 U50 ( .IN1(n112), .IN2(n24), .Q(n39) );
  NAND2X0 U51 ( .IN1(n40), .IN2(n2), .QN(N20) );
  XOR2X1 U52 ( .IN1(n126), .IN2(n26), .Q(n40) );
  NAND2X0 U53 ( .IN1(n41), .IN2(n2), .QN(N19) );
  XOR2X1 U54 ( .IN1(n113), .IN2(n27), .Q(n41) );
  NAND2X0 U55 ( .IN1(n42), .IN2(n2), .QN(N18) );
  XOR2X1 U56 ( .IN1(n114), .IN2(n22), .Q(n42) );
  NAND2X0 U57 ( .IN1(n43), .IN2(n2), .QN(N17) );
  XOR2X1 U58 ( .IN1(n115), .IN2(n34), .Q(n43) );
  NAND2X0 U59 ( .IN1(n44), .IN2(n2), .QN(N16) );
  XNOR2X1 U60 ( .IN1(n116), .IN2(n18), .Q(n44) );
  AOI22X1 U61 ( .IN1(n34), .IN2(n45), .IN3(n26), .IN4(n46), .QN(n18) );
  NOR2X0 U62 ( .IN1(n47), .IN2(n45), .QN(n26) );
  NAND2X0 U63 ( .IN1(n48), .IN2(n2), .QN(N15) );
  XNOR2X1 U64 ( .IN1(n117), .IN2(n19), .Q(n48) );
  AOI22X1 U65 ( .IN1(n24), .IN2(n49), .IN3(n20), .IN4(n50), .QN(n19) );
  NOR2X0 U66 ( .IN1(n47), .IN2(n50), .QN(n24) );
  NAND2X0 U67 ( .IN1(n51), .IN2(n2), .QN(N14) );
  XNOR2X1 U68 ( .IN1(n118), .IN2(n15), .Q(n51) );
  NAND2X0 U69 ( .IN1(n52), .IN2(n2), .QN(N13) );
  XNOR2X1 U70 ( .IN1(n119), .IN2(n17), .Q(n52) );
  NAND2X0 U71 ( .IN1(n53), .IN2(n2), .QN(N12) );
  XNOR2X1 U72 ( .IN1(n120), .IN2(n3), .Q(n53) );
  NAND2X0 U73 ( .IN1(Enable), .IN2(n54), .QN(n3) );
  XOR2X1 U74 ( .IN1(n45), .IN2(n50), .Q(n54) );
  NAND2X0 U75 ( .IN1(n55), .IN2(n2), .QN(N11) );
  XNOR2X1 U76 ( .IN1(n121), .IN2(n15), .Q(n55) );
  AOI22X1 U77 ( .IN1(n22), .IN2(n49), .IN3(n20), .IN4(n31), .QN(n15) );
  NOR2X0 U78 ( .IN1(n47), .IN2(n49), .QN(n20) );
  XNOR2X1 U79 ( .IN1(n32), .IN2(n45), .Q(n49) );
  XOR2X1 U80 ( .IN1(n122), .IN2(Data[1]), .Q(n45) );
  NOR2X0 U81 ( .IN1(n31), .IN2(n47), .QN(n22) );
  NAND2X0 U82 ( .IN1(n56), .IN2(n2), .QN(N10) );
  INVX0 U83 ( .INP(Initialize), .ZN(n2) );
  XNOR2X1 U84 ( .IN1(n123), .IN2(n17), .Q(n56) );
  AOI22X1 U85 ( .IN1(n34), .IN2(n32), .IN3(n27), .IN4(n46), .QN(n17) );
  NOR2X0 U86 ( .IN1(n32), .IN2(n47), .QN(n27) );
  XOR2X1 U87 ( .IN1(n124), .IN2(Data[0]), .Q(n32) );
  NOR2X0 U88 ( .IN1(n47), .IN2(n46), .QN(n34) );
  XNOR2X1 U89 ( .IN1(n31), .IN2(n50), .Q(n46) );
  XOR2X1 U90 ( .IN1(n66), .IN2(Data[2]), .Q(n50) );
  XOR2X1 U91 ( .IN1(n67), .IN2(Data[3]), .Q(n31) );
  INVX0 U92 ( .INP(Enable), .ZN(n47) );
endmodule


module eth_rxethmac_test_1 ( MRxClk, MRxDV, MRxD, Reset, Transmitting, MaxFL, 
        r_IFG, HugEn, DlyCrcEn, RxData, RxValid, RxStartFrm, RxEndFrm, ByteCnt, 
        ByteCntEq0, ByteCntGreat2, ByteCntMaxFrame, CrcError, StateIdle, 
        StatePreamble, StateSFD, StateData, MAC, r_Pro, r_Bro, r_HASH0, 
        r_HASH1, RxAbort, AddressMiss, PassAll, ControlFrmAddressOK, 
        eth_top_test_point_11887_in, test_si, test_se );
  input [3:0] MRxD;
  input [15:0] MaxFL;
  output [7:0] RxData;
  output [15:0] ByteCnt;
  output [1:0] StateData;
  input [47:0] MAC;
  input [31:0] r_HASH0;
  input [31:0] r_HASH1;
  input MRxClk, MRxDV, Reset, Transmitting, r_IFG, HugEn, DlyCrcEn, r_Pro,
         r_Bro, PassAll, ControlFrmAddressOK, eth_top_test_point_11887_in,
         test_si, test_se;
  output RxValid, RxStartFrm, RxEndFrm, ByteCntEq0, ByteCntGreat2,
         ByteCntMaxFrame, CrcError, StateIdle, StatePreamble, StateSFD,
         RxAbort, AddressMiss;
  wire   IFGCounterEq24, StateDrop, ByteCntEq1, ByteCntEq2, ByteCntEq3,
         ByteCntEq4, ByteCntEq5, ByteCntEq6, ByteCntEq7, ByteCntSmall7,
         Broadcast, CrcHashGood, Multicast, Enable_Crc, Initialize_Crc,
         DelayData, RxValid_d, GenerateRxStartFrm, RxStartFrm_d,
         GenerateRxEndFrm, N51, n55, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n1, n2, n3, n4,
         n76, n77, n78, n79, n80, n81, n82, n101, n105, n106, n107, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37;
  wire   [3:0] DlyCrcCnt;
  wire   [5:0] CrcHash;
  wire   [31:0] Crc;
  wire   [7:0] LatchedByte;
  wire   [7:0] RxData_d;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25;

  SDFFX1 CrcHashGood_reg ( .D(n37), .SI(Broadcast), .SE(test_se), .CLK(MRxClk), 
        .Q(CrcHashGood) );
  SDFFX1 \CrcHash_reg[5]  ( .D(n98), .SI(CrcHash[4]), .SE(test_se), .CLK(
        MRxClk), .Q(CrcHash[5]) );
  SDFFX1 \CrcHash_reg[4]  ( .D(n97), .SI(CrcHash[3]), .SE(test_se), .CLK(
        MRxClk), .Q(CrcHash[4]) );
  SDFFX1 \CrcHash_reg[3]  ( .D(n96), .SI(CrcHash[2]), .SE(test_se), .CLK(
        MRxClk), .Q(CrcHash[3]) );
  SDFFX1 \CrcHash_reg[2]  ( .D(n95), .SI(CrcHash[1]), .SE(test_se), .CLK(
        MRxClk), .Q(CrcHash[2]) );
  SDFFX1 \CrcHash_reg[1]  ( .D(n94), .SI(CrcHash[0]), .SE(test_se), .CLK(
        MRxClk), .Q(CrcHash[1]) );
  SDFFX1 \CrcHash_reg[0]  ( .D(n93), .SI(CrcHashGood), .SE(test_se), .CLK(
        MRxClk), .Q(CrcHash[0]) );
  SDFFARX1 \LatchedByte_reg[7]  ( .D(MRxD[3]), .SI(LatchedByte[6]), .SE(
        test_se), .CLK(MRxClk), .RSTB(n5), .Q(LatchedByte[7]), .QN(n77) );
  SDFFARX1 \LatchedByte_reg[6]  ( .D(MRxD[2]), .SI(LatchedByte[5]), .SE(
        test_se), .CLK(MRxClk), .RSTB(n6), .Q(LatchedByte[6]), .QN(n78) );
  SDFFARX1 \LatchedByte_reg[5]  ( .D(MRxD[1]), .SI(LatchedByte[4]), .SE(
        test_se), .CLK(MRxClk), .RSTB(n5), .Q(LatchedByte[5]), .QN(n79) );
  SDFFARX1 \LatchedByte_reg[4]  ( .D(MRxD[0]), .SI(n4), .SE(test_se), .CLK(
        MRxClk), .RSTB(n6), .Q(LatchedByte[4]), .QN(n80) );
  SDFFARX1 \LatchedByte_reg[3]  ( .D(LatchedByte[7]), .SI(n3), .SE(test_se), 
        .CLK(MRxClk), .RSTB(n5), .Q(n4), .QN(n81) );
  SDFFARX1 \LatchedByte_reg[2]  ( .D(LatchedByte[6]), .SI(n2), .SE(test_se), 
        .CLK(MRxClk), .RSTB(n6), .Q(n3), .QN(n82) );
  SDFFARX1 \LatchedByte_reg[1]  ( .D(LatchedByte[5]), .SI(n1), .SE(test_se), 
        .CLK(MRxClk), .RSTB(n5), .Q(n2) );
  SDFFARX1 \LatchedByte_reg[0]  ( .D(LatchedByte[4]), .SI(DelayData), .SE(
        test_se), .CLK(MRxClk), .RSTB(n6), .Q(n1) );
  SDFFARX1 DelayData_reg ( .D(StateData[0]), .SI(CrcHash[5]), .SE(test_se), 
        .CLK(MRxClk), .RSTB(n5), .Q(DelayData) );
  SDFFARX1 \RxData_d_reg[7]  ( .D(n85), .SI(RxData_d[6]), .SE(test_se), .CLK(
        MRxClk), .RSTB(n5), .Q(RxData_d[7]) );
  SDFFARX1 \RxData_reg[7]  ( .D(RxData_d[7]), .SI(RxData[6]), .SE(test_se), 
        .CLK(MRxClk), .RSTB(n6), .Q(RxData[7]) );
  SDFFARX1 \RxData_d_reg[6]  ( .D(n86), .SI(RxData_d[5]), .SE(test_se), .CLK(
        MRxClk), .RSTB(n6), .Q(RxData_d[6]) );
  SDFFARX1 \RxData_reg[6]  ( .D(RxData_d[6]), .SI(RxData[5]), .SE(test_se), 
        .CLK(MRxClk), .RSTB(n5), .Q(RxData[6]) );
  SDFFARX1 \RxData_d_reg[5]  ( .D(n87), .SI(RxData_d[4]), .SE(test_se), .CLK(
        MRxClk), .RSTB(n5), .Q(RxData_d[5]) );
  SDFFARX1 \RxData_reg[5]  ( .D(RxData_d[5]), .SI(RxData[4]), .SE(test_se), 
        .CLK(MRxClk), .RSTB(n6), .Q(RxData[5]) );
  SDFFARX1 \RxData_d_reg[4]  ( .D(n88), .SI(RxData_d[3]), .SE(test_se), .CLK(
        MRxClk), .RSTB(n6), .Q(RxData_d[4]) );
  SDFFARX1 \RxData_reg[4]  ( .D(RxData_d[4]), .SI(RxData[3]), .SE(test_se), 
        .CLK(MRxClk), .RSTB(n5), .Q(RxData[4]) );
  SDFFARX1 \RxData_d_reg[3]  ( .D(n89), .SI(RxData_d[2]), .SE(test_se), .CLK(
        MRxClk), .RSTB(n5), .Q(RxData_d[3]) );
  SDFFARX1 \RxData_reg[3]  ( .D(RxData_d[3]), .SI(RxData[2]), .SE(test_se), 
        .CLK(MRxClk), .RSTB(n6), .Q(RxData[3]) );
  SDFFARX1 \RxData_d_reg[2]  ( .D(n90), .SI(RxData_d[1]), .SE(test_se), .CLK(
        MRxClk), .RSTB(n6), .Q(RxData_d[2]) );
  SDFFARX1 \RxData_reg[2]  ( .D(RxData_d[2]), .SI(RxData[1]), .SE(test_se), 
        .CLK(MRxClk), .RSTB(n5), .Q(RxData[2]) );
  SDFFARX1 \RxData_d_reg[1]  ( .D(n91), .SI(RxData_d[0]), .SE(test_se), .CLK(
        MRxClk), .RSTB(n5), .Q(RxData_d[1]) );
  SDFFARX1 \RxData_reg[1]  ( .D(RxData_d[1]), .SI(RxData[0]), .SE(test_se), 
        .CLK(MRxClk), .RSTB(n6), .Q(RxData[1]) );
  SDFFARX1 \RxData_d_reg[0]  ( .D(n92), .SI(Multicast), .SE(test_se), .CLK(
        MRxClk), .RSTB(n6), .Q(RxData_d[0]) );
  SDFFARX1 \RxData_reg[0]  ( .D(RxData_d[0]), .SI(RxData_d[7]), .SE(test_se), 
        .CLK(MRxClk), .RSTB(n5), .Q(RxData[0]) );
  SDFFARX1 RxValid_d_reg ( .D(n36), .SI(RxStartFrm), .SE(test_se), .CLK(MRxClk), .RSTB(n5), .Q(RxValid_d) );
  SDFFARX1 RxValid_reg ( .D(RxValid_d), .SI(RxValid_d), .SE(test_se), .CLK(
        MRxClk), .RSTB(n6), .Q(RxValid) );
  SDFFARX1 RxStartFrm_d_reg ( .D(GenerateRxStartFrm), .SI(RxEndFrm), .SE(
        test_se), .CLK(MRxClk), .RSTB(n6), .Q(RxStartFrm_d) );
  SDFFARX1 RxStartFrm_reg ( .D(RxStartFrm_d), .SI(RxStartFrm_d), .SE(test_se), 
        .CLK(MRxClk), .RSTB(n5), .Q(RxStartFrm) );
  SDFFARX1 RxEndFrm_d_reg ( .D(GenerateRxEndFrm), .SI(RxData[7]), .SE(test_se), 
        .CLK(MRxClk), .RSTB(n5), .Q(n107), .QN(n101) );
  SDFFARX1 RxEndFrm_reg ( .D(N51), .SI(n107), .SE(test_se), .CLK(MRxClk), 
        .RSTB(n6), .Q(RxEndFrm), .QN(n55) );
  SDFFARX1 Multicast_reg ( .D(n83), .SI(LatchedByte[7]), .SE(test_se), .CLK(
        MRxClk), .RSTB(n5), .Q(Multicast), .QN(n76) );
  SDFFARX1 Broadcast_reg ( .D(n84), .SI(test_si), .SE(test_se), .CLK(MRxClk), 
        .RSTB(n6), .Q(Broadcast) );
  eth_rxstatem_test_1 rxstatem1 ( .MRxClk(MRxClk), .Reset(Reset), .MRxDV(MRxDV), .ByteCntEq0(ByteCntEq0), .ByteCntGreat2(ByteCntGreat2), .Transmitting(
        Transmitting), .MRxDEq5(n99), .MRxDEqD(n100), .IFGCounterEq24(
        IFGCounterEq24), .ByteCntMaxFrame(ByteCntMaxFrame), .StateData(
        StateData), .StateIdle(StateIdle), .StatePreamble(StatePreamble), 
        .StateSFD(StateSFD), .StateDrop(StateDrop), 
        .eth_top_test_point_11887_in(eth_top_test_point_11887_in), .test_si(
        n105), .test_se(test_se) );
  eth_rxcounters_test_1 rxcounters1 ( .MRxClk(MRxClk), .Reset(Reset), .MRxDV(
        MRxDV), .StateIdle(StateIdle), .StateSFD(StateSFD), .StateData(
        StateData), .StateDrop(StateDrop), .StatePreamble(StatePreamble), 
        .MRxDEqD(n100), .DlyCrcEn(DlyCrcEn), .DlyCrcCnt(DlyCrcCnt), 
        .Transmitting(Transmitting), .MaxFL(MaxFL), .r_IFG(r_IFG), .HugEn(
        HugEn), .IFGCounterEq24(IFGCounterEq24), .ByteCntEq0(ByteCntEq0), 
        .ByteCntEq1(ByteCntEq1), .ByteCntEq2(ByteCntEq2), .ByteCntEq3(
        ByteCntEq3), .ByteCntEq4(ByteCntEq4), .ByteCntEq5(ByteCntEq5), 
        .ByteCntEq6(ByteCntEq6), .ByteCntEq7(ByteCntEq7), .ByteCntGreat2(
        ByteCntGreat2), .ByteCntSmall7(ByteCntSmall7), .ByteCntMaxFrame(
        ByteCntMaxFrame), .ByteCntOut(ByteCnt), .eth_top_test_point_11887_in(
        eth_top_test_point_11887_in), .test_si(n106), .test_so(n105), 
        .test_se(test_se) );
  eth_rxaddrcheck_test_1 rxaddrcheck1 ( .MRxClk(MRxClk), .Reset(Reset), 
        .RxData(RxData), .Broadcast(Broadcast), .r_Bro(r_Bro), .r_Pro(r_Pro), 
        .ByteCntEq2(ByteCntEq2), .ByteCntEq3(ByteCntEq3), .ByteCntEq4(
        ByteCntEq4), .ByteCntEq5(ByteCntEq5), .ByteCntEq6(ByteCntEq6), 
        .ByteCntEq7(ByteCntEq7), .HASH0(r_HASH0), .HASH1(r_HASH1), .CrcHash(
        CrcHash), .CrcHashGood(CrcHashGood), .StateData(StateData), .RxEndFrm(
        RxEndFrm), .Multicast(Multicast), .MAC(MAC), .RxAbort(RxAbort), 
        .AddressMiss(AddressMiss), .PassAll(PassAll), .ControlFrmAddressOK(
        ControlFrmAddressOK), .eth_top_test_point_11887_in(
        eth_top_test_point_11887_in), .test_si(Crc[31]), .test_so(n106), 
        .test_se(test_se) );
  eth_crc_test_1 crcrx ( .Clk(MRxClk), .Reset(Reset), .Data({MRxD[0], MRxD[1], 
        MRxD[2], MRxD[3]}), .Enable(Enable_Crc), .Initialize(Initialize_Crc), 
        .Crc({Crc[31:26], SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25}), .CrcError(
        CrcError), .eth_top_test_point_11887_in(eth_top_test_point_11887_in), 
        .test_si(RxValid), .test_se(test_se) );
  INVX0 U3 ( .INP(eth_top_test_point_11887_in), .ZN(n5) );
  INVX0 U4 ( .INP(eth_top_test_point_11887_in), .ZN(n6) );
  INVX0 U5 ( .INP(n7), .ZN(n37) );
  NOR2X0 U6 ( .IN1(MRxD[3]), .IN2(n8), .QN(n99) );
  AO22X1 U7 ( .IN1(Crc[31]), .IN2(n9), .IN3(n10), .IN4(CrcHash[5]), .Q(n98) );
  AO22X1 U8 ( .IN1(Crc[30]), .IN2(n9), .IN3(n10), .IN4(CrcHash[4]), .Q(n97) );
  AO22X1 U9 ( .IN1(Crc[29]), .IN2(n9), .IN3(n10), .IN4(CrcHash[3]), .Q(n96) );
  AO22X1 U10 ( .IN1(Crc[28]), .IN2(n9), .IN3(n10), .IN4(CrcHash[2]), .Q(n95)
         );
  AO22X1 U11 ( .IN1(Crc[27]), .IN2(n9), .IN3(n10), .IN4(CrcHash[1]), .Q(n94)
         );
  AO22X1 U12 ( .IN1(Crc[26]), .IN2(n9), .IN3(n10), .IN4(CrcHash[0]), .Q(n93)
         );
  NOR3X0 U13 ( .IN1(Reset), .IN2(StateIdle), .IN3(n9), .QN(n10) );
  NOR3X0 U14 ( .IN1(Reset), .IN2(StateIdle), .IN3(n7), .QN(n9) );
  NAND2X0 U15 ( .IN1(ByteCntEq6), .IN2(StateData[0]), .QN(n7) );
  AO22X1 U16 ( .IN1(n36), .IN2(n1), .IN3(n11), .IN4(RxData_d[0]), .Q(n92) );
  AO22X1 U17 ( .IN1(n36), .IN2(n2), .IN3(n11), .IN4(RxData_d[1]), .Q(n91) );
  AO22X1 U18 ( .IN1(n36), .IN2(n3), .IN3(n11), .IN4(RxData_d[2]), .Q(n90) );
  AO22X1 U19 ( .IN1(n36), .IN2(n4), .IN3(n11), .IN4(RxData_d[3]), .Q(n89) );
  AO22X1 U20 ( .IN1(n36), .IN2(LatchedByte[4]), .IN3(n11), .IN4(RxData_d[4]), 
        .Q(n88) );
  AO22X1 U21 ( .IN1(n36), .IN2(LatchedByte[5]), .IN3(n11), .IN4(RxData_d[5]), 
        .Q(n87) );
  AO22X1 U22 ( .IN1(n36), .IN2(LatchedByte[6]), .IN3(n11), .IN4(RxData_d[6]), 
        .Q(n86) );
  AO22X1 U23 ( .IN1(n36), .IN2(LatchedByte[7]), .IN3(n11), .IN4(RxData_d[7]), 
        .Q(n85) );
  AND2X1 U24 ( .IN1(n12), .IN2(DelayData), .Q(n11) );
  INVX0 U25 ( .INP(n12), .ZN(n36) );
  NAND2X0 U26 ( .IN1(StateData[0]), .IN2(n13), .QN(n12) );
  NAND4X0 U27 ( .IN1(ByteCntEq0), .IN2(n14), .IN3(n15), .IN4(n16), .QN(n13) );
  INVX0 U28 ( .INP(DlyCrcCnt[2]), .ZN(n15) );
  OAI21X1 U29 ( .IN1(n17), .IN2(n18), .IN3(n19), .QN(n84) );
  NAND4X0 U30 ( .IN1(n55), .IN2(n20), .IN3(n21), .IN4(Broadcast), .QN(n19) );
  INVX0 U31 ( .INP(RxAbort), .ZN(n21) );
  NAND3X0 U32 ( .IN1(StateData[0]), .IN2(n17), .IN3(ByteCntSmall7), .QN(n20)
         );
  NAND4X0 U33 ( .IN1(n2), .IN2(n1), .IN3(n22), .IN4(n23), .QN(n17) );
  NOR4X0 U34 ( .IN1(n82), .IN2(n81), .IN3(n80), .IN4(n79), .QN(n23) );
  NOR2X0 U35 ( .IN1(n78), .IN2(n77), .QN(n22) );
  AO22X1 U36 ( .IN1(n24), .IN2(n1), .IN3(n25), .IN4(n55), .Q(n83) );
  NOR2X0 U37 ( .IN1(n76), .IN2(RxAbort), .QN(n25) );
  NOR2X0 U38 ( .IN1(n8), .IN2(n26), .QN(n100) );
  INVX0 U39 ( .INP(MRxD[3]), .ZN(n26) );
  NAND3X0 U40 ( .IN1(MRxD[0]), .IN2(n27), .IN3(MRxD[2]), .QN(n8) );
  INVX0 U41 ( .INP(MRxD[1]), .ZN(n27) );
  NAND2X0 U42 ( .IN1(n101), .IN2(n28), .QN(N51) );
  NAND3X0 U43 ( .IN1(ByteCntGreat2), .IN2(n29), .IN3(StateData[1]), .QN(n28)
         );
  AO21X1 U44 ( .IN1(n30), .IN2(DlyCrcEn), .IN3(StateSFD), .Q(Initialize_Crc)
         );
  XNOR2X1 U45 ( .IN1(n31), .IN2(n16), .Q(n30) );
  INVX0 U46 ( .INP(DlyCrcCnt[3]), .ZN(n16) );
  OR3X1 U47 ( .IN1(DlyCrcCnt[1]), .IN2(DlyCrcCnt[2]), .IN3(DlyCrcCnt[0]), .Q(
        n31) );
  MUX21X1 U48 ( .IN1(n24), .IN2(n32), .S(DlyCrcEn), .Q(GenerateRxStartFrm) );
  NOR4X0 U49 ( .IN1(DlyCrcCnt[3]), .IN2(DlyCrcCnt[2]), .IN3(n33), .IN4(n14), 
        .QN(n32) );
  NAND2X0 U50 ( .IN1(DlyCrcCnt[1]), .IN2(DlyCrcCnt[0]), .QN(n14) );
  INVX0 U51 ( .INP(n18), .ZN(n24) );
  NAND2X0 U52 ( .IN1(ByteCntEq1), .IN2(StateData[0]), .QN(n18) );
  NOR2X0 U53 ( .IN1(n34), .IN2(n33), .QN(GenerateRxEndFrm) );
  INVX0 U54 ( .INP(StateData[0]), .ZN(n33) );
  AOI21X1 U55 ( .IN1(n29), .IN2(ByteCntGreat2), .IN3(ByteCntMaxFrame), .QN(n34) );
  NOR3X0 U56 ( .IN1(n29), .IN2(ByteCntMaxFrame), .IN3(n35), .QN(Enable_Crc) );
  NOR2X0 U57 ( .IN1(StateData[0]), .IN2(StateData[1]), .QN(n35) );
  INVX0 U58 ( .INP(MRxDV), .ZN(n29) );
endmodule


module eth_spram_256x32_test_1 ( clk, rst, ce, we, oe, addr, di, do, test_si8, 
        test_si7, test_si6, test_si5, test_si4, test_si3, test_si2, test_si1, 
        test_so8, test_so7, test_so6, test_so5, test_so4, test_so3, test_so2, 
        test_so1, test_se );
  input [3:0] we;
  input [7:0] addr;
  input [31:0] di;
  output [31:0] do;
  input clk, rst, ce, oe, test_si8, test_si7, test_si6, test_si5, test_si4,
         test_si3, test_si2, test_si1, test_se;
  output test_so8, test_so7, test_so6, test_so5, test_so4, test_so3, test_so2,
         test_so1;
  wire   N54, N55, N56, N57, N58, N59, N60, N61, \mem3[255][31] ,
         \mem3[255][30] , \mem3[255][29] , \mem3[255][28] , \mem3[255][27] ,
         \mem3[255][26] , \mem3[255][25] , \mem3[255][24] , \mem3[254][31] ,
         \mem3[254][30] , \mem3[254][29] , \mem3[254][28] , \mem3[254][27] ,
         \mem3[254][26] , \mem3[254][25] , \mem3[254][24] , \mem3[253][31] ,
         \mem3[253][30] , \mem3[253][29] , \mem3[253][28] , \mem3[253][27] ,
         \mem3[253][26] , \mem3[253][25] , \mem3[253][24] , \mem3[252][31] ,
         \mem3[252][30] , \mem3[252][29] , \mem3[252][28] , \mem3[252][27] ,
         \mem3[252][26] , \mem3[252][25] , \mem3[252][24] , \mem3[251][31] ,
         \mem3[251][30] , \mem3[251][29] , \mem3[251][28] , \mem3[251][27] ,
         \mem3[251][26] , \mem3[251][25] , \mem3[251][24] , \mem3[250][31] ,
         \mem3[250][30] , \mem3[250][29] , \mem3[250][28] , \mem3[250][27] ,
         \mem3[250][26] , \mem3[250][25] , \mem3[250][24] , \mem3[249][31] ,
         \mem3[249][30] , \mem3[249][29] , \mem3[249][28] , \mem3[249][27] ,
         \mem3[249][26] , \mem3[249][25] , \mem3[249][24] , \mem3[248][31] ,
         \mem3[248][30] , \mem3[248][29] , \mem3[248][28] , \mem3[248][27] ,
         \mem3[248][26] , \mem3[248][25] , \mem3[248][24] , \mem3[247][31] ,
         \mem3[247][30] , \mem3[247][29] , \mem3[247][28] , \mem3[247][27] ,
         \mem3[247][26] , \mem3[247][25] , \mem3[247][24] , \mem3[246][31] ,
         \mem3[246][30] , \mem3[246][29] , \mem3[246][28] , \mem3[246][27] ,
         \mem3[246][26] , \mem3[246][25] , \mem3[246][24] , \mem3[245][31] ,
         \mem3[245][30] , \mem3[245][29] , \mem3[245][28] , \mem3[245][27] ,
         \mem3[245][26] , \mem3[245][25] , \mem3[245][24] , \mem3[244][31] ,
         \mem3[244][30] , \mem3[244][29] , \mem3[244][28] , \mem3[244][27] ,
         \mem3[244][26] , \mem3[244][25] , \mem3[244][24] , \mem3[243][31] ,
         \mem3[243][30] , \mem3[243][29] , \mem3[243][28] , \mem3[243][27] ,
         \mem3[243][26] , \mem3[243][25] , \mem3[243][24] , \mem3[242][31] ,
         \mem3[242][30] , \mem3[242][29] , \mem3[242][28] , \mem3[242][27] ,
         \mem3[242][26] , \mem3[242][25] , \mem3[242][24] , \mem3[241][31] ,
         \mem3[241][30] , \mem3[241][29] , \mem3[241][28] , \mem3[241][27] ,
         \mem3[241][26] , \mem3[241][25] , \mem3[241][24] , \mem3[240][31] ,
         \mem3[240][30] , \mem3[240][29] , \mem3[240][28] , \mem3[240][27] ,
         \mem3[240][26] , \mem3[240][25] , \mem3[240][24] , \mem3[239][31] ,
         \mem3[239][30] , \mem3[239][29] , \mem3[239][28] , \mem3[239][27] ,
         \mem3[239][26] , \mem3[239][25] , \mem3[239][24] , \mem3[238][31] ,
         \mem3[238][30] , \mem3[238][29] , \mem3[238][28] , \mem3[238][27] ,
         \mem3[238][26] , \mem3[238][25] , \mem3[238][24] , \mem3[237][31] ,
         \mem3[237][30] , \mem3[237][29] , \mem3[237][28] , \mem3[237][27] ,
         \mem3[237][26] , \mem3[237][25] , \mem3[237][24] , \mem3[236][31] ,
         \mem3[236][30] , \mem3[236][29] , \mem3[236][28] , \mem3[236][27] ,
         \mem3[236][26] , \mem3[236][25] , \mem3[236][24] , \mem3[235][31] ,
         \mem3[235][30] , \mem3[235][29] , \mem3[235][28] , \mem3[235][27] ,
         \mem3[235][26] , \mem3[235][25] , \mem3[235][24] , \mem3[234][31] ,
         \mem3[234][30] , \mem3[234][29] , \mem3[234][28] , \mem3[234][27] ,
         \mem3[234][26] , \mem3[234][25] , \mem3[234][24] , \mem3[233][31] ,
         \mem3[233][30] , \mem3[233][29] , \mem3[233][28] , \mem3[233][27] ,
         \mem3[233][26] , \mem3[233][25] , \mem3[233][24] , \mem3[232][31] ,
         \mem3[232][30] , \mem3[232][29] , \mem3[232][28] , \mem3[232][27] ,
         \mem3[232][26] , \mem3[232][25] , \mem3[232][24] , \mem3[231][31] ,
         \mem3[231][30] , \mem3[231][29] , \mem3[231][28] , \mem3[231][27] ,
         \mem3[231][26] , \mem3[231][25] , \mem3[231][24] , \mem3[230][31] ,
         \mem3[230][30] , \mem3[230][29] , \mem3[230][28] , \mem3[230][27] ,
         \mem3[230][26] , \mem3[230][25] , \mem3[230][24] , \mem3[229][31] ,
         \mem3[229][30] , \mem3[229][29] , \mem3[229][28] , \mem3[229][27] ,
         \mem3[229][26] , \mem3[229][25] , \mem3[229][24] , \mem3[228][31] ,
         \mem3[228][30] , \mem3[228][29] , \mem3[228][28] , \mem3[228][27] ,
         \mem3[228][26] , \mem3[228][25] , \mem3[228][24] , \mem3[227][31] ,
         \mem3[227][30] , \mem3[227][29] , \mem3[227][28] , \mem3[227][27] ,
         \mem3[227][26] , \mem3[227][25] , \mem3[227][24] , \mem3[226][31] ,
         \mem3[226][30] , \mem3[226][29] , \mem3[226][28] , \mem3[226][27] ,
         \mem3[226][26] , \mem3[226][25] , \mem3[226][24] , \mem3[225][31] ,
         \mem3[225][30] , \mem3[225][29] , \mem3[225][28] , \mem3[225][27] ,
         \mem3[225][26] , \mem3[225][25] , \mem3[225][24] , \mem3[224][31] ,
         \mem3[224][30] , \mem3[224][29] , \mem3[224][28] , \mem3[224][27] ,
         \mem3[224][26] , \mem3[224][25] , \mem3[224][24] , \mem3[223][31] ,
         \mem3[223][30] , \mem3[223][29] , \mem3[223][28] , \mem3[223][27] ,
         \mem3[223][26] , \mem3[223][25] , \mem3[223][24] , \mem3[222][31] ,
         \mem3[222][30] , \mem3[222][29] , \mem3[222][28] , \mem3[222][27] ,
         \mem3[222][26] , \mem3[222][25] , \mem3[222][24] , \mem3[221][31] ,
         \mem3[221][30] , \mem3[221][29] , \mem3[221][28] , \mem3[221][27] ,
         \mem3[221][26] , \mem3[221][25] , \mem3[221][24] , \mem3[220][31] ,
         \mem3[220][30] , \mem3[220][29] , \mem3[220][28] , \mem3[220][27] ,
         \mem3[220][26] , \mem3[220][25] , \mem3[220][24] , \mem3[219][31] ,
         \mem3[219][30] , \mem3[219][29] , \mem3[219][28] , \mem3[219][27] ,
         \mem3[219][26] , \mem3[219][25] , \mem3[219][24] , \mem3[218][31] ,
         \mem3[218][30] , \mem3[218][29] , \mem3[218][28] , \mem3[218][27] ,
         \mem3[218][26] , \mem3[218][25] , \mem3[218][24] , \mem3[217][31] ,
         \mem3[217][30] , \mem3[217][29] , \mem3[217][28] , \mem3[217][27] ,
         \mem3[217][26] , \mem3[217][25] , \mem3[217][24] , \mem3[216][31] ,
         \mem3[216][30] , \mem3[216][29] , \mem3[216][28] , \mem3[216][27] ,
         \mem3[216][26] , \mem3[216][25] , \mem3[216][24] , \mem3[215][31] ,
         \mem3[215][30] , \mem3[215][29] , \mem3[215][28] , \mem3[215][27] ,
         \mem3[215][26] , \mem3[215][25] , \mem3[215][24] , \mem3[214][31] ,
         \mem3[214][30] , \mem3[214][29] , \mem3[214][28] , \mem3[214][27] ,
         \mem3[214][26] , \mem3[214][25] , \mem3[214][24] , \mem3[213][31] ,
         \mem3[213][30] , \mem3[213][29] , \mem3[213][28] , \mem3[213][27] ,
         \mem3[213][26] , \mem3[213][25] , \mem3[213][24] , \mem3[212][31] ,
         \mem3[212][30] , \mem3[212][29] , \mem3[212][28] , \mem3[212][27] ,
         \mem3[212][26] , \mem3[212][25] , \mem3[212][24] , \mem3[211][31] ,
         \mem3[211][30] , \mem3[211][29] , \mem3[211][28] , \mem3[211][27] ,
         \mem3[211][26] , \mem3[211][25] , \mem3[211][24] , \mem3[210][31] ,
         \mem3[210][30] , \mem3[210][29] , \mem3[210][28] , \mem3[210][27] ,
         \mem3[210][26] , \mem3[210][25] , \mem3[210][24] , \mem3[209][31] ,
         \mem3[209][30] , \mem3[209][29] , \mem3[209][28] , \mem3[209][27] ,
         \mem3[209][26] , \mem3[209][25] , \mem3[209][24] , \mem3[208][31] ,
         \mem3[208][30] , \mem3[208][29] , \mem3[208][28] , \mem3[208][27] ,
         \mem3[208][26] , \mem3[208][25] , \mem3[208][24] , \mem3[207][31] ,
         \mem3[207][30] , \mem3[207][29] , \mem3[207][28] , \mem3[207][27] ,
         \mem3[207][26] , \mem3[207][25] , \mem3[207][24] , \mem3[206][31] ,
         \mem3[206][30] , \mem3[206][29] , \mem3[206][28] , \mem3[206][27] ,
         \mem3[206][26] , \mem3[206][25] , \mem3[206][24] , \mem3[205][31] ,
         \mem3[205][30] , \mem3[205][29] , \mem3[205][28] , \mem3[205][27] ,
         \mem3[205][26] , \mem3[205][25] , \mem3[205][24] , \mem3[204][31] ,
         \mem3[204][30] , \mem3[204][29] , \mem3[204][28] , \mem3[204][27] ,
         \mem3[204][26] , \mem3[204][25] , \mem3[204][24] , \mem3[203][31] ,
         \mem3[203][30] , \mem3[203][29] , \mem3[203][28] , \mem3[203][27] ,
         \mem3[203][26] , \mem3[203][25] , \mem3[203][24] , \mem3[202][31] ,
         \mem3[202][30] , \mem3[202][29] , \mem3[202][28] , \mem3[202][27] ,
         \mem3[202][26] , \mem3[202][25] , \mem3[202][24] , \mem3[201][31] ,
         \mem3[201][30] , \mem3[201][29] , \mem3[201][28] , \mem3[201][27] ,
         \mem3[201][26] , \mem3[201][25] , \mem3[201][24] , \mem3[200][31] ,
         \mem3[200][30] , \mem3[200][29] , \mem3[200][28] , \mem3[200][27] ,
         \mem3[200][26] , \mem3[200][25] , \mem3[200][24] , \mem3[199][31] ,
         \mem3[199][30] , \mem3[199][29] , \mem3[199][28] , \mem3[199][27] ,
         \mem3[199][26] , \mem3[199][25] , \mem3[199][24] , \mem3[198][31] ,
         \mem3[198][30] , \mem3[198][29] , \mem3[198][28] , \mem3[198][27] ,
         \mem3[198][26] , \mem3[198][25] , \mem3[198][24] , \mem3[197][31] ,
         \mem3[197][30] , \mem3[197][29] , \mem3[197][28] , \mem3[197][27] ,
         \mem3[197][26] , \mem3[197][25] , \mem3[197][24] , \mem3[196][31] ,
         \mem3[196][30] , \mem3[196][29] , \mem3[196][28] , \mem3[196][27] ,
         \mem3[196][26] , \mem3[196][25] , \mem3[196][24] , \mem3[195][31] ,
         \mem3[195][30] , \mem3[195][29] , \mem3[195][28] , \mem3[195][27] ,
         \mem3[195][26] , \mem3[195][25] , \mem3[195][24] , \mem3[194][31] ,
         \mem3[194][30] , \mem3[194][29] , \mem3[194][28] , \mem3[194][27] ,
         \mem3[194][26] , \mem3[194][25] , \mem3[194][24] , \mem3[193][31] ,
         \mem3[193][30] , \mem3[193][29] , \mem3[193][28] , \mem3[193][27] ,
         \mem3[193][26] , \mem3[193][25] , \mem3[193][24] , \mem3[192][31] ,
         \mem3[192][30] , \mem3[192][29] , \mem3[192][28] , \mem3[192][27] ,
         \mem3[192][26] , \mem3[192][25] , \mem3[192][24] , \mem3[191][31] ,
         \mem3[191][30] , \mem3[191][29] , \mem3[191][28] , \mem3[191][27] ,
         \mem3[191][26] , \mem3[191][25] , \mem3[191][24] , \mem3[190][31] ,
         \mem3[190][30] , \mem3[190][29] , \mem3[190][28] , \mem3[190][27] ,
         \mem3[190][26] , \mem3[190][25] , \mem3[190][24] , \mem3[189][31] ,
         \mem3[189][30] , \mem3[189][29] , \mem3[189][28] , \mem3[189][27] ,
         \mem3[189][26] , \mem3[189][25] , \mem3[189][24] , \mem3[188][31] ,
         \mem3[188][30] , \mem3[188][29] , \mem3[188][28] , \mem3[188][27] ,
         \mem3[188][26] , \mem3[188][25] , \mem3[188][24] , \mem3[187][31] ,
         \mem3[187][30] , \mem3[187][29] , \mem3[187][28] , \mem3[187][27] ,
         \mem3[187][26] , \mem3[187][25] , \mem3[187][24] , \mem3[186][31] ,
         \mem3[186][30] , \mem3[186][29] , \mem3[186][28] , \mem3[186][27] ,
         \mem3[186][26] , \mem3[186][25] , \mem3[186][24] , \mem3[185][31] ,
         \mem3[185][30] , \mem3[185][29] , \mem3[185][28] , \mem3[185][27] ,
         \mem3[185][26] , \mem3[185][25] , \mem3[185][24] , \mem3[184][31] ,
         \mem3[184][30] , \mem3[184][29] , \mem3[184][28] , \mem3[184][27] ,
         \mem3[184][26] , \mem3[184][25] , \mem3[184][24] , \mem3[183][31] ,
         \mem3[183][30] , \mem3[183][29] , \mem3[183][28] , \mem3[183][27] ,
         \mem3[183][26] , \mem3[183][25] , \mem3[183][24] , \mem3[182][31] ,
         \mem3[182][30] , \mem3[182][29] , \mem3[182][28] , \mem3[182][27] ,
         \mem3[182][26] , \mem3[182][25] , \mem3[182][24] , \mem3[181][31] ,
         \mem3[181][30] , \mem3[181][29] , \mem3[181][28] , \mem3[181][27] ,
         \mem3[181][26] , \mem3[181][25] , \mem3[181][24] , \mem3[180][31] ,
         \mem3[180][30] , \mem3[180][29] , \mem3[180][28] , \mem3[180][27] ,
         \mem3[180][26] , \mem3[180][25] , \mem3[180][24] , \mem3[179][31] ,
         \mem3[179][30] , \mem3[179][29] , \mem3[179][28] , \mem3[179][27] ,
         \mem3[179][26] , \mem3[179][25] , \mem3[179][24] , \mem3[178][31] ,
         \mem3[178][30] , \mem3[178][29] , \mem3[178][28] , \mem3[178][27] ,
         \mem3[178][26] , \mem3[178][25] , \mem3[178][24] , \mem3[177][31] ,
         \mem3[177][30] , \mem3[177][29] , \mem3[177][28] , \mem3[177][27] ,
         \mem3[177][26] , \mem3[177][25] , \mem3[177][24] , \mem3[176][31] ,
         \mem3[176][30] , \mem3[176][29] , \mem3[176][28] , \mem3[176][27] ,
         \mem3[176][26] , \mem3[176][25] , \mem3[176][24] , \mem3[175][31] ,
         \mem3[175][30] , \mem3[175][29] , \mem3[175][28] , \mem3[175][27] ,
         \mem3[175][26] , \mem3[175][25] , \mem3[175][24] , \mem3[174][31] ,
         \mem3[174][30] , \mem3[174][29] , \mem3[174][28] , \mem3[174][27] ,
         \mem3[174][26] , \mem3[174][25] , \mem3[174][24] , \mem3[173][31] ,
         \mem3[173][30] , \mem3[173][29] , \mem3[173][28] , \mem3[173][27] ,
         \mem3[173][26] , \mem3[173][25] , \mem3[173][24] , \mem3[172][31] ,
         \mem3[172][30] , \mem3[172][29] , \mem3[172][28] , \mem3[172][27] ,
         \mem3[172][26] , \mem3[172][25] , \mem3[172][24] , \mem3[171][31] ,
         \mem3[171][30] , \mem3[171][29] , \mem3[171][28] , \mem3[171][27] ,
         \mem3[171][26] , \mem3[171][25] , \mem3[171][24] , \mem3[170][31] ,
         \mem3[170][30] , \mem3[170][29] , \mem3[170][28] , \mem3[170][27] ,
         \mem3[170][26] , \mem3[170][25] , \mem3[170][24] , \mem3[169][31] ,
         \mem3[169][30] , \mem3[169][29] , \mem3[169][28] , \mem3[169][27] ,
         \mem3[169][26] , \mem3[169][25] , \mem3[169][24] , \mem3[168][31] ,
         \mem3[168][30] , \mem3[168][29] , \mem3[168][28] , \mem3[168][27] ,
         \mem3[168][26] , \mem3[168][25] , \mem3[168][24] , \mem3[167][31] ,
         \mem3[167][30] , \mem3[167][29] , \mem3[167][28] , \mem3[167][27] ,
         \mem3[167][26] , \mem3[167][25] , \mem3[167][24] , \mem3[166][31] ,
         \mem3[166][30] , \mem3[166][29] , \mem3[166][28] , \mem3[166][27] ,
         \mem3[166][26] , \mem3[166][25] , \mem3[166][24] , \mem3[165][31] ,
         \mem3[165][30] , \mem3[165][29] , \mem3[165][28] , \mem3[165][27] ,
         \mem3[165][26] , \mem3[165][25] , \mem3[165][24] , \mem3[164][31] ,
         \mem3[164][30] , \mem3[164][29] , \mem3[164][28] , \mem3[164][27] ,
         \mem3[164][26] , \mem3[164][25] , \mem3[164][24] , \mem3[163][31] ,
         \mem3[163][30] , \mem3[163][29] , \mem3[163][28] , \mem3[163][27] ,
         \mem3[163][26] , \mem3[163][25] , \mem3[163][24] , \mem3[162][31] ,
         \mem3[162][30] , \mem3[162][29] , \mem3[162][28] , \mem3[162][27] ,
         \mem3[162][26] , \mem3[162][25] , \mem3[162][24] , \mem3[161][31] ,
         \mem3[161][30] , \mem3[161][29] , \mem3[161][28] , \mem3[161][27] ,
         \mem3[161][26] , \mem3[161][25] , \mem3[161][24] , \mem3[160][31] ,
         \mem3[160][30] , \mem3[160][29] , \mem3[160][28] , \mem3[160][27] ,
         \mem3[160][26] , \mem3[160][25] , \mem3[160][24] , \mem3[159][31] ,
         \mem3[159][30] , \mem3[159][29] , \mem3[159][28] , \mem3[159][27] ,
         \mem3[159][26] , \mem3[159][25] , \mem3[159][24] , \mem3[158][31] ,
         \mem3[158][30] , \mem3[158][29] , \mem3[158][28] , \mem3[158][27] ,
         \mem3[158][26] , \mem3[158][25] , \mem3[158][24] , \mem3[157][31] ,
         \mem3[157][30] , \mem3[157][29] , \mem3[157][28] , \mem3[157][27] ,
         \mem3[157][26] , \mem3[157][25] , \mem3[157][24] , \mem3[156][31] ,
         \mem3[156][30] , \mem3[156][29] , \mem3[156][28] , \mem3[156][27] ,
         \mem3[156][26] , \mem3[156][25] , \mem3[156][24] , \mem3[155][31] ,
         \mem3[155][30] , \mem3[155][29] , \mem3[155][28] , \mem3[155][27] ,
         \mem3[155][26] , \mem3[155][25] , \mem3[155][24] , \mem3[154][31] ,
         \mem3[154][30] , \mem3[154][29] , \mem3[154][28] , \mem3[154][27] ,
         \mem3[154][26] , \mem3[154][25] , \mem3[154][24] , \mem3[153][31] ,
         \mem3[153][30] , \mem3[153][29] , \mem3[153][28] , \mem3[153][27] ,
         \mem3[153][26] , \mem3[153][25] , \mem3[153][24] , \mem3[152][31] ,
         \mem3[152][30] , \mem3[152][29] , \mem3[152][28] , \mem3[152][27] ,
         \mem3[152][26] , \mem3[152][25] , \mem3[152][24] , \mem3[151][31] ,
         \mem3[151][30] , \mem3[151][29] , \mem3[151][28] , \mem3[151][27] ,
         \mem3[151][26] , \mem3[151][25] , \mem3[151][24] , \mem3[150][31] ,
         \mem3[150][30] , \mem3[150][29] , \mem3[150][28] , \mem3[150][27] ,
         \mem3[150][26] , \mem3[150][25] , \mem3[150][24] , \mem3[149][31] ,
         \mem3[149][30] , \mem3[149][29] , \mem3[149][28] , \mem3[149][27] ,
         \mem3[149][26] , \mem3[149][25] , \mem3[149][24] , \mem3[148][31] ,
         \mem3[148][30] , \mem3[148][29] , \mem3[148][28] , \mem3[148][27] ,
         \mem3[148][26] , \mem3[148][25] , \mem3[148][24] , \mem3[147][31] ,
         \mem3[147][30] , \mem3[147][29] , \mem3[147][28] , \mem3[147][27] ,
         \mem3[147][26] , \mem3[147][25] , \mem3[147][24] , \mem3[146][31] ,
         \mem3[146][30] , \mem3[146][29] , \mem3[146][28] , \mem3[146][27] ,
         \mem3[146][26] , \mem3[146][25] , \mem3[146][24] , \mem3[145][31] ,
         \mem3[145][30] , \mem3[145][29] , \mem3[145][28] , \mem3[145][27] ,
         \mem3[145][26] , \mem3[145][25] , \mem3[145][24] , \mem3[144][31] ,
         \mem3[144][30] , \mem3[144][29] , \mem3[144][28] , \mem3[144][27] ,
         \mem3[144][26] , \mem3[144][25] , \mem3[144][24] , \mem3[143][31] ,
         \mem3[143][30] , \mem3[143][29] , \mem3[143][28] , \mem3[143][27] ,
         \mem3[143][26] , \mem3[143][25] , \mem3[143][24] , \mem3[142][31] ,
         \mem3[142][30] , \mem3[142][29] , \mem3[142][28] , \mem3[142][27] ,
         \mem3[142][26] , \mem3[142][25] , \mem3[142][24] , \mem3[141][31] ,
         \mem3[141][30] , \mem3[141][29] , \mem3[141][28] , \mem3[141][27] ,
         \mem3[141][26] , \mem3[141][25] , \mem3[141][24] , \mem3[140][31] ,
         \mem3[140][30] , \mem3[140][29] , \mem3[140][28] , \mem3[140][27] ,
         \mem3[140][26] , \mem3[140][25] , \mem3[140][24] , \mem3[139][31] ,
         \mem3[139][30] , \mem3[139][29] , \mem3[139][28] , \mem3[139][27] ,
         \mem3[139][26] , \mem3[139][25] , \mem3[139][24] , \mem3[138][31] ,
         \mem3[138][30] , \mem3[138][29] , \mem3[138][28] , \mem3[138][27] ,
         \mem3[138][26] , \mem3[138][25] , \mem3[138][24] , \mem3[137][31] ,
         \mem3[137][30] , \mem3[137][29] , \mem3[137][28] , \mem3[137][27] ,
         \mem3[137][26] , \mem3[137][25] , \mem3[137][24] , \mem3[136][31] ,
         \mem3[136][30] , \mem3[136][29] , \mem3[136][28] , \mem3[136][27] ,
         \mem3[136][26] , \mem3[136][25] , \mem3[136][24] , \mem3[135][31] ,
         \mem3[135][30] , \mem3[135][29] , \mem3[135][28] , \mem3[135][27] ,
         \mem3[135][26] , \mem3[135][25] , \mem3[135][24] , \mem3[134][31] ,
         \mem3[134][30] , \mem3[134][29] , \mem3[134][28] , \mem3[134][27] ,
         \mem3[134][26] , \mem3[134][25] , \mem3[134][24] , \mem3[133][31] ,
         \mem3[133][30] , \mem3[133][29] , \mem3[133][28] , \mem3[133][27] ,
         \mem3[133][26] , \mem3[133][25] , \mem3[133][24] , \mem3[132][31] ,
         \mem3[132][30] , \mem3[132][29] , \mem3[132][28] , \mem3[132][27] ,
         \mem3[132][26] , \mem3[132][25] , \mem3[132][24] , \mem3[131][31] ,
         \mem3[131][30] , \mem3[131][29] , \mem3[131][28] , \mem3[131][27] ,
         \mem3[131][26] , \mem3[131][25] , \mem3[131][24] , \mem3[130][31] ,
         \mem3[130][30] , \mem3[130][29] , \mem3[130][28] , \mem3[130][27] ,
         \mem3[130][26] , \mem3[130][25] , \mem3[130][24] , \mem3[129][31] ,
         \mem3[129][30] , \mem3[129][29] , \mem3[129][28] , \mem3[129][27] ,
         \mem3[129][26] , \mem3[129][25] , \mem3[129][24] , \mem3[128][31] ,
         \mem3[128][30] , \mem3[128][29] , \mem3[128][28] , \mem3[128][27] ,
         \mem3[128][26] , \mem3[128][25] , \mem3[128][24] , \mem3[127][31] ,
         \mem3[127][30] , \mem3[127][29] , \mem3[127][28] , \mem3[127][27] ,
         \mem3[127][26] , \mem3[127][25] , \mem3[127][24] , \mem3[126][31] ,
         \mem3[126][30] , \mem3[126][29] , \mem3[126][28] , \mem3[126][27] ,
         \mem3[126][26] , \mem3[126][25] , \mem3[126][24] , \mem3[125][31] ,
         \mem3[125][30] , \mem3[125][29] , \mem3[125][28] , \mem3[125][27] ,
         \mem3[125][26] , \mem3[125][25] , \mem3[125][24] , \mem3[124][31] ,
         \mem3[124][30] , \mem3[124][29] , \mem3[124][28] , \mem3[124][27] ,
         \mem3[124][26] , \mem3[124][25] , \mem3[124][24] , \mem3[123][31] ,
         \mem3[123][30] , \mem3[123][29] , \mem3[123][28] , \mem3[123][27] ,
         \mem3[123][26] , \mem3[123][25] , \mem3[123][24] , \mem3[122][31] ,
         \mem3[122][30] , \mem3[122][29] , \mem3[122][28] , \mem3[122][27] ,
         \mem3[122][26] , \mem3[122][25] , \mem3[122][24] , \mem3[121][31] ,
         \mem3[121][30] , \mem3[121][29] , \mem3[121][28] , \mem3[121][27] ,
         \mem3[121][26] , \mem3[121][25] , \mem3[121][24] , \mem3[120][31] ,
         \mem3[120][30] , \mem3[120][29] , \mem3[120][28] , \mem3[120][27] ,
         \mem3[120][26] , \mem3[120][25] , \mem3[120][24] , \mem3[119][31] ,
         \mem3[119][30] , \mem3[119][29] , \mem3[119][28] , \mem3[119][27] ,
         \mem3[119][26] , \mem3[119][25] , \mem3[119][24] , \mem3[118][31] ,
         \mem3[118][30] , \mem3[118][29] , \mem3[118][28] , \mem3[118][27] ,
         \mem3[118][26] , \mem3[118][25] , \mem3[118][24] , \mem3[117][31] ,
         \mem3[117][30] , \mem3[117][29] , \mem3[117][28] , \mem3[117][27] ,
         \mem3[117][26] , \mem3[117][25] , \mem3[117][24] , \mem3[116][31] ,
         \mem3[116][30] , \mem3[116][29] , \mem3[116][28] , \mem3[116][27] ,
         \mem3[116][26] , \mem3[116][25] , \mem3[116][24] , \mem3[115][31] ,
         \mem3[115][30] , \mem3[115][29] , \mem3[115][28] , \mem3[115][27] ,
         \mem3[115][26] , \mem3[115][25] , \mem3[115][24] , \mem3[114][31] ,
         \mem3[114][30] , \mem3[114][29] , \mem3[114][28] , \mem3[114][27] ,
         \mem3[114][26] , \mem3[114][25] , \mem3[114][24] , \mem3[113][31] ,
         \mem3[113][30] , \mem3[113][29] , \mem3[113][28] , \mem3[113][27] ,
         \mem3[113][26] , \mem3[113][25] , \mem3[113][24] , \mem3[112][31] ,
         \mem3[112][30] , \mem3[112][29] , \mem3[112][28] , \mem3[112][27] ,
         \mem3[112][26] , \mem3[112][25] , \mem3[112][24] , \mem3[111][31] ,
         \mem3[111][30] , \mem3[111][29] , \mem3[111][28] , \mem3[111][27] ,
         \mem3[111][26] , \mem3[111][25] , \mem3[111][24] , \mem3[110][31] ,
         \mem3[110][30] , \mem3[110][29] , \mem3[110][28] , \mem3[110][27] ,
         \mem3[110][26] , \mem3[110][25] , \mem3[110][24] , \mem3[109][31] ,
         \mem3[109][30] , \mem3[109][29] , \mem3[109][28] , \mem3[109][27] ,
         \mem3[109][26] , \mem3[109][25] , \mem3[109][24] , \mem3[108][31] ,
         \mem3[108][30] , \mem3[108][29] , \mem3[108][28] , \mem3[108][27] ,
         \mem3[108][26] , \mem3[108][25] , \mem3[108][24] , \mem3[107][31] ,
         \mem3[107][30] , \mem3[107][29] , \mem3[107][28] , \mem3[107][27] ,
         \mem3[107][26] , \mem3[107][25] , \mem3[107][24] , \mem3[106][31] ,
         \mem3[106][30] , \mem3[106][29] , \mem3[106][28] , \mem3[106][27] ,
         \mem3[106][26] , \mem3[106][25] , \mem3[106][24] , \mem3[105][31] ,
         \mem3[105][30] , \mem3[105][29] , \mem3[105][28] , \mem3[105][27] ,
         \mem3[105][26] , \mem3[105][25] , \mem3[105][24] , \mem3[104][31] ,
         \mem3[104][30] , \mem3[104][29] , \mem3[104][28] , \mem3[104][27] ,
         \mem3[104][26] , \mem3[104][25] , \mem3[104][24] , \mem3[103][31] ,
         \mem3[103][30] , \mem3[103][29] , \mem3[103][28] , \mem3[103][27] ,
         \mem3[103][26] , \mem3[103][25] , \mem3[103][24] , \mem3[102][31] ,
         \mem3[102][30] , \mem3[102][29] , \mem3[102][28] , \mem3[102][27] ,
         \mem3[102][26] , \mem3[102][25] , \mem3[102][24] , \mem3[101][31] ,
         \mem3[101][30] , \mem3[101][29] , \mem3[101][28] , \mem3[101][27] ,
         \mem3[101][26] , \mem3[101][25] , \mem3[101][24] , \mem3[100][31] ,
         \mem3[100][30] , \mem3[100][29] , \mem3[100][28] , \mem3[100][27] ,
         \mem3[100][26] , \mem3[100][25] , \mem3[100][24] , \mem3[99][31] ,
         \mem3[99][30] , \mem3[99][29] , \mem3[99][28] , \mem3[99][27] ,
         \mem3[99][26] , \mem3[99][25] , \mem3[99][24] , \mem3[98][31] ,
         \mem3[98][30] , \mem3[98][29] , \mem3[98][28] , \mem3[98][27] ,
         \mem3[98][26] , \mem3[98][25] , \mem3[98][24] , \mem3[97][31] ,
         \mem3[97][30] , \mem3[97][29] , \mem3[97][28] , \mem3[97][27] ,
         \mem3[97][26] , \mem3[97][25] , \mem3[97][24] , \mem3[96][31] ,
         \mem3[96][30] , \mem3[96][29] , \mem3[96][28] , \mem3[96][27] ,
         \mem3[96][26] , \mem3[96][25] , \mem3[96][24] , \mem3[95][31] ,
         \mem3[95][30] , \mem3[95][29] , \mem3[95][28] , \mem3[95][27] ,
         \mem3[95][26] , \mem3[95][25] , \mem3[95][24] , \mem3[94][31] ,
         \mem3[94][30] , \mem3[94][29] , \mem3[94][28] , \mem3[94][27] ,
         \mem3[94][26] , \mem3[94][25] , \mem3[94][24] , \mem3[93][31] ,
         \mem3[93][30] , \mem3[93][29] , \mem3[93][28] , \mem3[93][27] ,
         \mem3[93][26] , \mem3[93][25] , \mem3[93][24] , \mem3[92][31] ,
         \mem3[92][30] , \mem3[92][29] , \mem3[92][28] , \mem3[92][27] ,
         \mem3[92][26] , \mem3[92][25] , \mem3[92][24] , \mem3[91][31] ,
         \mem3[91][30] , \mem3[91][29] , \mem3[91][28] , \mem3[91][27] ,
         \mem3[91][26] , \mem3[91][25] , \mem3[91][24] , \mem3[90][31] ,
         \mem3[90][30] , \mem3[90][29] , \mem3[90][28] , \mem3[90][27] ,
         \mem3[90][26] , \mem3[90][25] , \mem3[90][24] , \mem3[89][31] ,
         \mem3[89][30] , \mem3[89][29] , \mem3[89][28] , \mem3[89][27] ,
         \mem3[89][26] , \mem3[89][25] , \mem3[89][24] , \mem3[88][31] ,
         \mem3[88][30] , \mem3[88][29] , \mem3[88][28] , \mem3[88][27] ,
         \mem3[88][26] , \mem3[88][25] , \mem3[88][24] , \mem3[87][31] ,
         \mem3[87][30] , \mem3[87][29] , \mem3[87][28] , \mem3[87][27] ,
         \mem3[87][26] , \mem3[87][25] , \mem3[87][24] , \mem3[86][31] ,
         \mem3[86][30] , \mem3[86][29] , \mem3[86][28] , \mem3[86][27] ,
         \mem3[86][26] , \mem3[86][25] , \mem3[86][24] , \mem3[85][31] ,
         \mem3[85][30] , \mem3[85][29] , \mem3[85][28] , \mem3[85][27] ,
         \mem3[85][26] , \mem3[85][25] , \mem3[85][24] , \mem3[84][31] ,
         \mem3[84][30] , \mem3[84][29] , \mem3[84][28] , \mem3[84][27] ,
         \mem3[84][26] , \mem3[84][25] , \mem3[84][24] , \mem3[83][31] ,
         \mem3[83][30] , \mem3[83][29] , \mem3[83][28] , \mem3[83][27] ,
         \mem3[83][26] , \mem3[83][25] , \mem3[83][24] , \mem3[82][31] ,
         \mem3[82][30] , \mem3[82][29] , \mem3[82][28] , \mem3[82][27] ,
         \mem3[82][26] , \mem3[82][25] , \mem3[82][24] , \mem3[81][31] ,
         \mem3[81][30] , \mem3[81][29] , \mem3[81][28] , \mem3[81][27] ,
         \mem3[81][26] , \mem3[81][25] , \mem3[81][24] , \mem3[80][31] ,
         \mem3[80][30] , \mem3[80][29] , \mem3[80][28] , \mem3[80][27] ,
         \mem3[80][26] , \mem3[80][25] , \mem3[80][24] , \mem3[79][31] ,
         \mem3[79][30] , \mem3[79][29] , \mem3[79][28] , \mem3[79][27] ,
         \mem3[79][26] , \mem3[79][25] , \mem3[79][24] , \mem3[78][31] ,
         \mem3[78][30] , \mem3[78][29] , \mem3[78][28] , \mem3[78][27] ,
         \mem3[78][26] , \mem3[78][25] , \mem3[78][24] , \mem3[77][31] ,
         \mem3[77][30] , \mem3[77][29] , \mem3[77][28] , \mem3[77][27] ,
         \mem3[77][26] , \mem3[77][25] , \mem3[77][24] , \mem3[76][31] ,
         \mem3[76][30] , \mem3[76][29] , \mem3[76][28] , \mem3[76][27] ,
         \mem3[76][26] , \mem3[76][25] , \mem3[76][24] , \mem3[75][31] ,
         \mem3[75][30] , \mem3[75][29] , \mem3[75][28] , \mem3[75][27] ,
         \mem3[75][26] , \mem3[75][25] , \mem3[75][24] , \mem3[74][31] ,
         \mem3[74][30] , \mem3[74][29] , \mem3[74][28] , \mem3[74][27] ,
         \mem3[74][26] , \mem3[74][25] , \mem3[74][24] , \mem3[73][31] ,
         \mem3[73][30] , \mem3[73][29] , \mem3[73][28] , \mem3[73][27] ,
         \mem3[73][26] , \mem3[73][25] , \mem3[73][24] , \mem3[72][31] ,
         \mem3[72][30] , \mem3[72][29] , \mem3[72][28] , \mem3[72][27] ,
         \mem3[72][26] , \mem3[72][25] , \mem3[72][24] , \mem3[71][31] ,
         \mem3[71][30] , \mem3[71][29] , \mem3[71][28] , \mem3[71][27] ,
         \mem3[71][26] , \mem3[71][25] , \mem3[71][24] , \mem3[70][31] ,
         \mem3[70][30] , \mem3[70][29] , \mem3[70][28] , \mem3[70][27] ,
         \mem3[70][26] , \mem3[70][25] , \mem3[70][24] , \mem3[69][31] ,
         \mem3[69][30] , \mem3[69][29] , \mem3[69][28] , \mem3[69][27] ,
         \mem3[69][26] , \mem3[69][25] , \mem3[69][24] , \mem3[68][31] ,
         \mem3[68][30] , \mem3[68][29] , \mem3[68][28] , \mem3[68][27] ,
         \mem3[68][26] , \mem3[68][25] , \mem3[68][24] , \mem3[67][31] ,
         \mem3[67][30] , \mem3[67][29] , \mem3[67][28] , \mem3[67][27] ,
         \mem3[67][26] , \mem3[67][25] , \mem3[67][24] , \mem3[66][31] ,
         \mem3[66][30] , \mem3[66][29] , \mem3[66][28] , \mem3[66][27] ,
         \mem3[66][26] , \mem3[66][25] , \mem3[66][24] , \mem3[65][31] ,
         \mem3[65][30] , \mem3[65][29] , \mem3[65][28] , \mem3[65][27] ,
         \mem3[65][26] , \mem3[65][25] , \mem3[65][24] , \mem3[64][31] ,
         \mem3[64][30] , \mem3[64][29] , \mem3[64][28] , \mem3[64][27] ,
         \mem3[64][26] , \mem3[64][25] , \mem3[64][24] , \mem3[63][31] ,
         \mem3[63][30] , \mem3[63][29] , \mem3[63][28] , \mem3[63][27] ,
         \mem3[63][26] , \mem3[63][25] , \mem3[63][24] , \mem3[62][31] ,
         \mem3[62][30] , \mem3[62][29] , \mem3[62][28] , \mem3[62][27] ,
         \mem3[62][26] , \mem3[62][25] , \mem3[62][24] , \mem3[61][31] ,
         \mem3[61][30] , \mem3[61][29] , \mem3[61][28] , \mem3[61][27] ,
         \mem3[61][26] , \mem3[61][25] , \mem3[61][24] , \mem3[60][31] ,
         \mem3[60][30] , \mem3[60][29] , \mem3[60][28] , \mem3[60][27] ,
         \mem3[60][26] , \mem3[60][25] , \mem3[60][24] , \mem3[59][31] ,
         \mem3[59][30] , \mem3[59][29] , \mem3[59][28] , \mem3[59][27] ,
         \mem3[59][26] , \mem3[59][25] , \mem3[59][24] , \mem3[58][31] ,
         \mem3[58][30] , \mem3[58][29] , \mem3[58][28] , \mem3[58][27] ,
         \mem3[58][26] , \mem3[58][25] , \mem3[58][24] , \mem3[57][31] ,
         \mem3[57][30] , \mem3[57][29] , \mem3[57][28] , \mem3[57][27] ,
         \mem3[57][26] , \mem3[57][25] , \mem3[57][24] , \mem3[56][31] ,
         \mem3[56][30] , \mem3[56][29] , \mem3[56][28] , \mem3[56][27] ,
         \mem3[56][26] , \mem3[56][25] , \mem3[56][24] , \mem3[55][31] ,
         \mem3[55][30] , \mem3[55][29] , \mem3[55][28] , \mem3[55][27] ,
         \mem3[55][26] , \mem3[55][25] , \mem3[55][24] , \mem3[54][31] ,
         \mem3[54][30] , \mem3[54][29] , \mem3[54][28] , \mem3[54][27] ,
         \mem3[54][26] , \mem3[54][25] , \mem3[54][24] , \mem3[53][31] ,
         \mem3[53][30] , \mem3[53][29] , \mem3[53][28] , \mem3[53][27] ,
         \mem3[53][26] , \mem3[53][25] , \mem3[53][24] , \mem3[52][31] ,
         \mem3[52][30] , \mem3[52][29] , \mem3[52][28] , \mem3[52][27] ,
         \mem3[52][26] , \mem3[52][25] , \mem3[52][24] , \mem3[51][31] ,
         \mem3[51][30] , \mem3[51][29] , \mem3[51][28] , \mem3[51][27] ,
         \mem3[51][26] , \mem3[51][25] , \mem3[51][24] , \mem3[50][31] ,
         \mem3[50][30] , \mem3[50][29] , \mem3[50][28] , \mem3[50][27] ,
         \mem3[50][26] , \mem3[50][25] , \mem3[50][24] , \mem3[49][31] ,
         \mem3[49][30] , \mem3[49][29] , \mem3[49][28] , \mem3[49][27] ,
         \mem3[49][26] , \mem3[49][25] , \mem3[49][24] , \mem3[48][31] ,
         \mem3[48][30] , \mem3[48][29] , \mem3[48][28] , \mem3[48][27] ,
         \mem3[48][26] , \mem3[48][25] , \mem3[48][24] , \mem3[47][31] ,
         \mem3[47][30] , \mem3[47][29] , \mem3[47][28] , \mem3[47][27] ,
         \mem3[47][26] , \mem3[47][25] , \mem3[47][24] , \mem3[46][31] ,
         \mem3[46][30] , \mem3[46][29] , \mem3[46][28] , \mem3[46][27] ,
         \mem3[46][26] , \mem3[46][25] , \mem3[46][24] , \mem3[45][31] ,
         \mem3[45][30] , \mem3[45][29] , \mem3[45][28] , \mem3[45][27] ,
         \mem3[45][26] , \mem3[45][25] , \mem3[45][24] , \mem3[44][31] ,
         \mem3[44][30] , \mem3[44][29] , \mem3[44][28] , \mem3[44][27] ,
         \mem3[44][26] , \mem3[44][25] , \mem3[44][24] , \mem3[43][31] ,
         \mem3[43][30] , \mem3[43][29] , \mem3[43][28] , \mem3[43][27] ,
         \mem3[43][26] , \mem3[43][25] , \mem3[43][24] , \mem3[42][31] ,
         \mem3[42][30] , \mem3[42][29] , \mem3[42][28] , \mem3[42][27] ,
         \mem3[42][26] , \mem3[42][25] , \mem3[42][24] , \mem3[41][31] ,
         \mem3[41][30] , \mem3[41][29] , \mem3[41][28] , \mem3[41][27] ,
         \mem3[41][26] , \mem3[41][25] , \mem3[41][24] , \mem3[40][31] ,
         \mem3[40][30] , \mem3[40][29] , \mem3[40][28] , \mem3[40][27] ,
         \mem3[40][26] , \mem3[40][25] , \mem3[40][24] , \mem3[39][31] ,
         \mem3[39][30] , \mem3[39][29] , \mem3[39][28] , \mem3[39][27] ,
         \mem3[39][26] , \mem3[39][25] , \mem3[39][24] , \mem3[38][31] ,
         \mem3[38][30] , \mem3[38][29] , \mem3[38][28] , \mem3[38][27] ,
         \mem3[38][26] , \mem3[38][25] , \mem3[38][24] , \mem3[37][31] ,
         \mem3[37][30] , \mem3[37][29] , \mem3[37][28] , \mem3[37][27] ,
         \mem3[37][26] , \mem3[37][25] , \mem3[37][24] , \mem3[36][31] ,
         \mem3[36][30] , \mem3[36][29] , \mem3[36][28] , \mem3[36][27] ,
         \mem3[36][26] , \mem3[36][25] , \mem3[36][24] , \mem3[35][31] ,
         \mem3[35][30] , \mem3[35][29] , \mem3[35][28] , \mem3[35][27] ,
         \mem3[35][26] , \mem3[35][25] , \mem3[35][24] , \mem3[34][31] ,
         \mem3[34][30] , \mem3[34][29] , \mem3[34][28] , \mem3[34][27] ,
         \mem3[34][26] , \mem3[34][25] , \mem3[34][24] , \mem3[33][31] ,
         \mem3[33][30] , \mem3[33][29] , \mem3[33][28] , \mem3[33][27] ,
         \mem3[33][26] , \mem3[33][25] , \mem3[33][24] , \mem3[32][31] ,
         \mem3[32][30] , \mem3[32][29] , \mem3[32][28] , \mem3[32][27] ,
         \mem3[32][26] , \mem3[32][25] , \mem3[32][24] , \mem3[31][31] ,
         \mem3[31][30] , \mem3[31][29] , \mem3[31][28] , \mem3[31][27] ,
         \mem3[31][26] , \mem3[31][25] , \mem3[31][24] , \mem3[30][31] ,
         \mem3[30][30] , \mem3[30][29] , \mem3[30][28] , \mem3[30][27] ,
         \mem3[30][26] , \mem3[30][25] , \mem3[30][24] , \mem3[29][31] ,
         \mem3[29][30] , \mem3[29][29] , \mem3[29][28] , \mem3[29][27] ,
         \mem3[29][26] , \mem3[29][25] , \mem3[29][24] , \mem3[28][31] ,
         \mem3[28][30] , \mem3[28][29] , \mem3[28][28] , \mem3[28][27] ,
         \mem3[28][26] , \mem3[28][25] , \mem3[28][24] , \mem3[27][31] ,
         \mem3[27][30] , \mem3[27][29] , \mem3[27][28] , \mem3[27][27] ,
         \mem3[27][26] , \mem3[27][25] , \mem3[27][24] , \mem3[26][31] ,
         \mem3[26][30] , \mem3[26][29] , \mem3[26][28] , \mem3[26][27] ,
         \mem3[26][26] , \mem3[26][25] , \mem3[26][24] , \mem3[25][31] ,
         \mem3[25][30] , \mem3[25][29] , \mem3[25][28] , \mem3[25][27] ,
         \mem3[25][26] , \mem3[25][25] , \mem3[25][24] , \mem3[24][31] ,
         \mem3[24][30] , \mem3[24][29] , \mem3[24][28] , \mem3[24][27] ,
         \mem3[24][26] , \mem3[24][25] , \mem3[24][24] , \mem3[23][31] ,
         \mem3[23][30] , \mem3[23][29] , \mem3[23][28] , \mem3[23][27] ,
         \mem3[23][26] , \mem3[23][25] , \mem3[23][24] , \mem3[22][31] ,
         \mem3[22][30] , \mem3[22][29] , \mem3[22][28] , \mem3[22][27] ,
         \mem3[22][26] , \mem3[22][25] , \mem3[22][24] , \mem3[21][31] ,
         \mem3[21][30] , \mem3[21][29] , \mem3[21][28] , \mem3[21][27] ,
         \mem3[21][26] , \mem3[21][25] , \mem3[21][24] , \mem3[20][31] ,
         \mem3[20][30] , \mem3[20][29] , \mem3[20][28] , \mem3[20][27] ,
         \mem3[20][26] , \mem3[20][25] , \mem3[20][24] , \mem3[19][31] ,
         \mem3[19][30] , \mem3[19][29] , \mem3[19][28] , \mem3[19][27] ,
         \mem3[19][26] , \mem3[19][25] , \mem3[19][24] , \mem3[18][31] ,
         \mem3[18][30] , \mem3[18][29] , \mem3[18][28] , \mem3[18][27] ,
         \mem3[18][26] , \mem3[18][25] , \mem3[18][24] , \mem3[17][31] ,
         \mem3[17][30] , \mem3[17][29] , \mem3[17][28] , \mem3[17][27] ,
         \mem3[17][26] , \mem3[17][25] , \mem3[17][24] , \mem3[16][31] ,
         \mem3[16][30] , \mem3[16][29] , \mem3[16][28] , \mem3[16][27] ,
         \mem3[16][26] , \mem3[16][25] , \mem3[16][24] , \mem3[15][31] ,
         \mem3[15][30] , \mem3[15][29] , \mem3[15][28] , \mem3[15][27] ,
         \mem3[15][26] , \mem3[15][25] , \mem3[15][24] , \mem3[14][31] ,
         \mem3[14][30] , \mem3[14][29] , \mem3[14][28] , \mem3[14][27] ,
         \mem3[14][26] , \mem3[14][25] , \mem3[14][24] , \mem3[13][31] ,
         \mem3[13][30] , \mem3[13][29] , \mem3[13][28] , \mem3[13][27] ,
         \mem3[13][26] , \mem3[13][25] , \mem3[13][24] , \mem3[12][31] ,
         \mem3[12][30] , \mem3[12][29] , \mem3[12][28] , \mem3[12][27] ,
         \mem3[12][26] , \mem3[12][25] , \mem3[12][24] , \mem3[11][31] ,
         \mem3[11][30] , \mem3[11][29] , \mem3[11][28] , \mem3[11][27] ,
         \mem3[11][26] , \mem3[11][25] , \mem3[11][24] , \mem3[10][31] ,
         \mem3[10][30] , \mem3[10][29] , \mem3[10][28] , \mem3[10][27] ,
         \mem3[10][26] , \mem3[10][25] , \mem3[10][24] , \mem3[9][31] ,
         \mem3[9][30] , \mem3[9][29] , \mem3[9][28] , \mem3[9][27] ,
         \mem3[9][26] , \mem3[9][25] , \mem3[9][24] , \mem3[8][31] ,
         \mem3[8][30] , \mem3[8][29] , \mem3[8][28] , \mem3[8][27] ,
         \mem3[8][26] , \mem3[8][25] , \mem3[8][24] , \mem3[7][31] ,
         \mem3[7][30] , \mem3[7][29] , \mem3[7][28] , \mem3[7][27] ,
         \mem3[7][26] , \mem3[7][25] , \mem3[7][24] , \mem3[6][31] ,
         \mem3[6][30] , \mem3[6][29] , \mem3[6][28] , \mem3[6][27] ,
         \mem3[6][26] , \mem3[6][25] , \mem3[6][24] , \mem3[5][31] ,
         \mem3[5][30] , \mem3[5][29] , \mem3[5][28] , \mem3[5][27] ,
         \mem3[5][26] , \mem3[5][25] , \mem3[5][24] , \mem3[4][31] ,
         \mem3[4][30] , \mem3[4][29] , \mem3[4][28] , \mem3[4][27] ,
         \mem3[4][26] , \mem3[4][25] , \mem3[4][24] , \mem3[3][31] ,
         \mem3[3][30] , \mem3[3][29] , \mem3[3][28] , \mem3[3][27] ,
         \mem3[3][26] , \mem3[3][25] , \mem3[3][24] , \mem3[2][31] ,
         \mem3[2][30] , \mem3[2][29] , \mem3[2][28] , \mem3[2][27] ,
         \mem3[2][26] , \mem3[2][25] , \mem3[2][24] , \mem3[1][31] ,
         \mem3[1][30] , \mem3[1][29] , \mem3[1][28] , \mem3[1][27] ,
         \mem3[1][26] , \mem3[1][25] , \mem3[1][24] , \mem3[0][31] ,
         \mem3[0][30] , \mem3[0][29] , \mem3[0][28] , \mem3[0][27] ,
         \mem3[0][26] , \mem3[0][25] , \mem3[0][24] , \mem2[255][23] ,
         \mem2[255][22] , \mem2[255][21] , \mem2[255][20] , \mem2[255][19] ,
         \mem2[255][18] , \mem2[255][17] , \mem2[255][16] , \mem2[254][23] ,
         \mem2[254][22] , \mem2[254][21] , \mem2[254][20] , \mem2[254][19] ,
         \mem2[254][18] , \mem2[254][17] , \mem2[254][16] , \mem2[253][23] ,
         \mem2[253][22] , \mem2[253][21] , \mem2[253][20] , \mem2[253][19] ,
         \mem2[253][18] , \mem2[253][17] , \mem2[253][16] , \mem2[252][23] ,
         \mem2[252][22] , \mem2[252][21] , \mem2[252][20] , \mem2[252][19] ,
         \mem2[252][18] , \mem2[252][17] , \mem2[252][16] , \mem2[251][23] ,
         \mem2[251][22] , \mem2[251][21] , \mem2[251][20] , \mem2[251][19] ,
         \mem2[251][18] , \mem2[251][17] , \mem2[251][16] , \mem2[250][23] ,
         \mem2[250][22] , \mem2[250][21] , \mem2[250][20] , \mem2[250][19] ,
         \mem2[250][18] , \mem2[250][17] , \mem2[250][16] , \mem2[249][23] ,
         \mem2[249][22] , \mem2[249][21] , \mem2[249][20] , \mem2[249][19] ,
         \mem2[249][18] , \mem2[249][17] , \mem2[249][16] , \mem2[248][23] ,
         \mem2[248][22] , \mem2[248][21] , \mem2[248][20] , \mem2[248][19] ,
         \mem2[248][18] , \mem2[248][17] , \mem2[248][16] , \mem2[247][23] ,
         \mem2[247][22] , \mem2[247][21] , \mem2[247][20] , \mem2[247][19] ,
         \mem2[247][18] , \mem2[247][17] , \mem2[247][16] , \mem2[246][23] ,
         \mem2[246][22] , \mem2[246][21] , \mem2[246][20] , \mem2[246][19] ,
         \mem2[246][18] , \mem2[246][17] , \mem2[246][16] , \mem2[245][23] ,
         \mem2[245][22] , \mem2[245][21] , \mem2[245][20] , \mem2[245][19] ,
         \mem2[245][18] , \mem2[245][17] , \mem2[245][16] , \mem2[244][23] ,
         \mem2[244][22] , \mem2[244][21] , \mem2[244][20] , \mem2[244][19] ,
         \mem2[244][18] , \mem2[244][17] , \mem2[244][16] , \mem2[243][23] ,
         \mem2[243][22] , \mem2[243][21] , \mem2[243][20] , \mem2[243][19] ,
         \mem2[243][18] , \mem2[243][17] , \mem2[243][16] , \mem2[242][23] ,
         \mem2[242][22] , \mem2[242][21] , \mem2[242][20] , \mem2[242][19] ,
         \mem2[242][18] , \mem2[242][17] , \mem2[242][16] , \mem2[241][23] ,
         \mem2[241][22] , \mem2[241][21] , \mem2[241][20] , \mem2[241][19] ,
         \mem2[241][18] , \mem2[241][17] , \mem2[241][16] , \mem2[240][23] ,
         \mem2[240][22] , \mem2[240][21] , \mem2[240][20] , \mem2[240][19] ,
         \mem2[240][18] , \mem2[240][17] , \mem2[240][16] , \mem2[239][23] ,
         \mem2[239][22] , \mem2[239][21] , \mem2[239][20] , \mem2[239][19] ,
         \mem2[239][18] , \mem2[239][17] , \mem2[239][16] , \mem2[238][23] ,
         \mem2[238][22] , \mem2[238][21] , \mem2[238][20] , \mem2[238][19] ,
         \mem2[238][18] , \mem2[238][17] , \mem2[238][16] , \mem2[237][23] ,
         \mem2[237][22] , \mem2[237][21] , \mem2[237][20] , \mem2[237][19] ,
         \mem2[237][18] , \mem2[237][17] , \mem2[237][16] , \mem2[236][23] ,
         \mem2[236][22] , \mem2[236][21] , \mem2[236][20] , \mem2[236][19] ,
         \mem2[236][18] , \mem2[236][17] , \mem2[236][16] , \mem2[235][23] ,
         \mem2[235][22] , \mem2[235][21] , \mem2[235][20] , \mem2[235][19] ,
         \mem2[235][18] , \mem2[235][17] , \mem2[235][16] , \mem2[234][23] ,
         \mem2[234][22] , \mem2[234][21] , \mem2[234][20] , \mem2[234][19] ,
         \mem2[234][18] , \mem2[234][17] , \mem2[234][16] , \mem2[233][23] ,
         \mem2[233][22] , \mem2[233][21] , \mem2[233][20] , \mem2[233][19] ,
         \mem2[233][18] , \mem2[233][17] , \mem2[233][16] , \mem2[232][23] ,
         \mem2[232][22] , \mem2[232][21] , \mem2[232][20] , \mem2[232][19] ,
         \mem2[232][18] , \mem2[232][17] , \mem2[232][16] , \mem2[231][23] ,
         \mem2[231][22] , \mem2[231][21] , \mem2[231][20] , \mem2[231][19] ,
         \mem2[231][18] , \mem2[231][17] , \mem2[231][16] , \mem2[230][23] ,
         \mem2[230][22] , \mem2[230][21] , \mem2[230][20] , \mem2[230][19] ,
         \mem2[230][18] , \mem2[230][17] , \mem2[230][16] , \mem2[229][23] ,
         \mem2[229][22] , \mem2[229][21] , \mem2[229][20] , \mem2[229][19] ,
         \mem2[229][18] , \mem2[229][17] , \mem2[229][16] , \mem2[228][23] ,
         \mem2[228][22] , \mem2[228][21] , \mem2[228][20] , \mem2[228][19] ,
         \mem2[228][18] , \mem2[228][17] , \mem2[228][16] , \mem2[227][23] ,
         \mem2[227][22] , \mem2[227][21] , \mem2[227][20] , \mem2[227][19] ,
         \mem2[227][18] , \mem2[227][17] , \mem2[227][16] , \mem2[226][23] ,
         \mem2[226][22] , \mem2[226][21] , \mem2[226][20] , \mem2[226][19] ,
         \mem2[226][18] , \mem2[226][17] , \mem2[226][16] , \mem2[225][23] ,
         \mem2[225][22] , \mem2[225][21] , \mem2[225][20] , \mem2[225][19] ,
         \mem2[225][18] , \mem2[225][17] , \mem2[225][16] , \mem2[224][23] ,
         \mem2[224][22] , \mem2[224][21] , \mem2[224][20] , \mem2[224][19] ,
         \mem2[224][18] , \mem2[224][17] , \mem2[224][16] , \mem2[223][23] ,
         \mem2[223][22] , \mem2[223][21] , \mem2[223][20] , \mem2[223][19] ,
         \mem2[223][18] , \mem2[223][17] , \mem2[223][16] , \mem2[222][23] ,
         \mem2[222][22] , \mem2[222][21] , \mem2[222][20] , \mem2[222][19] ,
         \mem2[222][18] , \mem2[222][17] , \mem2[222][16] , \mem2[221][23] ,
         \mem2[221][22] , \mem2[221][21] , \mem2[221][20] , \mem2[221][19] ,
         \mem2[221][18] , \mem2[221][17] , \mem2[221][16] , \mem2[220][23] ,
         \mem2[220][22] , \mem2[220][21] , \mem2[220][20] , \mem2[220][19] ,
         \mem2[220][18] , \mem2[220][17] , \mem2[220][16] , \mem2[219][23] ,
         \mem2[219][22] , \mem2[219][21] , \mem2[219][20] , \mem2[219][19] ,
         \mem2[219][18] , \mem2[219][17] , \mem2[219][16] , \mem2[218][23] ,
         \mem2[218][22] , \mem2[218][21] , \mem2[218][20] , \mem2[218][19] ,
         \mem2[218][18] , \mem2[218][17] , \mem2[218][16] , \mem2[217][23] ,
         \mem2[217][22] , \mem2[217][21] , \mem2[217][20] , \mem2[217][19] ,
         \mem2[217][18] , \mem2[217][17] , \mem2[217][16] , \mem2[216][23] ,
         \mem2[216][22] , \mem2[216][21] , \mem2[216][20] , \mem2[216][19] ,
         \mem2[216][18] , \mem2[216][17] , \mem2[216][16] , \mem2[215][23] ,
         \mem2[215][22] , \mem2[215][21] , \mem2[215][20] , \mem2[215][19] ,
         \mem2[215][18] , \mem2[215][17] , \mem2[215][16] , \mem2[214][23] ,
         \mem2[214][22] , \mem2[214][21] , \mem2[214][20] , \mem2[214][19] ,
         \mem2[214][18] , \mem2[214][17] , \mem2[214][16] , \mem2[213][23] ,
         \mem2[213][22] , \mem2[213][21] , \mem2[213][20] , \mem2[213][19] ,
         \mem2[213][18] , \mem2[213][17] , \mem2[213][16] , \mem2[212][23] ,
         \mem2[212][22] , \mem2[212][21] , \mem2[212][20] , \mem2[212][19] ,
         \mem2[212][18] , \mem2[212][17] , \mem2[212][16] , \mem2[211][23] ,
         \mem2[211][22] , \mem2[211][21] , \mem2[211][20] , \mem2[211][19] ,
         \mem2[211][18] , \mem2[211][17] , \mem2[211][16] , \mem2[210][23] ,
         \mem2[210][22] , \mem2[210][21] , \mem2[210][20] , \mem2[210][19] ,
         \mem2[210][18] , \mem2[210][17] , \mem2[210][16] , \mem2[209][23] ,
         \mem2[209][22] , \mem2[209][21] , \mem2[209][20] , \mem2[209][19] ,
         \mem2[209][18] , \mem2[209][17] , \mem2[209][16] , \mem2[208][23] ,
         \mem2[208][22] , \mem2[208][21] , \mem2[208][20] , \mem2[208][19] ,
         \mem2[208][18] , \mem2[208][17] , \mem2[208][16] , \mem2[207][23] ,
         \mem2[207][22] , \mem2[207][21] , \mem2[207][20] , \mem2[207][19] ,
         \mem2[207][18] , \mem2[207][17] , \mem2[207][16] , \mem2[206][23] ,
         \mem2[206][22] , \mem2[206][21] , \mem2[206][20] , \mem2[206][19] ,
         \mem2[206][18] , \mem2[206][17] , \mem2[206][16] , \mem2[205][23] ,
         \mem2[205][22] , \mem2[205][21] , \mem2[205][20] , \mem2[205][19] ,
         \mem2[205][18] , \mem2[205][17] , \mem2[205][16] , \mem2[204][23] ,
         \mem2[204][22] , \mem2[204][21] , \mem2[204][20] , \mem2[204][19] ,
         \mem2[204][18] , \mem2[204][17] , \mem2[204][16] , \mem2[203][23] ,
         \mem2[203][22] , \mem2[203][21] , \mem2[203][20] , \mem2[203][19] ,
         \mem2[203][18] , \mem2[203][17] , \mem2[203][16] , \mem2[202][23] ,
         \mem2[202][22] , \mem2[202][21] , \mem2[202][20] , \mem2[202][19] ,
         \mem2[202][18] , \mem2[202][17] , \mem2[202][16] , \mem2[201][23] ,
         \mem2[201][22] , \mem2[201][21] , \mem2[201][20] , \mem2[201][19] ,
         \mem2[201][18] , \mem2[201][17] , \mem2[201][16] , \mem2[200][23] ,
         \mem2[200][22] , \mem2[200][21] , \mem2[200][20] , \mem2[200][19] ,
         \mem2[200][18] , \mem2[200][17] , \mem2[200][16] , \mem2[199][23] ,
         \mem2[199][22] , \mem2[199][21] , \mem2[199][20] , \mem2[199][19] ,
         \mem2[199][18] , \mem2[199][17] , \mem2[199][16] , \mem2[198][23] ,
         \mem2[198][22] , \mem2[198][21] , \mem2[198][20] , \mem2[198][19] ,
         \mem2[198][18] , \mem2[198][17] , \mem2[198][16] , \mem2[197][23] ,
         \mem2[197][22] , \mem2[197][21] , \mem2[197][20] , \mem2[197][19] ,
         \mem2[197][18] , \mem2[197][17] , \mem2[197][16] , \mem2[196][23] ,
         \mem2[196][22] , \mem2[196][21] , \mem2[196][20] , \mem2[196][19] ,
         \mem2[196][18] , \mem2[196][17] , \mem2[196][16] , \mem2[195][23] ,
         \mem2[195][22] , \mem2[195][21] , \mem2[195][20] , \mem2[195][19] ,
         \mem2[195][18] , \mem2[195][17] , \mem2[195][16] , \mem2[194][23] ,
         \mem2[194][22] , \mem2[194][21] , \mem2[194][20] , \mem2[194][19] ,
         \mem2[194][18] , \mem2[194][17] , \mem2[194][16] , \mem2[193][23] ,
         \mem2[193][22] , \mem2[193][21] , \mem2[193][20] , \mem2[193][19] ,
         \mem2[193][18] , \mem2[193][17] , \mem2[193][16] , \mem2[192][23] ,
         \mem2[192][22] , \mem2[192][21] , \mem2[192][20] , \mem2[192][19] ,
         \mem2[192][18] , \mem2[192][17] , \mem2[192][16] , \mem2[191][23] ,
         \mem2[191][22] , \mem2[191][21] , \mem2[191][20] , \mem2[191][19] ,
         \mem2[191][18] , \mem2[191][17] , \mem2[191][16] , \mem2[190][23] ,
         \mem2[190][22] , \mem2[190][21] , \mem2[190][20] , \mem2[190][19] ,
         \mem2[190][18] , \mem2[190][17] , \mem2[190][16] , \mem2[189][23] ,
         \mem2[189][22] , \mem2[189][21] , \mem2[189][20] , \mem2[189][19] ,
         \mem2[189][18] , \mem2[189][17] , \mem2[189][16] , \mem2[188][23] ,
         \mem2[188][22] , \mem2[188][21] , \mem2[188][20] , \mem2[188][19] ,
         \mem2[188][18] , \mem2[188][17] , \mem2[188][16] , \mem2[187][23] ,
         \mem2[187][22] , \mem2[187][21] , \mem2[187][20] , \mem2[187][19] ,
         \mem2[187][18] , \mem2[187][17] , \mem2[187][16] , \mem2[186][23] ,
         \mem2[186][22] , \mem2[186][21] , \mem2[186][20] , \mem2[186][19] ,
         \mem2[186][18] , \mem2[186][17] , \mem2[186][16] , \mem2[185][23] ,
         \mem2[185][22] , \mem2[185][21] , \mem2[185][20] , \mem2[185][19] ,
         \mem2[185][18] , \mem2[185][17] , \mem2[185][16] , \mem2[184][23] ,
         \mem2[184][22] , \mem2[184][21] , \mem2[184][20] , \mem2[184][19] ,
         \mem2[184][18] , \mem2[184][17] , \mem2[184][16] , \mem2[183][23] ,
         \mem2[183][22] , \mem2[183][21] , \mem2[183][20] , \mem2[183][19] ,
         \mem2[183][18] , \mem2[183][17] , \mem2[183][16] , \mem2[182][23] ,
         \mem2[182][22] , \mem2[182][21] , \mem2[182][20] , \mem2[182][19] ,
         \mem2[182][18] , \mem2[182][17] , \mem2[182][16] , \mem2[181][23] ,
         \mem2[181][22] , \mem2[181][21] , \mem2[181][20] , \mem2[181][19] ,
         \mem2[181][18] , \mem2[181][17] , \mem2[181][16] , \mem2[180][23] ,
         \mem2[180][22] , \mem2[180][21] , \mem2[180][20] , \mem2[180][19] ,
         \mem2[180][18] , \mem2[180][17] , \mem2[180][16] , \mem2[179][23] ,
         \mem2[179][22] , \mem2[179][21] , \mem2[179][20] , \mem2[179][19] ,
         \mem2[179][18] , \mem2[179][17] , \mem2[179][16] , \mem2[178][23] ,
         \mem2[178][22] , \mem2[178][21] , \mem2[178][20] , \mem2[178][19] ,
         \mem2[178][18] , \mem2[178][17] , \mem2[178][16] , \mem2[177][23] ,
         \mem2[177][22] , \mem2[177][21] , \mem2[177][20] , \mem2[177][19] ,
         \mem2[177][18] , \mem2[177][17] , \mem2[177][16] , \mem2[176][23] ,
         \mem2[176][22] , \mem2[176][21] , \mem2[176][20] , \mem2[176][19] ,
         \mem2[176][18] , \mem2[176][17] , \mem2[176][16] , \mem2[175][23] ,
         \mem2[175][22] , \mem2[175][21] , \mem2[175][20] , \mem2[175][19] ,
         \mem2[175][18] , \mem2[175][17] , \mem2[175][16] , \mem2[174][23] ,
         \mem2[174][22] , \mem2[174][21] , \mem2[174][20] , \mem2[174][19] ,
         \mem2[174][18] , \mem2[174][17] , \mem2[174][16] , \mem2[173][23] ,
         \mem2[173][22] , \mem2[173][21] , \mem2[173][20] , \mem2[173][19] ,
         \mem2[173][18] , \mem2[173][17] , \mem2[173][16] , \mem2[172][23] ,
         \mem2[172][22] , \mem2[172][21] , \mem2[172][20] , \mem2[172][19] ,
         \mem2[172][18] , \mem2[172][17] , \mem2[172][16] , \mem2[171][23] ,
         \mem2[171][22] , \mem2[171][21] , \mem2[171][20] , \mem2[171][19] ,
         \mem2[171][18] , \mem2[171][17] , \mem2[171][16] , \mem2[170][23] ,
         \mem2[170][22] , \mem2[170][21] , \mem2[170][20] , \mem2[170][19] ,
         \mem2[170][18] , \mem2[170][17] , \mem2[170][16] , \mem2[169][23] ,
         \mem2[169][22] , \mem2[169][21] , \mem2[169][20] , \mem2[169][19] ,
         \mem2[169][18] , \mem2[169][17] , \mem2[169][16] , \mem2[168][23] ,
         \mem2[168][22] , \mem2[168][21] , \mem2[168][20] , \mem2[168][19] ,
         \mem2[168][18] , \mem2[168][17] , \mem2[168][16] , \mem2[167][23] ,
         \mem2[167][22] , \mem2[167][21] , \mem2[167][20] , \mem2[167][19] ,
         \mem2[167][18] , \mem2[167][17] , \mem2[167][16] , \mem2[166][23] ,
         \mem2[166][22] , \mem2[166][21] , \mem2[166][20] , \mem2[166][19] ,
         \mem2[166][18] , \mem2[166][17] , \mem2[166][16] , \mem2[165][23] ,
         \mem2[165][22] , \mem2[165][21] , \mem2[165][20] , \mem2[165][19] ,
         \mem2[165][18] , \mem2[165][17] , \mem2[165][16] , \mem2[164][23] ,
         \mem2[164][22] , \mem2[164][21] , \mem2[164][20] , \mem2[164][19] ,
         \mem2[164][18] , \mem2[164][17] , \mem2[164][16] , \mem2[163][23] ,
         \mem2[163][22] , \mem2[163][21] , \mem2[163][20] , \mem2[163][19] ,
         \mem2[163][18] , \mem2[163][17] , \mem2[163][16] , \mem2[162][23] ,
         \mem2[162][22] , \mem2[162][21] , \mem2[162][20] , \mem2[162][19] ,
         \mem2[162][18] , \mem2[162][17] , \mem2[162][16] , \mem2[161][23] ,
         \mem2[161][22] , \mem2[161][21] , \mem2[161][20] , \mem2[161][19] ,
         \mem2[161][18] , \mem2[161][17] , \mem2[161][16] , \mem2[160][23] ,
         \mem2[160][22] , \mem2[160][21] , \mem2[160][20] , \mem2[160][19] ,
         \mem2[160][18] , \mem2[160][17] , \mem2[160][16] , \mem2[159][23] ,
         \mem2[159][22] , \mem2[159][21] , \mem2[159][20] , \mem2[159][19] ,
         \mem2[159][18] , \mem2[159][17] , \mem2[159][16] , \mem2[158][23] ,
         \mem2[158][22] , \mem2[158][21] , \mem2[158][20] , \mem2[158][19] ,
         \mem2[158][18] , \mem2[158][17] , \mem2[158][16] , \mem2[157][23] ,
         \mem2[157][22] , \mem2[157][21] , \mem2[157][20] , \mem2[157][19] ,
         \mem2[157][18] , \mem2[157][17] , \mem2[157][16] , \mem2[156][23] ,
         \mem2[156][22] , \mem2[156][21] , \mem2[156][20] , \mem2[156][19] ,
         \mem2[156][18] , \mem2[156][17] , \mem2[156][16] , \mem2[155][23] ,
         \mem2[155][22] , \mem2[155][21] , \mem2[155][20] , \mem2[155][19] ,
         \mem2[155][18] , \mem2[155][17] , \mem2[155][16] , \mem2[154][23] ,
         \mem2[154][22] , \mem2[154][21] , \mem2[154][20] , \mem2[154][19] ,
         \mem2[154][18] , \mem2[154][17] , \mem2[154][16] , \mem2[153][23] ,
         \mem2[153][22] , \mem2[153][21] , \mem2[153][20] , \mem2[153][19] ,
         \mem2[153][18] , \mem2[153][17] , \mem2[153][16] , \mem2[152][23] ,
         \mem2[152][22] , \mem2[152][21] , \mem2[152][20] , \mem2[152][19] ,
         \mem2[152][18] , \mem2[152][17] , \mem2[152][16] , \mem2[151][23] ,
         \mem2[151][22] , \mem2[151][21] , \mem2[151][20] , \mem2[151][19] ,
         \mem2[151][18] , \mem2[151][17] , \mem2[151][16] , \mem2[150][23] ,
         \mem2[150][22] , \mem2[150][21] , \mem2[150][20] , \mem2[150][19] ,
         \mem2[150][18] , \mem2[150][17] , \mem2[150][16] , \mem2[149][23] ,
         \mem2[149][22] , \mem2[149][21] , \mem2[149][20] , \mem2[149][19] ,
         \mem2[149][18] , \mem2[149][17] , \mem2[149][16] , \mem2[148][23] ,
         \mem2[148][22] , \mem2[148][21] , \mem2[148][20] , \mem2[148][19] ,
         \mem2[148][18] , \mem2[148][17] , \mem2[148][16] , \mem2[147][23] ,
         \mem2[147][22] , \mem2[147][21] , \mem2[147][20] , \mem2[147][19] ,
         \mem2[147][18] , \mem2[147][17] , \mem2[147][16] , \mem2[146][23] ,
         \mem2[146][22] , \mem2[146][21] , \mem2[146][20] , \mem2[146][19] ,
         \mem2[146][18] , \mem2[146][17] , \mem2[146][16] , \mem2[145][23] ,
         \mem2[145][22] , \mem2[145][21] , \mem2[145][20] , \mem2[145][19] ,
         \mem2[145][18] , \mem2[145][17] , \mem2[145][16] , \mem2[144][23] ,
         \mem2[144][22] , \mem2[144][21] , \mem2[144][20] , \mem2[144][19] ,
         \mem2[144][18] , \mem2[144][17] , \mem2[144][16] , \mem2[143][23] ,
         \mem2[143][22] , \mem2[143][21] , \mem2[143][20] , \mem2[143][19] ,
         \mem2[143][18] , \mem2[143][17] , \mem2[143][16] , \mem2[142][23] ,
         \mem2[142][22] , \mem2[142][21] , \mem2[142][20] , \mem2[142][19] ,
         \mem2[142][18] , \mem2[142][17] , \mem2[142][16] , \mem2[141][23] ,
         \mem2[141][22] , \mem2[141][21] , \mem2[141][20] , \mem2[141][19] ,
         \mem2[141][18] , \mem2[141][17] , \mem2[141][16] , \mem2[140][23] ,
         \mem2[140][22] , \mem2[140][21] , \mem2[140][20] , \mem2[140][19] ,
         \mem2[140][18] , \mem2[140][17] , \mem2[140][16] , \mem2[139][23] ,
         \mem2[139][22] , \mem2[139][21] , \mem2[139][20] , \mem2[139][19] ,
         \mem2[139][18] , \mem2[139][17] , \mem2[139][16] , \mem2[138][23] ,
         \mem2[138][22] , \mem2[138][21] , \mem2[138][20] , \mem2[138][19] ,
         \mem2[138][18] , \mem2[138][17] , \mem2[138][16] , \mem2[137][23] ,
         \mem2[137][22] , \mem2[137][21] , \mem2[137][20] , \mem2[137][19] ,
         \mem2[137][18] , \mem2[137][17] , \mem2[137][16] , \mem2[136][23] ,
         \mem2[136][22] , \mem2[136][21] , \mem2[136][20] , \mem2[136][19] ,
         \mem2[136][18] , \mem2[136][17] , \mem2[136][16] , \mem2[135][23] ,
         \mem2[135][22] , \mem2[135][21] , \mem2[135][20] , \mem2[135][19] ,
         \mem2[135][18] , \mem2[135][17] , \mem2[135][16] , \mem2[134][23] ,
         \mem2[134][22] , \mem2[134][21] , \mem2[134][20] , \mem2[134][19] ,
         \mem2[134][18] , \mem2[134][17] , \mem2[134][16] , \mem2[133][23] ,
         \mem2[133][22] , \mem2[133][21] , \mem2[133][20] , \mem2[133][19] ,
         \mem2[133][18] , \mem2[133][17] , \mem2[133][16] , \mem2[132][23] ,
         \mem2[132][22] , \mem2[132][21] , \mem2[132][20] , \mem2[132][19] ,
         \mem2[132][18] , \mem2[132][17] , \mem2[132][16] , \mem2[131][23] ,
         \mem2[131][22] , \mem2[131][21] , \mem2[131][20] , \mem2[131][19] ,
         \mem2[131][18] , \mem2[131][17] , \mem2[131][16] , \mem2[130][23] ,
         \mem2[130][22] , \mem2[130][21] , \mem2[130][20] , \mem2[130][19] ,
         \mem2[130][18] , \mem2[130][17] , \mem2[130][16] , \mem2[129][23] ,
         \mem2[129][22] , \mem2[129][21] , \mem2[129][20] , \mem2[129][19] ,
         \mem2[129][18] , \mem2[129][17] , \mem2[129][16] , \mem2[128][23] ,
         \mem2[128][22] , \mem2[128][21] , \mem2[128][20] , \mem2[128][19] ,
         \mem2[128][18] , \mem2[128][17] , \mem2[128][16] , \mem2[127][23] ,
         \mem2[127][22] , \mem2[127][21] , \mem2[127][20] , \mem2[127][19] ,
         \mem2[127][18] , \mem2[127][17] , \mem2[127][16] , \mem2[126][23] ,
         \mem2[126][22] , \mem2[126][21] , \mem2[126][20] , \mem2[126][19] ,
         \mem2[126][18] , \mem2[126][17] , \mem2[126][16] , \mem2[125][23] ,
         \mem2[125][22] , \mem2[125][21] , \mem2[125][20] , \mem2[125][19] ,
         \mem2[125][18] , \mem2[125][17] , \mem2[125][16] , \mem2[124][23] ,
         \mem2[124][22] , \mem2[124][21] , \mem2[124][20] , \mem2[124][19] ,
         \mem2[124][18] , \mem2[124][17] , \mem2[124][16] , \mem2[123][23] ,
         \mem2[123][22] , \mem2[123][21] , \mem2[123][20] , \mem2[123][19] ,
         \mem2[123][18] , \mem2[123][17] , \mem2[123][16] , \mem2[122][23] ,
         \mem2[122][22] , \mem2[122][21] , \mem2[122][20] , \mem2[122][19] ,
         \mem2[122][18] , \mem2[122][17] , \mem2[122][16] , \mem2[121][23] ,
         \mem2[121][22] , \mem2[121][21] , \mem2[121][20] , \mem2[121][19] ,
         \mem2[121][18] , \mem2[121][17] , \mem2[121][16] , \mem2[120][23] ,
         \mem2[120][22] , \mem2[120][21] , \mem2[120][20] , \mem2[120][19] ,
         \mem2[120][18] , \mem2[120][17] , \mem2[120][16] , \mem2[119][23] ,
         \mem2[119][22] , \mem2[119][21] , \mem2[119][20] , \mem2[119][19] ,
         \mem2[119][18] , \mem2[119][17] , \mem2[119][16] , \mem2[118][23] ,
         \mem2[118][22] , \mem2[118][21] , \mem2[118][20] , \mem2[118][19] ,
         \mem2[118][18] , \mem2[118][17] , \mem2[118][16] , \mem2[117][23] ,
         \mem2[117][22] , \mem2[117][21] , \mem2[117][20] , \mem2[117][19] ,
         \mem2[117][18] , \mem2[117][17] , \mem2[117][16] , \mem2[116][23] ,
         \mem2[116][22] , \mem2[116][21] , \mem2[116][20] , \mem2[116][19] ,
         \mem2[116][18] , \mem2[116][17] , \mem2[116][16] , \mem2[115][23] ,
         \mem2[115][22] , \mem2[115][21] , \mem2[115][20] , \mem2[115][19] ,
         \mem2[115][18] , \mem2[115][17] , \mem2[115][16] , \mem2[114][23] ,
         \mem2[114][22] , \mem2[114][21] , \mem2[114][20] , \mem2[114][19] ,
         \mem2[114][18] , \mem2[114][17] , \mem2[114][16] , \mem2[113][23] ,
         \mem2[113][22] , \mem2[113][21] , \mem2[113][20] , \mem2[113][19] ,
         \mem2[113][18] , \mem2[113][17] , \mem2[113][16] , \mem2[112][23] ,
         \mem2[112][22] , \mem2[112][21] , \mem2[112][20] , \mem2[112][19] ,
         \mem2[112][18] , \mem2[112][17] , \mem2[112][16] , \mem2[111][23] ,
         \mem2[111][22] , \mem2[111][21] , \mem2[111][20] , \mem2[111][19] ,
         \mem2[111][18] , \mem2[111][17] , \mem2[111][16] , \mem2[110][23] ,
         \mem2[110][22] , \mem2[110][21] , \mem2[110][20] , \mem2[110][19] ,
         \mem2[110][18] , \mem2[110][17] , \mem2[110][16] , \mem2[109][23] ,
         \mem2[109][22] , \mem2[109][21] , \mem2[109][20] , \mem2[109][19] ,
         \mem2[109][18] , \mem2[109][17] , \mem2[109][16] , \mem2[108][23] ,
         \mem2[108][22] , \mem2[108][21] , \mem2[108][20] , \mem2[108][19] ,
         \mem2[108][18] , \mem2[108][17] , \mem2[108][16] , \mem2[107][23] ,
         \mem2[107][22] , \mem2[107][21] , \mem2[107][20] , \mem2[107][19] ,
         \mem2[107][18] , \mem2[107][17] , \mem2[107][16] , \mem2[106][23] ,
         \mem2[106][22] , \mem2[106][21] , \mem2[106][20] , \mem2[106][19] ,
         \mem2[106][18] , \mem2[106][17] , \mem2[106][16] , \mem2[105][23] ,
         \mem2[105][22] , \mem2[105][21] , \mem2[105][20] , \mem2[105][19] ,
         \mem2[105][18] , \mem2[105][17] , \mem2[105][16] , \mem2[104][23] ,
         \mem2[104][22] , \mem2[104][21] , \mem2[104][20] , \mem2[104][19] ,
         \mem2[104][18] , \mem2[104][17] , \mem2[104][16] , \mem2[103][23] ,
         \mem2[103][22] , \mem2[103][21] , \mem2[103][20] , \mem2[103][19] ,
         \mem2[103][18] , \mem2[103][17] , \mem2[103][16] , \mem2[102][23] ,
         \mem2[102][22] , \mem2[102][21] , \mem2[102][20] , \mem2[102][19] ,
         \mem2[102][18] , \mem2[102][17] , \mem2[102][16] , \mem2[101][23] ,
         \mem2[101][22] , \mem2[101][21] , \mem2[101][20] , \mem2[101][19] ,
         \mem2[101][18] , \mem2[101][17] , \mem2[101][16] , \mem2[100][23] ,
         \mem2[100][22] , \mem2[100][21] , \mem2[100][20] , \mem2[100][19] ,
         \mem2[100][18] , \mem2[100][17] , \mem2[100][16] , \mem2[99][23] ,
         \mem2[99][22] , \mem2[99][21] , \mem2[99][20] , \mem2[99][19] ,
         \mem2[99][18] , \mem2[99][17] , \mem2[99][16] , \mem2[98][23] ,
         \mem2[98][22] , \mem2[98][21] , \mem2[98][20] , \mem2[98][19] ,
         \mem2[98][18] , \mem2[98][17] , \mem2[98][16] , \mem2[97][23] ,
         \mem2[97][22] , \mem2[97][21] , \mem2[97][20] , \mem2[97][19] ,
         \mem2[97][18] , \mem2[97][17] , \mem2[97][16] , \mem2[96][23] ,
         \mem2[96][22] , \mem2[96][21] , \mem2[96][20] , \mem2[96][19] ,
         \mem2[96][18] , \mem2[96][17] , \mem2[96][16] , \mem2[95][23] ,
         \mem2[95][22] , \mem2[95][21] , \mem2[95][20] , \mem2[95][19] ,
         \mem2[95][18] , \mem2[95][17] , \mem2[95][16] , \mem2[94][23] ,
         \mem2[94][22] , \mem2[94][21] , \mem2[94][20] , \mem2[94][19] ,
         \mem2[94][18] , \mem2[94][17] , \mem2[94][16] , \mem2[93][23] ,
         \mem2[93][22] , \mem2[93][21] , \mem2[93][20] , \mem2[93][19] ,
         \mem2[93][18] , \mem2[93][17] , \mem2[93][16] , \mem2[92][23] ,
         \mem2[92][22] , \mem2[92][21] , \mem2[92][20] , \mem2[92][19] ,
         \mem2[92][18] , \mem2[92][17] , \mem2[92][16] , \mem2[91][23] ,
         \mem2[91][22] , \mem2[91][21] , \mem2[91][20] , \mem2[91][19] ,
         \mem2[91][18] , \mem2[91][17] , \mem2[91][16] , \mem2[90][23] ,
         \mem2[90][22] , \mem2[90][21] , \mem2[90][20] , \mem2[90][19] ,
         \mem2[90][18] , \mem2[90][17] , \mem2[90][16] , \mem2[89][23] ,
         \mem2[89][22] , \mem2[89][21] , \mem2[89][20] , \mem2[89][19] ,
         \mem2[89][18] , \mem2[89][17] , \mem2[89][16] , \mem2[88][23] ,
         \mem2[88][22] , \mem2[88][21] , \mem2[88][20] , \mem2[88][19] ,
         \mem2[88][18] , \mem2[88][17] , \mem2[88][16] , \mem2[87][23] ,
         \mem2[87][22] , \mem2[87][21] , \mem2[87][20] , \mem2[87][19] ,
         \mem2[87][18] , \mem2[87][17] , \mem2[87][16] , \mem2[86][23] ,
         \mem2[86][22] , \mem2[86][21] , \mem2[86][20] , \mem2[86][19] ,
         \mem2[86][18] , \mem2[86][17] , \mem2[86][16] , \mem2[85][23] ,
         \mem2[85][22] , \mem2[85][21] , \mem2[85][20] , \mem2[85][19] ,
         \mem2[85][18] , \mem2[85][17] , \mem2[85][16] , \mem2[84][23] ,
         \mem2[84][22] , \mem2[84][21] , \mem2[84][20] , \mem2[84][19] ,
         \mem2[84][18] , \mem2[84][17] , \mem2[84][16] , \mem2[83][23] ,
         \mem2[83][22] , \mem2[83][21] , \mem2[83][20] , \mem2[83][19] ,
         \mem2[83][18] , \mem2[83][17] , \mem2[83][16] , \mem2[82][23] ,
         \mem2[82][22] , \mem2[82][21] , \mem2[82][20] , \mem2[82][19] ,
         \mem2[82][18] , \mem2[82][17] , \mem2[82][16] , \mem2[81][23] ,
         \mem2[81][22] , \mem2[81][21] , \mem2[81][20] , \mem2[81][19] ,
         \mem2[81][18] , \mem2[81][17] , \mem2[81][16] , \mem2[80][23] ,
         \mem2[80][22] , \mem2[80][21] , \mem2[80][20] , \mem2[80][19] ,
         \mem2[80][18] , \mem2[80][17] , \mem2[80][16] , \mem2[79][23] ,
         \mem2[79][22] , \mem2[79][21] , \mem2[79][20] , \mem2[79][19] ,
         \mem2[79][18] , \mem2[79][17] , \mem2[79][16] , \mem2[78][23] ,
         \mem2[78][22] , \mem2[78][21] , \mem2[78][20] , \mem2[78][19] ,
         \mem2[78][18] , \mem2[78][17] , \mem2[78][16] , \mem2[77][23] ,
         \mem2[77][22] , \mem2[77][21] , \mem2[77][20] , \mem2[77][19] ,
         \mem2[77][18] , \mem2[77][17] , \mem2[77][16] , \mem2[76][23] ,
         \mem2[76][22] , \mem2[76][21] , \mem2[76][20] , \mem2[76][19] ,
         \mem2[76][18] , \mem2[76][17] , \mem2[76][16] , \mem2[75][23] ,
         \mem2[75][22] , \mem2[75][21] , \mem2[75][20] , \mem2[75][19] ,
         \mem2[75][18] , \mem2[75][17] , \mem2[75][16] , \mem2[74][23] ,
         \mem2[74][22] , \mem2[74][21] , \mem2[74][20] , \mem2[74][19] ,
         \mem2[74][18] , \mem2[74][17] , \mem2[74][16] , \mem2[73][23] ,
         \mem2[73][22] , \mem2[73][21] , \mem2[73][20] , \mem2[73][19] ,
         \mem2[73][18] , \mem2[73][17] , \mem2[73][16] , \mem2[72][23] ,
         \mem2[72][22] , \mem2[72][21] , \mem2[72][20] , \mem2[72][19] ,
         \mem2[72][18] , \mem2[72][17] , \mem2[72][16] , \mem2[71][23] ,
         \mem2[71][22] , \mem2[71][21] , \mem2[71][20] , \mem2[71][19] ,
         \mem2[71][18] , \mem2[71][17] , \mem2[71][16] , \mem2[70][23] ,
         \mem2[70][22] , \mem2[70][21] , \mem2[70][20] , \mem2[70][19] ,
         \mem2[70][18] , \mem2[70][17] , \mem2[70][16] , \mem2[69][23] ,
         \mem2[69][22] , \mem2[69][21] , \mem2[69][20] , \mem2[69][19] ,
         \mem2[69][18] , \mem2[69][17] , \mem2[69][16] , \mem2[68][23] ,
         \mem2[68][22] , \mem2[68][21] , \mem2[68][20] , \mem2[68][19] ,
         \mem2[68][18] , \mem2[68][17] , \mem2[68][16] , \mem2[67][23] ,
         \mem2[67][22] , \mem2[67][21] , \mem2[67][20] , \mem2[67][19] ,
         \mem2[67][18] , \mem2[67][17] , \mem2[67][16] , \mem2[66][23] ,
         \mem2[66][22] , \mem2[66][21] , \mem2[66][20] , \mem2[66][19] ,
         \mem2[66][18] , \mem2[66][17] , \mem2[66][16] , \mem2[65][23] ,
         \mem2[65][22] , \mem2[65][21] , \mem2[65][20] , \mem2[65][19] ,
         \mem2[65][18] , \mem2[65][17] , \mem2[65][16] , \mem2[64][23] ,
         \mem2[64][22] , \mem2[64][21] , \mem2[64][20] , \mem2[64][19] ,
         \mem2[64][18] , \mem2[64][17] , \mem2[64][16] , \mem2[63][23] ,
         \mem2[63][22] , \mem2[63][21] , \mem2[63][20] , \mem2[63][19] ,
         \mem2[63][18] , \mem2[63][17] , \mem2[63][16] , \mem2[62][23] ,
         \mem2[62][22] , \mem2[62][21] , \mem2[62][20] , \mem2[62][19] ,
         \mem2[62][18] , \mem2[62][17] , \mem2[62][16] , \mem2[61][23] ,
         \mem2[61][22] , \mem2[61][21] , \mem2[61][20] , \mem2[61][19] ,
         \mem2[61][18] , \mem2[61][17] , \mem2[61][16] , \mem2[60][23] ,
         \mem2[60][22] , \mem2[60][21] , \mem2[60][20] , \mem2[60][19] ,
         \mem2[60][18] , \mem2[60][17] , \mem2[60][16] , \mem2[59][23] ,
         \mem2[59][22] , \mem2[59][21] , \mem2[59][20] , \mem2[59][19] ,
         \mem2[59][18] , \mem2[59][17] , \mem2[59][16] , \mem2[58][23] ,
         \mem2[58][22] , \mem2[58][21] , \mem2[58][20] , \mem2[58][19] ,
         \mem2[58][18] , \mem2[58][17] , \mem2[58][16] , \mem2[57][23] ,
         \mem2[57][22] , \mem2[57][21] , \mem2[57][20] , \mem2[57][19] ,
         \mem2[57][18] , \mem2[57][17] , \mem2[57][16] , \mem2[56][23] ,
         \mem2[56][22] , \mem2[56][21] , \mem2[56][20] , \mem2[56][19] ,
         \mem2[56][18] , \mem2[56][17] , \mem2[56][16] , \mem2[55][23] ,
         \mem2[55][22] , \mem2[55][21] , \mem2[55][20] , \mem2[55][19] ,
         \mem2[55][18] , \mem2[55][17] , \mem2[55][16] , \mem2[54][23] ,
         \mem2[54][22] , \mem2[54][21] , \mem2[54][20] , \mem2[54][19] ,
         \mem2[54][18] , \mem2[54][17] , \mem2[54][16] , \mem2[53][23] ,
         \mem2[53][22] , \mem2[53][21] , \mem2[53][20] , \mem2[53][19] ,
         \mem2[53][18] , \mem2[53][17] , \mem2[53][16] , \mem2[52][23] ,
         \mem2[52][22] , \mem2[52][21] , \mem2[52][20] , \mem2[52][19] ,
         \mem2[52][18] , \mem2[52][17] , \mem2[52][16] , \mem2[51][23] ,
         \mem2[51][22] , \mem2[51][21] , \mem2[51][20] , \mem2[51][19] ,
         \mem2[51][18] , \mem2[51][17] , \mem2[51][16] , \mem2[50][23] ,
         \mem2[50][22] , \mem2[50][21] , \mem2[50][20] , \mem2[50][19] ,
         \mem2[50][18] , \mem2[50][17] , \mem2[50][16] , \mem2[49][23] ,
         \mem2[49][22] , \mem2[49][21] , \mem2[49][20] , \mem2[49][19] ,
         \mem2[49][18] , \mem2[49][17] , \mem2[49][16] , \mem2[48][23] ,
         \mem2[48][22] , \mem2[48][21] , \mem2[48][20] , \mem2[48][19] ,
         \mem2[48][18] , \mem2[48][17] , \mem2[48][16] , \mem2[47][23] ,
         \mem2[47][22] , \mem2[47][21] , \mem2[47][20] , \mem2[47][19] ,
         \mem2[47][18] , \mem2[47][17] , \mem2[47][16] , \mem2[46][23] ,
         \mem2[46][22] , \mem2[46][21] , \mem2[46][20] , \mem2[46][19] ,
         \mem2[46][18] , \mem2[46][17] , \mem2[46][16] , \mem2[45][23] ,
         \mem2[45][22] , \mem2[45][21] , \mem2[45][20] , \mem2[45][19] ,
         \mem2[45][18] , \mem2[45][17] , \mem2[45][16] , \mem2[44][23] ,
         \mem2[44][22] , \mem2[44][21] , \mem2[44][20] , \mem2[44][19] ,
         \mem2[44][18] , \mem2[44][17] , \mem2[44][16] , \mem2[43][23] ,
         \mem2[43][22] , \mem2[43][21] , \mem2[43][20] , \mem2[43][19] ,
         \mem2[43][18] , \mem2[43][17] , \mem2[43][16] , \mem2[42][23] ,
         \mem2[42][22] , \mem2[42][21] , \mem2[42][20] , \mem2[42][19] ,
         \mem2[42][18] , \mem2[42][17] , \mem2[42][16] , \mem2[41][23] ,
         \mem2[41][22] , \mem2[41][21] , \mem2[41][20] , \mem2[41][19] ,
         \mem2[41][18] , \mem2[41][17] , \mem2[41][16] , \mem2[40][23] ,
         \mem2[40][22] , \mem2[40][21] , \mem2[40][20] , \mem2[40][19] ,
         \mem2[40][18] , \mem2[40][17] , \mem2[40][16] , \mem2[39][23] ,
         \mem2[39][22] , \mem2[39][21] , \mem2[39][20] , \mem2[39][19] ,
         \mem2[39][18] , \mem2[39][17] , \mem2[39][16] , \mem2[38][23] ,
         \mem2[38][22] , \mem2[38][21] , \mem2[38][20] , \mem2[38][19] ,
         \mem2[38][18] , \mem2[38][17] , \mem2[38][16] , \mem2[37][23] ,
         \mem2[37][22] , \mem2[37][21] , \mem2[37][20] , \mem2[37][19] ,
         \mem2[37][18] , \mem2[37][17] , \mem2[37][16] , \mem2[36][23] ,
         \mem2[36][22] , \mem2[36][21] , \mem2[36][20] , \mem2[36][19] ,
         \mem2[36][18] , \mem2[36][17] , \mem2[36][16] , \mem2[35][23] ,
         \mem2[35][22] , \mem2[35][21] , \mem2[35][20] , \mem2[35][19] ,
         \mem2[35][18] , \mem2[35][17] , \mem2[35][16] , \mem2[34][23] ,
         \mem2[34][22] , \mem2[34][21] , \mem2[34][20] , \mem2[34][19] ,
         \mem2[34][18] , \mem2[34][17] , \mem2[34][16] , \mem2[33][23] ,
         \mem2[33][22] , \mem2[33][21] , \mem2[33][20] , \mem2[33][19] ,
         \mem2[33][18] , \mem2[33][17] , \mem2[33][16] , \mem2[32][23] ,
         \mem2[32][22] , \mem2[32][21] , \mem2[32][20] , \mem2[32][19] ,
         \mem2[32][18] , \mem2[32][17] , \mem2[32][16] , \mem2[31][23] ,
         \mem2[31][22] , \mem2[31][21] , \mem2[31][20] , \mem2[31][19] ,
         \mem2[31][18] , \mem2[31][17] , \mem2[31][16] , \mem2[30][23] ,
         \mem2[30][22] , \mem2[30][21] , \mem2[30][20] , \mem2[30][19] ,
         \mem2[30][18] , \mem2[30][17] , \mem2[30][16] , \mem2[29][23] ,
         \mem2[29][22] , \mem2[29][21] , \mem2[29][20] , \mem2[29][19] ,
         \mem2[29][18] , \mem2[29][17] , \mem2[29][16] , \mem2[28][23] ,
         \mem2[28][22] , \mem2[28][21] , \mem2[28][20] , \mem2[28][19] ,
         \mem2[28][18] , \mem2[28][17] , \mem2[28][16] , \mem2[27][23] ,
         \mem2[27][22] , \mem2[27][21] , \mem2[27][20] , \mem2[27][19] ,
         \mem2[27][18] , \mem2[27][17] , \mem2[27][16] , \mem2[26][23] ,
         \mem2[26][22] , \mem2[26][21] , \mem2[26][20] , \mem2[26][19] ,
         \mem2[26][18] , \mem2[26][17] , \mem2[26][16] , \mem2[25][23] ,
         \mem2[25][22] , \mem2[25][21] , \mem2[25][20] , \mem2[25][19] ,
         \mem2[25][18] , \mem2[25][17] , \mem2[25][16] , \mem2[24][23] ,
         \mem2[24][22] , \mem2[24][21] , \mem2[24][20] , \mem2[24][19] ,
         \mem2[24][18] , \mem2[24][17] , \mem2[24][16] , \mem2[23][23] ,
         \mem2[23][22] , \mem2[23][21] , \mem2[23][20] , \mem2[23][19] ,
         \mem2[23][18] , \mem2[23][17] , \mem2[23][16] , \mem2[22][23] ,
         \mem2[22][22] , \mem2[22][21] , \mem2[22][20] , \mem2[22][19] ,
         \mem2[22][18] , \mem2[22][17] , \mem2[22][16] , \mem2[21][23] ,
         \mem2[21][22] , \mem2[21][21] , \mem2[21][20] , \mem2[21][19] ,
         \mem2[21][18] , \mem2[21][17] , \mem2[21][16] , \mem2[20][23] ,
         \mem2[20][22] , \mem2[20][21] , \mem2[20][20] , \mem2[20][19] ,
         \mem2[20][18] , \mem2[20][17] , \mem2[20][16] , \mem2[19][23] ,
         \mem2[19][22] , \mem2[19][21] , \mem2[19][20] , \mem2[19][19] ,
         \mem2[19][18] , \mem2[19][17] , \mem2[19][16] , \mem2[18][23] ,
         \mem2[18][22] , \mem2[18][21] , \mem2[18][20] , \mem2[18][19] ,
         \mem2[18][18] , \mem2[18][17] , \mem2[18][16] , \mem2[17][23] ,
         \mem2[17][22] , \mem2[17][21] , \mem2[17][20] , \mem2[17][19] ,
         \mem2[17][18] , \mem2[17][17] , \mem2[17][16] , \mem2[16][23] ,
         \mem2[16][22] , \mem2[16][21] , \mem2[16][20] , \mem2[16][19] ,
         \mem2[16][18] , \mem2[16][17] , \mem2[16][16] , \mem2[15][23] ,
         \mem2[15][22] , \mem2[15][21] , \mem2[15][20] , \mem2[15][19] ,
         \mem2[15][18] , \mem2[15][17] , \mem2[15][16] , \mem2[14][23] ,
         \mem2[14][22] , \mem2[14][21] , \mem2[14][20] , \mem2[14][19] ,
         \mem2[14][18] , \mem2[14][17] , \mem2[14][16] , \mem2[13][23] ,
         \mem2[13][22] , \mem2[13][21] , \mem2[13][20] , \mem2[13][19] ,
         \mem2[13][18] , \mem2[13][17] , \mem2[13][16] , \mem2[12][23] ,
         \mem2[12][22] , \mem2[12][21] , \mem2[12][20] , \mem2[12][19] ,
         \mem2[12][18] , \mem2[12][17] , \mem2[12][16] , \mem2[11][23] ,
         \mem2[11][22] , \mem2[11][21] , \mem2[11][20] , \mem2[11][19] ,
         \mem2[11][18] , \mem2[11][17] , \mem2[11][16] , \mem2[10][23] ,
         \mem2[10][22] , \mem2[10][21] , \mem2[10][20] , \mem2[10][19] ,
         \mem2[10][18] , \mem2[10][17] , \mem2[10][16] , \mem2[9][23] ,
         \mem2[9][22] , \mem2[9][21] , \mem2[9][20] , \mem2[9][19] ,
         \mem2[9][18] , \mem2[9][17] , \mem2[9][16] , \mem2[8][23] ,
         \mem2[8][22] , \mem2[8][21] , \mem2[8][20] , \mem2[8][19] ,
         \mem2[8][18] , \mem2[8][17] , \mem2[8][16] , \mem2[7][23] ,
         \mem2[7][22] , \mem2[7][21] , \mem2[7][20] , \mem2[7][19] ,
         \mem2[7][18] , \mem2[7][17] , \mem2[7][16] , \mem2[6][23] ,
         \mem2[6][22] , \mem2[6][21] , \mem2[6][20] , \mem2[6][19] ,
         \mem2[6][18] , \mem2[6][17] , \mem2[6][16] , \mem2[5][23] ,
         \mem2[5][22] , \mem2[5][21] , \mem2[5][20] , \mem2[5][19] ,
         \mem2[5][18] , \mem2[5][17] , \mem2[5][16] , \mem2[4][23] ,
         \mem2[4][22] , \mem2[4][21] , \mem2[4][20] , \mem2[4][19] ,
         \mem2[4][18] , \mem2[4][17] , \mem2[4][16] , \mem2[3][23] ,
         \mem2[3][22] , \mem2[3][21] , \mem2[3][20] , \mem2[3][19] ,
         \mem2[3][18] , \mem2[3][17] , \mem2[3][16] , \mem2[2][23] ,
         \mem2[2][22] , \mem2[2][21] , \mem2[2][20] , \mem2[2][19] ,
         \mem2[2][18] , \mem2[2][17] , \mem2[2][16] , \mem2[1][23] ,
         \mem2[1][22] , \mem2[1][21] , \mem2[1][20] , \mem2[1][19] ,
         \mem2[1][18] , \mem2[1][17] , \mem2[1][16] , \mem2[0][23] ,
         \mem2[0][22] , \mem2[0][21] , \mem2[0][20] , \mem2[0][19] ,
         \mem2[0][18] , \mem2[0][17] , \mem2[0][16] , \mem1[255][15] ,
         \mem1[255][14] , \mem1[255][13] , \mem1[255][12] , \mem1[255][11] ,
         \mem1[255][10] , \mem1[255][9] , \mem1[255][8] , \mem1[254][15] ,
         \mem1[254][14] , \mem1[254][13] , \mem1[254][12] , \mem1[254][11] ,
         \mem1[254][10] , \mem1[254][9] , \mem1[254][8] , \mem1[253][15] ,
         \mem1[253][14] , \mem1[253][13] , \mem1[253][12] , \mem1[253][11] ,
         \mem1[253][10] , \mem1[253][9] , \mem1[253][8] , \mem1[252][15] ,
         \mem1[252][14] , \mem1[252][13] , \mem1[252][12] , \mem1[252][11] ,
         \mem1[252][10] , \mem1[252][9] , \mem1[252][8] , \mem1[251][15] ,
         \mem1[251][14] , \mem1[251][13] , \mem1[251][12] , \mem1[251][11] ,
         \mem1[251][10] , \mem1[251][9] , \mem1[251][8] , \mem1[250][15] ,
         \mem1[250][14] , \mem1[250][13] , \mem1[250][12] , \mem1[250][11] ,
         \mem1[250][10] , \mem1[250][9] , \mem1[250][8] , \mem1[249][15] ,
         \mem1[249][14] , \mem1[249][13] , \mem1[249][12] , \mem1[249][11] ,
         \mem1[249][10] , \mem1[249][9] , \mem1[249][8] , \mem1[248][15] ,
         \mem1[248][14] , \mem1[248][13] , \mem1[248][12] , \mem1[248][11] ,
         \mem1[248][10] , \mem1[248][9] , \mem1[248][8] , \mem1[247][15] ,
         \mem1[247][14] , \mem1[247][13] , \mem1[247][12] , \mem1[247][11] ,
         \mem1[247][10] , \mem1[247][9] , \mem1[247][8] , \mem1[246][15] ,
         \mem1[246][14] , \mem1[246][13] , \mem1[246][12] , \mem1[246][11] ,
         \mem1[246][10] , \mem1[246][9] , \mem1[246][8] , \mem1[245][15] ,
         \mem1[245][14] , \mem1[245][13] , \mem1[245][12] , \mem1[245][11] ,
         \mem1[245][10] , \mem1[245][9] , \mem1[245][8] , \mem1[244][15] ,
         \mem1[244][14] , \mem1[244][13] , \mem1[244][12] , \mem1[244][11] ,
         \mem1[244][10] , \mem1[244][9] , \mem1[244][8] , \mem1[243][15] ,
         \mem1[243][14] , \mem1[243][13] , \mem1[243][12] , \mem1[243][11] ,
         \mem1[243][10] , \mem1[243][9] , \mem1[243][8] , \mem1[242][15] ,
         \mem1[242][14] , \mem1[242][13] , \mem1[242][12] , \mem1[242][11] ,
         \mem1[242][10] , \mem1[242][9] , \mem1[242][8] , \mem1[241][15] ,
         \mem1[241][14] , \mem1[241][13] , \mem1[241][12] , \mem1[241][11] ,
         \mem1[241][10] , \mem1[241][9] , \mem1[241][8] , \mem1[240][15] ,
         \mem1[240][14] , \mem1[240][13] , \mem1[240][12] , \mem1[240][11] ,
         \mem1[240][10] , \mem1[240][9] , \mem1[240][8] , \mem1[239][15] ,
         \mem1[239][14] , \mem1[239][13] , \mem1[239][12] , \mem1[239][11] ,
         \mem1[239][10] , \mem1[239][9] , \mem1[239][8] , \mem1[238][15] ,
         \mem1[238][14] , \mem1[238][13] , \mem1[238][12] , \mem1[238][11] ,
         \mem1[238][10] , \mem1[238][9] , \mem1[238][8] , \mem1[237][15] ,
         \mem1[237][14] , \mem1[237][13] , \mem1[237][12] , \mem1[237][11] ,
         \mem1[237][10] , \mem1[237][9] , \mem1[237][8] , \mem1[236][15] ,
         \mem1[236][14] , \mem1[236][13] , \mem1[236][12] , \mem1[236][11] ,
         \mem1[236][10] , \mem1[236][9] , \mem1[236][8] , \mem1[235][15] ,
         \mem1[235][14] , \mem1[235][13] , \mem1[235][12] , \mem1[235][11] ,
         \mem1[235][10] , \mem1[235][9] , \mem1[235][8] , \mem1[234][15] ,
         \mem1[234][14] , \mem1[234][13] , \mem1[234][12] , \mem1[234][11] ,
         \mem1[234][10] , \mem1[234][9] , \mem1[234][8] , \mem1[233][15] ,
         \mem1[233][14] , \mem1[233][13] , \mem1[233][12] , \mem1[233][11] ,
         \mem1[233][10] , \mem1[233][9] , \mem1[233][8] , \mem1[232][15] ,
         \mem1[232][14] , \mem1[232][13] , \mem1[232][12] , \mem1[232][11] ,
         \mem1[232][10] , \mem1[232][9] , \mem1[232][8] , \mem1[231][15] ,
         \mem1[231][14] , \mem1[231][13] , \mem1[231][12] , \mem1[231][11] ,
         \mem1[231][10] , \mem1[231][9] , \mem1[231][8] , \mem1[230][15] ,
         \mem1[230][14] , \mem1[230][13] , \mem1[230][12] , \mem1[230][11] ,
         \mem1[230][10] , \mem1[230][9] , \mem1[230][8] , \mem1[229][15] ,
         \mem1[229][14] , \mem1[229][13] , \mem1[229][12] , \mem1[229][11] ,
         \mem1[229][10] , \mem1[229][9] , \mem1[229][8] , \mem1[228][15] ,
         \mem1[228][14] , \mem1[228][13] , \mem1[228][12] , \mem1[228][11] ,
         \mem1[228][10] , \mem1[228][9] , \mem1[228][8] , \mem1[227][15] ,
         \mem1[227][14] , \mem1[227][13] , \mem1[227][12] , \mem1[227][11] ,
         \mem1[227][10] , \mem1[227][9] , \mem1[227][8] , \mem1[226][15] ,
         \mem1[226][14] , \mem1[226][13] , \mem1[226][12] , \mem1[226][11] ,
         \mem1[226][10] , \mem1[226][9] , \mem1[226][8] , \mem1[225][15] ,
         \mem1[225][14] , \mem1[225][13] , \mem1[225][12] , \mem1[225][11] ,
         \mem1[225][10] , \mem1[225][9] , \mem1[225][8] , \mem1[224][15] ,
         \mem1[224][14] , \mem1[224][13] , \mem1[224][12] , \mem1[224][11] ,
         \mem1[224][10] , \mem1[224][9] , \mem1[224][8] , \mem1[223][15] ,
         \mem1[223][14] , \mem1[223][13] , \mem1[223][12] , \mem1[223][11] ,
         \mem1[223][10] , \mem1[223][9] , \mem1[223][8] , \mem1[222][15] ,
         \mem1[222][14] , \mem1[222][13] , \mem1[222][12] , \mem1[222][11] ,
         \mem1[222][10] , \mem1[222][9] , \mem1[222][8] , \mem1[221][15] ,
         \mem1[221][14] , \mem1[221][13] , \mem1[221][12] , \mem1[221][11] ,
         \mem1[221][10] , \mem1[221][9] , \mem1[221][8] , \mem1[220][15] ,
         \mem1[220][14] , \mem1[220][13] , \mem1[220][12] , \mem1[220][11] ,
         \mem1[220][10] , \mem1[220][9] , \mem1[220][8] , \mem1[219][15] ,
         \mem1[219][14] , \mem1[219][13] , \mem1[219][12] , \mem1[219][11] ,
         \mem1[219][10] , \mem1[219][9] , \mem1[219][8] , \mem1[218][15] ,
         \mem1[218][14] , \mem1[218][13] , \mem1[218][12] , \mem1[218][11] ,
         \mem1[218][10] , \mem1[218][9] , \mem1[218][8] , \mem1[217][15] ,
         \mem1[217][14] , \mem1[217][13] , \mem1[217][12] , \mem1[217][11] ,
         \mem1[217][10] , \mem1[217][9] , \mem1[217][8] , \mem1[216][15] ,
         \mem1[216][14] , \mem1[216][13] , \mem1[216][12] , \mem1[216][11] ,
         \mem1[216][10] , \mem1[216][9] , \mem1[216][8] , \mem1[215][15] ,
         \mem1[215][14] , \mem1[215][13] , \mem1[215][12] , \mem1[215][11] ,
         \mem1[215][10] , \mem1[215][9] , \mem1[215][8] , \mem1[214][15] ,
         \mem1[214][14] , \mem1[214][13] , \mem1[214][12] , \mem1[214][11] ,
         \mem1[214][10] , \mem1[214][9] , \mem1[214][8] , \mem1[213][15] ,
         \mem1[213][14] , \mem1[213][13] , \mem1[213][12] , \mem1[213][11] ,
         \mem1[213][10] , \mem1[213][9] , \mem1[213][8] , \mem1[212][15] ,
         \mem1[212][14] , \mem1[212][13] , \mem1[212][12] , \mem1[212][11] ,
         \mem1[212][10] , \mem1[212][9] , \mem1[212][8] , \mem1[211][15] ,
         \mem1[211][14] , \mem1[211][13] , \mem1[211][12] , \mem1[211][11] ,
         \mem1[211][10] , \mem1[211][9] , \mem1[211][8] , \mem1[210][15] ,
         \mem1[210][14] , \mem1[210][13] , \mem1[210][12] , \mem1[210][11] ,
         \mem1[210][10] , \mem1[210][9] , \mem1[210][8] , \mem1[209][15] ,
         \mem1[209][14] , \mem1[209][13] , \mem1[209][12] , \mem1[209][11] ,
         \mem1[209][10] , \mem1[209][9] , \mem1[209][8] , \mem1[208][15] ,
         \mem1[208][14] , \mem1[208][13] , \mem1[208][12] , \mem1[208][11] ,
         \mem1[208][10] , \mem1[208][9] , \mem1[208][8] , \mem1[207][15] ,
         \mem1[207][14] , \mem1[207][13] , \mem1[207][12] , \mem1[207][11] ,
         \mem1[207][10] , \mem1[207][9] , \mem1[207][8] , \mem1[206][15] ,
         \mem1[206][14] , \mem1[206][13] , \mem1[206][12] , \mem1[206][11] ,
         \mem1[206][10] , \mem1[206][9] , \mem1[206][8] , \mem1[205][15] ,
         \mem1[205][14] , \mem1[205][13] , \mem1[205][12] , \mem1[205][11] ,
         \mem1[205][10] , \mem1[205][9] , \mem1[205][8] , \mem1[204][15] ,
         \mem1[204][14] , \mem1[204][13] , \mem1[204][12] , \mem1[204][11] ,
         \mem1[204][10] , \mem1[204][9] , \mem1[204][8] , \mem1[203][15] ,
         \mem1[203][14] , \mem1[203][13] , \mem1[203][12] , \mem1[203][11] ,
         \mem1[203][10] , \mem1[203][9] , \mem1[203][8] , \mem1[202][15] ,
         \mem1[202][14] , \mem1[202][13] , \mem1[202][12] , \mem1[202][11] ,
         \mem1[202][10] , \mem1[202][9] , \mem1[202][8] , \mem1[201][15] ,
         \mem1[201][14] , \mem1[201][13] , \mem1[201][12] , \mem1[201][11] ,
         \mem1[201][10] , \mem1[201][9] , \mem1[201][8] , \mem1[200][15] ,
         \mem1[200][14] , \mem1[200][13] , \mem1[200][12] , \mem1[200][11] ,
         \mem1[200][10] , \mem1[200][9] , \mem1[200][8] , \mem1[199][15] ,
         \mem1[199][14] , \mem1[199][13] , \mem1[199][12] , \mem1[199][11] ,
         \mem1[199][10] , \mem1[199][9] , \mem1[199][8] , \mem1[198][15] ,
         \mem1[198][14] , \mem1[198][13] , \mem1[198][12] , \mem1[198][11] ,
         \mem1[198][10] , \mem1[198][9] , \mem1[198][8] , \mem1[197][15] ,
         \mem1[197][14] , \mem1[197][13] , \mem1[197][12] , \mem1[197][11] ,
         \mem1[197][10] , \mem1[197][9] , \mem1[197][8] , \mem1[196][15] ,
         \mem1[196][14] , \mem1[196][13] , \mem1[196][12] , \mem1[196][11] ,
         \mem1[196][10] , \mem1[196][9] , \mem1[196][8] , \mem1[195][15] ,
         \mem1[195][14] , \mem1[195][13] , \mem1[195][12] , \mem1[195][11] ,
         \mem1[195][10] , \mem1[195][9] , \mem1[195][8] , \mem1[194][15] ,
         \mem1[194][14] , \mem1[194][13] , \mem1[194][12] , \mem1[194][11] ,
         \mem1[194][10] , \mem1[194][9] , \mem1[194][8] , \mem1[193][15] ,
         \mem1[193][14] , \mem1[193][13] , \mem1[193][12] , \mem1[193][11] ,
         \mem1[193][10] , \mem1[193][9] , \mem1[193][8] , \mem1[192][15] ,
         \mem1[192][14] , \mem1[192][13] , \mem1[192][12] , \mem1[192][11] ,
         \mem1[192][10] , \mem1[192][9] , \mem1[192][8] , \mem1[191][15] ,
         \mem1[191][14] , \mem1[191][13] , \mem1[191][12] , \mem1[191][11] ,
         \mem1[191][10] , \mem1[191][9] , \mem1[191][8] , \mem1[190][15] ,
         \mem1[190][14] , \mem1[190][13] , \mem1[190][12] , \mem1[190][11] ,
         \mem1[190][10] , \mem1[190][9] , \mem1[190][8] , \mem1[189][15] ,
         \mem1[189][14] , \mem1[189][13] , \mem1[189][12] , \mem1[189][11] ,
         \mem1[189][10] , \mem1[189][9] , \mem1[189][8] , \mem1[188][15] ,
         \mem1[188][14] , \mem1[188][13] , \mem1[188][12] , \mem1[188][11] ,
         \mem1[188][10] , \mem1[188][9] , \mem1[188][8] , \mem1[187][15] ,
         \mem1[187][14] , \mem1[187][13] , \mem1[187][12] , \mem1[187][11] ,
         \mem1[187][10] , \mem1[187][9] , \mem1[187][8] , \mem1[186][15] ,
         \mem1[186][14] , \mem1[186][13] , \mem1[186][12] , \mem1[186][11] ,
         \mem1[186][10] , \mem1[186][9] , \mem1[186][8] , \mem1[185][15] ,
         \mem1[185][14] , \mem1[185][13] , \mem1[185][12] , \mem1[185][11] ,
         \mem1[185][10] , \mem1[185][9] , \mem1[185][8] , \mem1[184][15] ,
         \mem1[184][14] , \mem1[184][13] , \mem1[184][12] , \mem1[184][11] ,
         \mem1[184][10] , \mem1[184][9] , \mem1[184][8] , \mem1[183][15] ,
         \mem1[183][14] , \mem1[183][13] , \mem1[183][12] , \mem1[183][11] ,
         \mem1[183][10] , \mem1[183][9] , \mem1[183][8] , \mem1[182][15] ,
         \mem1[182][14] , \mem1[182][13] , \mem1[182][12] , \mem1[182][11] ,
         \mem1[182][10] , \mem1[182][9] , \mem1[182][8] , \mem1[181][15] ,
         \mem1[181][14] , \mem1[181][13] , \mem1[181][12] , \mem1[181][11] ,
         \mem1[181][10] , \mem1[181][9] , \mem1[181][8] , \mem1[180][15] ,
         \mem1[180][14] , \mem1[180][13] , \mem1[180][12] , \mem1[180][11] ,
         \mem1[180][10] , \mem1[180][9] , \mem1[180][8] , \mem1[179][15] ,
         \mem1[179][14] , \mem1[179][13] , \mem1[179][12] , \mem1[179][11] ,
         \mem1[179][10] , \mem1[179][9] , \mem1[179][8] , \mem1[178][15] ,
         \mem1[178][14] , \mem1[178][13] , \mem1[178][12] , \mem1[178][11] ,
         \mem1[178][10] , \mem1[178][9] , \mem1[178][8] , \mem1[177][15] ,
         \mem1[177][14] , \mem1[177][13] , \mem1[177][12] , \mem1[177][11] ,
         \mem1[177][10] , \mem1[177][9] , \mem1[177][8] , \mem1[176][15] ,
         \mem1[176][14] , \mem1[176][13] , \mem1[176][12] , \mem1[176][11] ,
         \mem1[176][10] , \mem1[176][9] , \mem1[176][8] , \mem1[175][15] ,
         \mem1[175][14] , \mem1[175][13] , \mem1[175][12] , \mem1[175][11] ,
         \mem1[175][10] , \mem1[175][9] , \mem1[175][8] , \mem1[174][15] ,
         \mem1[174][14] , \mem1[174][13] , \mem1[174][12] , \mem1[174][11] ,
         \mem1[174][10] , \mem1[174][9] , \mem1[174][8] , \mem1[173][15] ,
         \mem1[173][14] , \mem1[173][13] , \mem1[173][12] , \mem1[173][11] ,
         \mem1[173][10] , \mem1[173][9] , \mem1[173][8] , \mem1[172][15] ,
         \mem1[172][14] , \mem1[172][13] , \mem1[172][12] , \mem1[172][11] ,
         \mem1[172][10] , \mem1[172][9] , \mem1[172][8] , \mem1[171][15] ,
         \mem1[171][14] , \mem1[171][13] , \mem1[171][12] , \mem1[171][11] ,
         \mem1[171][10] , \mem1[171][9] , \mem1[171][8] , \mem1[170][15] ,
         \mem1[170][14] , \mem1[170][13] , \mem1[170][12] , \mem1[170][11] ,
         \mem1[170][10] , \mem1[170][9] , \mem1[170][8] , \mem1[169][15] ,
         \mem1[169][14] , \mem1[169][13] , \mem1[169][12] , \mem1[169][11] ,
         \mem1[169][10] , \mem1[169][9] , \mem1[169][8] , \mem1[168][15] ,
         \mem1[168][14] , \mem1[168][13] , \mem1[168][12] , \mem1[168][11] ,
         \mem1[168][10] , \mem1[168][9] , \mem1[168][8] , \mem1[167][15] ,
         \mem1[167][14] , \mem1[167][13] , \mem1[167][12] , \mem1[167][11] ,
         \mem1[167][10] , \mem1[167][9] , \mem1[167][8] , \mem1[166][15] ,
         \mem1[166][14] , \mem1[166][13] , \mem1[166][12] , \mem1[166][11] ,
         \mem1[166][10] , \mem1[166][9] , \mem1[166][8] , \mem1[165][15] ,
         \mem1[165][14] , \mem1[165][13] , \mem1[165][12] , \mem1[165][11] ,
         \mem1[165][10] , \mem1[165][9] , \mem1[165][8] , \mem1[164][15] ,
         \mem1[164][14] , \mem1[164][13] , \mem1[164][12] , \mem1[164][11] ,
         \mem1[164][10] , \mem1[164][9] , \mem1[164][8] , \mem1[163][15] ,
         \mem1[163][14] , \mem1[163][13] , \mem1[163][12] , \mem1[163][11] ,
         \mem1[163][10] , \mem1[163][9] , \mem1[163][8] , \mem1[162][15] ,
         \mem1[162][14] , \mem1[162][13] , \mem1[162][12] , \mem1[162][11] ,
         \mem1[162][10] , \mem1[162][9] , \mem1[162][8] , \mem1[161][15] ,
         \mem1[161][14] , \mem1[161][13] , \mem1[161][12] , \mem1[161][11] ,
         \mem1[161][10] , \mem1[161][9] , \mem1[161][8] , \mem1[160][15] ,
         \mem1[160][14] , \mem1[160][13] , \mem1[160][12] , \mem1[160][11] ,
         \mem1[160][10] , \mem1[160][9] , \mem1[160][8] , \mem1[159][15] ,
         \mem1[159][14] , \mem1[159][13] , \mem1[159][12] , \mem1[159][11] ,
         \mem1[159][10] , \mem1[159][9] , \mem1[159][8] , \mem1[158][15] ,
         \mem1[158][14] , \mem1[158][13] , \mem1[158][12] , \mem1[158][11] ,
         \mem1[158][10] , \mem1[158][9] , \mem1[158][8] , \mem1[157][15] ,
         \mem1[157][14] , \mem1[157][13] , \mem1[157][12] , \mem1[157][11] ,
         \mem1[157][10] , \mem1[157][9] , \mem1[157][8] , \mem1[156][15] ,
         \mem1[156][14] , \mem1[156][13] , \mem1[156][12] , \mem1[156][11] ,
         \mem1[156][10] , \mem1[156][9] , \mem1[156][8] , \mem1[155][15] ,
         \mem1[155][14] , \mem1[155][13] , \mem1[155][12] , \mem1[155][11] ,
         \mem1[155][10] , \mem1[155][9] , \mem1[155][8] , \mem1[154][15] ,
         \mem1[154][14] , \mem1[154][13] , \mem1[154][12] , \mem1[154][11] ,
         \mem1[154][10] , \mem1[154][9] , \mem1[154][8] , \mem1[153][15] ,
         \mem1[153][14] , \mem1[153][13] , \mem1[153][12] , \mem1[153][11] ,
         \mem1[153][10] , \mem1[153][9] , \mem1[153][8] , \mem1[152][15] ,
         \mem1[152][14] , \mem1[152][13] , \mem1[152][12] , \mem1[152][11] ,
         \mem1[152][10] , \mem1[152][9] , \mem1[152][8] , \mem1[151][15] ,
         \mem1[151][14] , \mem1[151][13] , \mem1[151][12] , \mem1[151][11] ,
         \mem1[151][10] , \mem1[151][9] , \mem1[151][8] , \mem1[150][15] ,
         \mem1[150][14] , \mem1[150][13] , \mem1[150][12] , \mem1[150][11] ,
         \mem1[150][10] , \mem1[150][9] , \mem1[150][8] , \mem1[149][15] ,
         \mem1[149][14] , \mem1[149][13] , \mem1[149][12] , \mem1[149][11] ,
         \mem1[149][10] , \mem1[149][9] , \mem1[149][8] , \mem1[148][15] ,
         \mem1[148][14] , \mem1[148][13] , \mem1[148][12] , \mem1[148][11] ,
         \mem1[148][10] , \mem1[148][9] , \mem1[148][8] , \mem1[147][15] ,
         \mem1[147][14] , \mem1[147][13] , \mem1[147][12] , \mem1[147][11] ,
         \mem1[147][10] , \mem1[147][9] , \mem1[147][8] , \mem1[146][15] ,
         \mem1[146][14] , \mem1[146][13] , \mem1[146][12] , \mem1[146][11] ,
         \mem1[146][10] , \mem1[146][9] , \mem1[146][8] , \mem1[145][15] ,
         \mem1[145][14] , \mem1[145][13] , \mem1[145][12] , \mem1[145][11] ,
         \mem1[145][10] , \mem1[145][9] , \mem1[145][8] , \mem1[144][15] ,
         \mem1[144][14] , \mem1[144][13] , \mem1[144][12] , \mem1[144][11] ,
         \mem1[144][10] , \mem1[144][9] , \mem1[144][8] , \mem1[143][15] ,
         \mem1[143][14] , \mem1[143][13] , \mem1[143][12] , \mem1[143][11] ,
         \mem1[143][10] , \mem1[143][9] , \mem1[143][8] , \mem1[142][15] ,
         \mem1[142][14] , \mem1[142][13] , \mem1[142][12] , \mem1[142][11] ,
         \mem1[142][10] , \mem1[142][9] , \mem1[142][8] , \mem1[141][15] ,
         \mem1[141][14] , \mem1[141][13] , \mem1[141][12] , \mem1[141][11] ,
         \mem1[141][10] , \mem1[141][9] , \mem1[141][8] , \mem1[140][15] ,
         \mem1[140][14] , \mem1[140][13] , \mem1[140][12] , \mem1[140][11] ,
         \mem1[140][10] , \mem1[140][9] , \mem1[140][8] , \mem1[139][15] ,
         \mem1[139][14] , \mem1[139][13] , \mem1[139][12] , \mem1[139][11] ,
         \mem1[139][10] , \mem1[139][9] , \mem1[139][8] , \mem1[138][15] ,
         \mem1[138][14] , \mem1[138][13] , \mem1[138][12] , \mem1[138][11] ,
         \mem1[138][10] , \mem1[138][9] , \mem1[138][8] , \mem1[137][15] ,
         \mem1[137][14] , \mem1[137][13] , \mem1[137][12] , \mem1[137][11] ,
         \mem1[137][10] , \mem1[137][9] , \mem1[137][8] , \mem1[136][15] ,
         \mem1[136][14] , \mem1[136][13] , \mem1[136][12] , \mem1[136][11] ,
         \mem1[136][10] , \mem1[136][9] , \mem1[136][8] , \mem1[135][15] ,
         \mem1[135][14] , \mem1[135][13] , \mem1[135][12] , \mem1[135][11] ,
         \mem1[135][10] , \mem1[135][9] , \mem1[135][8] , \mem1[134][15] ,
         \mem1[134][14] , \mem1[134][13] , \mem1[134][12] , \mem1[134][11] ,
         \mem1[134][10] , \mem1[134][9] , \mem1[134][8] , \mem1[133][15] ,
         \mem1[133][14] , \mem1[133][13] , \mem1[133][12] , \mem1[133][11] ,
         \mem1[133][10] , \mem1[133][9] , \mem1[133][8] , \mem1[132][15] ,
         \mem1[132][14] , \mem1[132][13] , \mem1[132][12] , \mem1[132][11] ,
         \mem1[132][10] , \mem1[132][9] , \mem1[132][8] , \mem1[131][15] ,
         \mem1[131][14] , \mem1[131][13] , \mem1[131][12] , \mem1[131][11] ,
         \mem1[131][10] , \mem1[131][9] , \mem1[131][8] , \mem1[130][15] ,
         \mem1[130][14] , \mem1[130][13] , \mem1[130][12] , \mem1[130][11] ,
         \mem1[130][10] , \mem1[130][9] , \mem1[130][8] , \mem1[129][15] ,
         \mem1[129][14] , \mem1[129][13] , \mem1[129][12] , \mem1[129][11] ,
         \mem1[129][10] , \mem1[129][9] , \mem1[129][8] , \mem1[128][15] ,
         \mem1[128][14] , \mem1[128][13] , \mem1[128][12] , \mem1[128][11] ,
         \mem1[128][10] , \mem1[128][9] , \mem1[128][8] , \mem1[127][15] ,
         \mem1[127][14] , \mem1[127][13] , \mem1[127][12] , \mem1[127][11] ,
         \mem1[127][10] , \mem1[127][9] , \mem1[127][8] , \mem1[126][15] ,
         \mem1[126][14] , \mem1[126][13] , \mem1[126][12] , \mem1[126][11] ,
         \mem1[126][10] , \mem1[126][9] , \mem1[126][8] , \mem1[125][15] ,
         \mem1[125][14] , \mem1[125][13] , \mem1[125][12] , \mem1[125][11] ,
         \mem1[125][10] , \mem1[125][9] , \mem1[125][8] , \mem1[124][15] ,
         \mem1[124][14] , \mem1[124][13] , \mem1[124][12] , \mem1[124][11] ,
         \mem1[124][10] , \mem1[124][9] , \mem1[124][8] , \mem1[123][15] ,
         \mem1[123][14] , \mem1[123][13] , \mem1[123][12] , \mem1[123][11] ,
         \mem1[123][10] , \mem1[123][9] , \mem1[123][8] , \mem1[122][15] ,
         \mem1[122][14] , \mem1[122][13] , \mem1[122][12] , \mem1[122][11] ,
         \mem1[122][10] , \mem1[122][9] , \mem1[122][8] , \mem1[121][15] ,
         \mem1[121][14] , \mem1[121][13] , \mem1[121][12] , \mem1[121][11] ,
         \mem1[121][10] , \mem1[121][9] , \mem1[121][8] , \mem1[120][15] ,
         \mem1[120][14] , \mem1[120][13] , \mem1[120][12] , \mem1[120][11] ,
         \mem1[120][10] , \mem1[120][9] , \mem1[120][8] , \mem1[119][15] ,
         \mem1[119][14] , \mem1[119][13] , \mem1[119][12] , \mem1[119][11] ,
         \mem1[119][10] , \mem1[119][9] , \mem1[119][8] , \mem1[118][15] ,
         \mem1[118][14] , \mem1[118][13] , \mem1[118][12] , \mem1[118][11] ,
         \mem1[118][10] , \mem1[118][9] , \mem1[118][8] , \mem1[117][15] ,
         \mem1[117][14] , \mem1[117][13] , \mem1[117][12] , \mem1[117][11] ,
         \mem1[117][10] , \mem1[117][9] , \mem1[117][8] , \mem1[116][15] ,
         \mem1[116][14] , \mem1[116][13] , \mem1[116][12] , \mem1[116][11] ,
         \mem1[116][10] , \mem1[116][9] , \mem1[116][8] , \mem1[115][15] ,
         \mem1[115][14] , \mem1[115][13] , \mem1[115][12] , \mem1[115][11] ,
         \mem1[115][10] , \mem1[115][9] , \mem1[115][8] , \mem1[114][15] ,
         \mem1[114][14] , \mem1[114][13] , \mem1[114][12] , \mem1[114][11] ,
         \mem1[114][10] , \mem1[114][9] , \mem1[114][8] , \mem1[113][15] ,
         \mem1[113][14] , \mem1[113][13] , \mem1[113][12] , \mem1[113][11] ,
         \mem1[113][10] , \mem1[113][9] , \mem1[113][8] , \mem1[112][15] ,
         \mem1[112][14] , \mem1[112][13] , \mem1[112][12] , \mem1[112][11] ,
         \mem1[112][10] , \mem1[112][9] , \mem1[112][8] , \mem1[111][15] ,
         \mem1[111][14] , \mem1[111][13] , \mem1[111][12] , \mem1[111][11] ,
         \mem1[111][10] , \mem1[111][9] , \mem1[111][8] , \mem1[110][15] ,
         \mem1[110][14] , \mem1[110][13] , \mem1[110][12] , \mem1[110][11] ,
         \mem1[110][10] , \mem1[110][9] , \mem1[110][8] , \mem1[109][15] ,
         \mem1[109][14] , \mem1[109][13] , \mem1[109][12] , \mem1[109][11] ,
         \mem1[109][10] , \mem1[109][9] , \mem1[109][8] , \mem1[108][15] ,
         \mem1[108][14] , \mem1[108][13] , \mem1[108][12] , \mem1[108][11] ,
         \mem1[108][10] , \mem1[108][9] , \mem1[108][8] , \mem1[107][15] ,
         \mem1[107][14] , \mem1[107][13] , \mem1[107][12] , \mem1[107][11] ,
         \mem1[107][10] , \mem1[107][9] , \mem1[107][8] , \mem1[106][15] ,
         \mem1[106][14] , \mem1[106][13] , \mem1[106][12] , \mem1[106][11] ,
         \mem1[106][10] , \mem1[106][9] , \mem1[106][8] , \mem1[105][15] ,
         \mem1[105][14] , \mem1[105][13] , \mem1[105][12] , \mem1[105][11] ,
         \mem1[105][10] , \mem1[105][9] , \mem1[105][8] , \mem1[104][15] ,
         \mem1[104][14] , \mem1[104][13] , \mem1[104][12] , \mem1[104][11] ,
         \mem1[104][10] , \mem1[104][9] , \mem1[104][8] , \mem1[103][15] ,
         \mem1[103][14] , \mem1[103][13] , \mem1[103][12] , \mem1[103][11] ,
         \mem1[103][10] , \mem1[103][9] , \mem1[103][8] , \mem1[102][15] ,
         \mem1[102][14] , \mem1[102][13] , \mem1[102][12] , \mem1[102][11] ,
         \mem1[102][10] , \mem1[102][9] , \mem1[102][8] , \mem1[101][15] ,
         \mem1[101][14] , \mem1[101][13] , \mem1[101][12] , \mem1[101][11] ,
         \mem1[101][10] , \mem1[101][9] , \mem1[101][8] , \mem1[100][15] ,
         \mem1[100][14] , \mem1[100][13] , \mem1[100][12] , \mem1[100][11] ,
         \mem1[100][10] , \mem1[100][9] , \mem1[100][8] , \mem1[99][15] ,
         \mem1[99][14] , \mem1[99][13] , \mem1[99][12] , \mem1[99][11] ,
         \mem1[99][10] , \mem1[99][9] , \mem1[99][8] , \mem1[98][15] ,
         \mem1[98][14] , \mem1[98][13] , \mem1[98][12] , \mem1[98][11] ,
         \mem1[98][10] , \mem1[98][9] , \mem1[98][8] , \mem1[97][15] ,
         \mem1[97][14] , \mem1[97][13] , \mem1[97][12] , \mem1[97][11] ,
         \mem1[97][10] , \mem1[97][9] , \mem1[97][8] , \mem1[96][15] ,
         \mem1[96][14] , \mem1[96][13] , \mem1[96][12] , \mem1[96][11] ,
         \mem1[96][10] , \mem1[96][9] , \mem1[96][8] , \mem1[95][15] ,
         \mem1[95][14] , \mem1[95][13] , \mem1[95][12] , \mem1[95][11] ,
         \mem1[95][10] , \mem1[95][9] , \mem1[95][8] , \mem1[94][15] ,
         \mem1[94][14] , \mem1[94][13] , \mem1[94][12] , \mem1[94][11] ,
         \mem1[94][10] , \mem1[94][9] , \mem1[94][8] , \mem1[93][15] ,
         \mem1[93][14] , \mem1[93][13] , \mem1[93][12] , \mem1[93][11] ,
         \mem1[93][10] , \mem1[93][9] , \mem1[93][8] , \mem1[92][15] ,
         \mem1[92][14] , \mem1[92][13] , \mem1[92][12] , \mem1[92][11] ,
         \mem1[92][10] , \mem1[92][9] , \mem1[92][8] , \mem1[91][15] ,
         \mem1[91][14] , \mem1[91][13] , \mem1[91][12] , \mem1[91][11] ,
         \mem1[91][10] , \mem1[91][9] , \mem1[91][8] , \mem1[90][15] ,
         \mem1[90][14] , \mem1[90][13] , \mem1[90][12] , \mem1[90][11] ,
         \mem1[90][10] , \mem1[90][9] , \mem1[90][8] , \mem1[89][15] ,
         \mem1[89][14] , \mem1[89][13] , \mem1[89][12] , \mem1[89][11] ,
         \mem1[89][10] , \mem1[89][9] , \mem1[89][8] , \mem1[88][15] ,
         \mem1[88][14] , \mem1[88][13] , \mem1[88][12] , \mem1[88][11] ,
         \mem1[88][10] , \mem1[88][9] , \mem1[88][8] , \mem1[87][15] ,
         \mem1[87][14] , \mem1[87][13] , \mem1[87][12] , \mem1[87][11] ,
         \mem1[87][10] , \mem1[87][9] , \mem1[87][8] , \mem1[86][15] ,
         \mem1[86][14] , \mem1[86][13] , \mem1[86][12] , \mem1[86][11] ,
         \mem1[86][10] , \mem1[86][9] , \mem1[86][8] , \mem1[85][15] ,
         \mem1[85][14] , \mem1[85][13] , \mem1[85][12] , \mem1[85][11] ,
         \mem1[85][10] , \mem1[85][9] , \mem1[85][8] , \mem1[84][15] ,
         \mem1[84][14] , \mem1[84][13] , \mem1[84][12] , \mem1[84][11] ,
         \mem1[84][10] , \mem1[84][9] , \mem1[84][8] , \mem1[83][15] ,
         \mem1[83][14] , \mem1[83][13] , \mem1[83][12] , \mem1[83][11] ,
         \mem1[83][10] , \mem1[83][9] , \mem1[83][8] , \mem1[82][15] ,
         \mem1[82][14] , \mem1[82][13] , \mem1[82][12] , \mem1[82][11] ,
         \mem1[82][10] , \mem1[82][9] , \mem1[82][8] , \mem1[81][15] ,
         \mem1[81][14] , \mem1[81][13] , \mem1[81][12] , \mem1[81][11] ,
         \mem1[81][10] , \mem1[81][9] , \mem1[81][8] , \mem1[80][15] ,
         \mem1[80][14] , \mem1[80][13] , \mem1[80][12] , \mem1[80][11] ,
         \mem1[80][10] , \mem1[80][9] , \mem1[80][8] , \mem1[79][15] ,
         \mem1[79][14] , \mem1[79][13] , \mem1[79][12] , \mem1[79][11] ,
         \mem1[79][10] , \mem1[79][9] , \mem1[79][8] , \mem1[78][15] ,
         \mem1[78][14] , \mem1[78][13] , \mem1[78][12] , \mem1[78][11] ,
         \mem1[78][10] , \mem1[78][9] , \mem1[78][8] , \mem1[77][15] ,
         \mem1[77][14] , \mem1[77][13] , \mem1[77][12] , \mem1[77][11] ,
         \mem1[77][10] , \mem1[77][9] , \mem1[77][8] , \mem1[76][15] ,
         \mem1[76][14] , \mem1[76][13] , \mem1[76][12] , \mem1[76][11] ,
         \mem1[76][10] , \mem1[76][9] , \mem1[76][8] , \mem1[75][15] ,
         \mem1[75][14] , \mem1[75][13] , \mem1[75][12] , \mem1[75][11] ,
         \mem1[75][10] , \mem1[75][9] , \mem1[75][8] , \mem1[74][15] ,
         \mem1[74][14] , \mem1[74][13] , \mem1[74][12] , \mem1[74][11] ,
         \mem1[74][10] , \mem1[74][9] , \mem1[74][8] , \mem1[73][15] ,
         \mem1[73][14] , \mem1[73][13] , \mem1[73][12] , \mem1[73][11] ,
         \mem1[73][10] , \mem1[73][9] , \mem1[73][8] , \mem1[72][15] ,
         \mem1[72][14] , \mem1[72][13] , \mem1[72][12] , \mem1[72][11] ,
         \mem1[72][10] , \mem1[72][9] , \mem1[72][8] , \mem1[71][15] ,
         \mem1[71][14] , \mem1[71][13] , \mem1[71][12] , \mem1[71][11] ,
         \mem1[71][10] , \mem1[71][9] , \mem1[71][8] , \mem1[70][15] ,
         \mem1[70][14] , \mem1[70][13] , \mem1[70][12] , \mem1[70][11] ,
         \mem1[70][10] , \mem1[70][9] , \mem1[70][8] , \mem1[69][15] ,
         \mem1[69][14] , \mem1[69][13] , \mem1[69][12] , \mem1[69][11] ,
         \mem1[69][10] , \mem1[69][9] , \mem1[69][8] , \mem1[68][15] ,
         \mem1[68][14] , \mem1[68][13] , \mem1[68][12] , \mem1[68][11] ,
         \mem1[68][10] , \mem1[68][9] , \mem1[68][8] , \mem1[67][15] ,
         \mem1[67][14] , \mem1[67][13] , \mem1[67][12] , \mem1[67][11] ,
         \mem1[67][10] , \mem1[67][9] , \mem1[67][8] , \mem1[66][15] ,
         \mem1[66][14] , \mem1[66][13] , \mem1[66][12] , \mem1[66][11] ,
         \mem1[66][10] , \mem1[66][9] , \mem1[66][8] , \mem1[65][15] ,
         \mem1[65][14] , \mem1[65][13] , \mem1[65][12] , \mem1[65][11] ,
         \mem1[65][10] , \mem1[65][9] , \mem1[65][8] , \mem1[64][15] ,
         \mem1[64][14] , \mem1[64][13] , \mem1[64][12] , \mem1[64][11] ,
         \mem1[64][10] , \mem1[64][9] , \mem1[64][8] , \mem1[63][15] ,
         \mem1[63][14] , \mem1[63][13] , \mem1[63][12] , \mem1[63][11] ,
         \mem1[63][10] , \mem1[63][9] , \mem1[63][8] , \mem1[62][15] ,
         \mem1[62][14] , \mem1[62][13] , \mem1[62][12] , \mem1[62][11] ,
         \mem1[62][10] , \mem1[62][9] , \mem1[62][8] , \mem1[61][15] ,
         \mem1[61][14] , \mem1[61][13] , \mem1[61][12] , \mem1[61][11] ,
         \mem1[61][10] , \mem1[61][9] , \mem1[61][8] , \mem1[60][15] ,
         \mem1[60][14] , \mem1[60][13] , \mem1[60][12] , \mem1[60][11] ,
         \mem1[60][10] , \mem1[60][9] , \mem1[60][8] , \mem1[59][15] ,
         \mem1[59][14] , \mem1[59][13] , \mem1[59][12] , \mem1[59][11] ,
         \mem1[59][10] , \mem1[59][9] , \mem1[59][8] , \mem1[58][15] ,
         \mem1[58][14] , \mem1[58][13] , \mem1[58][12] , \mem1[58][11] ,
         \mem1[58][10] , \mem1[58][9] , \mem1[58][8] , \mem1[57][15] ,
         \mem1[57][14] , \mem1[57][13] , \mem1[57][12] , \mem1[57][11] ,
         \mem1[57][10] , \mem1[57][9] , \mem1[57][8] , \mem1[56][15] ,
         \mem1[56][14] , \mem1[56][13] , \mem1[56][12] , \mem1[56][11] ,
         \mem1[56][10] , \mem1[56][9] , \mem1[56][8] , \mem1[55][15] ,
         \mem1[55][14] , \mem1[55][13] , \mem1[55][12] , \mem1[55][11] ,
         \mem1[55][10] , \mem1[55][9] , \mem1[55][8] , \mem1[54][15] ,
         \mem1[54][14] , \mem1[54][13] , \mem1[54][12] , \mem1[54][11] ,
         \mem1[54][10] , \mem1[54][9] , \mem1[54][8] , \mem1[53][15] ,
         \mem1[53][14] , \mem1[53][13] , \mem1[53][12] , \mem1[53][11] ,
         \mem1[53][10] , \mem1[53][9] , \mem1[53][8] , \mem1[52][15] ,
         \mem1[52][14] , \mem1[52][13] , \mem1[52][12] , \mem1[52][11] ,
         \mem1[52][10] , \mem1[52][9] , \mem1[52][8] , \mem1[51][15] ,
         \mem1[51][14] , \mem1[51][13] , \mem1[51][12] , \mem1[51][11] ,
         \mem1[51][10] , \mem1[51][9] , \mem1[51][8] , \mem1[50][15] ,
         \mem1[50][14] , \mem1[50][13] , \mem1[50][12] , \mem1[50][11] ,
         \mem1[50][10] , \mem1[50][9] , \mem1[50][8] , \mem1[49][15] ,
         \mem1[49][14] , \mem1[49][13] , \mem1[49][12] , \mem1[49][11] ,
         \mem1[49][10] , \mem1[49][9] , \mem1[49][8] , \mem1[48][15] ,
         \mem1[48][14] , \mem1[48][13] , \mem1[48][12] , \mem1[48][11] ,
         \mem1[48][10] , \mem1[48][9] , \mem1[48][8] , \mem1[47][15] ,
         \mem1[47][14] , \mem1[47][13] , \mem1[47][12] , \mem1[47][11] ,
         \mem1[47][10] , \mem1[47][9] , \mem1[47][8] , \mem1[46][15] ,
         \mem1[46][14] , \mem1[46][13] , \mem1[46][12] , \mem1[46][11] ,
         \mem1[46][10] , \mem1[46][9] , \mem1[46][8] , \mem1[45][15] ,
         \mem1[45][14] , \mem1[45][13] , \mem1[45][12] , \mem1[45][11] ,
         \mem1[45][10] , \mem1[45][9] , \mem1[45][8] , \mem1[44][15] ,
         \mem1[44][14] , \mem1[44][13] , \mem1[44][12] , \mem1[44][11] ,
         \mem1[44][10] , \mem1[44][9] , \mem1[44][8] , \mem1[43][15] ,
         \mem1[43][14] , \mem1[43][13] , \mem1[43][12] , \mem1[43][11] ,
         \mem1[43][10] , \mem1[43][9] , \mem1[43][8] , \mem1[42][15] ,
         \mem1[42][14] , \mem1[42][13] , \mem1[42][12] , \mem1[42][11] ,
         \mem1[42][10] , \mem1[42][9] , \mem1[42][8] , \mem1[41][15] ,
         \mem1[41][14] , \mem1[41][13] , \mem1[41][12] , \mem1[41][11] ,
         \mem1[41][10] , \mem1[41][9] , \mem1[41][8] , \mem1[40][15] ,
         \mem1[40][14] , \mem1[40][13] , \mem1[40][12] , \mem1[40][11] ,
         \mem1[40][10] , \mem1[40][9] , \mem1[40][8] , \mem1[39][15] ,
         \mem1[39][14] , \mem1[39][13] , \mem1[39][12] , \mem1[39][11] ,
         \mem1[39][10] , \mem1[39][9] , \mem1[39][8] , \mem1[38][15] ,
         \mem1[38][14] , \mem1[38][13] , \mem1[38][12] , \mem1[38][11] ,
         \mem1[38][10] , \mem1[38][9] , \mem1[38][8] , \mem1[37][15] ,
         \mem1[37][14] , \mem1[37][13] , \mem1[37][12] , \mem1[37][11] ,
         \mem1[37][10] , \mem1[37][9] , \mem1[37][8] , \mem1[36][15] ,
         \mem1[36][14] , \mem1[36][13] , \mem1[36][12] , \mem1[36][11] ,
         \mem1[36][10] , \mem1[36][9] , \mem1[36][8] , \mem1[35][15] ,
         \mem1[35][14] , \mem1[35][13] , \mem1[35][12] , \mem1[35][11] ,
         \mem1[35][10] , \mem1[35][9] , \mem1[35][8] , \mem1[34][15] ,
         \mem1[34][14] , \mem1[34][13] , \mem1[34][12] , \mem1[34][11] ,
         \mem1[34][10] , \mem1[34][9] , \mem1[34][8] , \mem1[33][15] ,
         \mem1[33][14] , \mem1[33][13] , \mem1[33][12] , \mem1[33][11] ,
         \mem1[33][10] , \mem1[33][9] , \mem1[33][8] , \mem1[32][15] ,
         \mem1[32][14] , \mem1[32][13] , \mem1[32][12] , \mem1[32][11] ,
         \mem1[32][10] , \mem1[32][9] , \mem1[32][8] , \mem1[31][15] ,
         \mem1[31][14] , \mem1[31][13] , \mem1[31][12] , \mem1[31][11] ,
         \mem1[31][10] , \mem1[31][9] , \mem1[31][8] , \mem1[30][15] ,
         \mem1[30][14] , \mem1[30][13] , \mem1[30][12] , \mem1[30][11] ,
         \mem1[30][10] , \mem1[30][9] , \mem1[30][8] , \mem1[29][15] ,
         \mem1[29][14] , \mem1[29][13] , \mem1[29][12] , \mem1[29][11] ,
         \mem1[29][10] , \mem1[29][9] , \mem1[29][8] , \mem1[28][15] ,
         \mem1[28][14] , \mem1[28][13] , \mem1[28][12] , \mem1[28][11] ,
         \mem1[28][10] , \mem1[28][9] , \mem1[28][8] , \mem1[27][15] ,
         \mem1[27][14] , \mem1[27][13] , \mem1[27][12] , \mem1[27][11] ,
         \mem1[27][10] , \mem1[27][9] , \mem1[27][8] , \mem1[26][15] ,
         \mem1[26][14] , \mem1[26][13] , \mem1[26][12] , \mem1[26][11] ,
         \mem1[26][10] , \mem1[26][9] , \mem1[26][8] , \mem1[25][15] ,
         \mem1[25][14] , \mem1[25][13] , \mem1[25][12] , \mem1[25][11] ,
         \mem1[25][10] , \mem1[25][9] , \mem1[25][8] , \mem1[24][15] ,
         \mem1[24][14] , \mem1[24][13] , \mem1[24][12] , \mem1[24][11] ,
         \mem1[24][10] , \mem1[24][9] , \mem1[24][8] , \mem1[23][15] ,
         \mem1[23][14] , \mem1[23][13] , \mem1[23][12] , \mem1[23][11] ,
         \mem1[23][10] , \mem1[23][9] , \mem1[23][8] , \mem1[22][15] ,
         \mem1[22][14] , \mem1[22][13] , \mem1[22][12] , \mem1[22][11] ,
         \mem1[22][10] , \mem1[22][9] , \mem1[22][8] , \mem1[21][15] ,
         \mem1[21][14] , \mem1[21][13] , \mem1[21][12] , \mem1[21][11] ,
         \mem1[21][10] , \mem1[21][9] , \mem1[21][8] , \mem1[20][15] ,
         \mem1[20][14] , \mem1[20][13] , \mem1[20][12] , \mem1[20][11] ,
         \mem1[20][10] , \mem1[20][9] , \mem1[20][8] , \mem1[19][15] ,
         \mem1[19][14] , \mem1[19][13] , \mem1[19][12] , \mem1[19][11] ,
         \mem1[19][10] , \mem1[19][9] , \mem1[19][8] , \mem1[18][15] ,
         \mem1[18][14] , \mem1[18][13] , \mem1[18][12] , \mem1[18][11] ,
         \mem1[18][10] , \mem1[18][9] , \mem1[18][8] , \mem1[17][15] ,
         \mem1[17][14] , \mem1[17][13] , \mem1[17][12] , \mem1[17][11] ,
         \mem1[17][10] , \mem1[17][9] , \mem1[17][8] , \mem1[16][15] ,
         \mem1[16][14] , \mem1[16][13] , \mem1[16][12] , \mem1[16][11] ,
         \mem1[16][10] , \mem1[16][9] , \mem1[16][8] , \mem1[15][15] ,
         \mem1[15][14] , \mem1[15][13] , \mem1[15][12] , \mem1[15][11] ,
         \mem1[15][10] , \mem1[15][9] , \mem1[15][8] , \mem1[14][15] ,
         \mem1[14][14] , \mem1[14][13] , \mem1[14][12] , \mem1[14][11] ,
         \mem1[14][10] , \mem1[14][9] , \mem1[14][8] , \mem1[13][15] ,
         \mem1[13][14] , \mem1[13][13] , \mem1[13][12] , \mem1[13][11] ,
         \mem1[13][10] , \mem1[13][9] , \mem1[13][8] , \mem1[12][15] ,
         \mem1[12][14] , \mem1[12][13] , \mem1[12][12] , \mem1[12][11] ,
         \mem1[12][10] , \mem1[12][9] , \mem1[12][8] , \mem1[11][15] ,
         \mem1[11][14] , \mem1[11][13] , \mem1[11][12] , \mem1[11][11] ,
         \mem1[11][10] , \mem1[11][9] , \mem1[11][8] , \mem1[10][15] ,
         \mem1[10][14] , \mem1[10][13] , \mem1[10][12] , \mem1[10][11] ,
         \mem1[10][10] , \mem1[10][9] , \mem1[10][8] , \mem1[9][15] ,
         \mem1[9][14] , \mem1[9][13] , \mem1[9][12] , \mem1[9][11] ,
         \mem1[9][10] , \mem1[9][9] , \mem1[9][8] , \mem1[8][15] ,
         \mem1[8][14] , \mem1[8][13] , \mem1[8][12] , \mem1[8][11] ,
         \mem1[8][10] , \mem1[8][9] , \mem1[8][8] , \mem1[7][15] ,
         \mem1[7][14] , \mem1[7][13] , \mem1[7][12] , \mem1[7][11] ,
         \mem1[7][10] , \mem1[7][9] , \mem1[7][8] , \mem1[6][15] ,
         \mem1[6][14] , \mem1[6][13] , \mem1[6][12] , \mem1[6][11] ,
         \mem1[6][10] , \mem1[6][9] , \mem1[6][8] , \mem1[5][15] ,
         \mem1[5][14] , \mem1[5][13] , \mem1[5][12] , \mem1[5][11] ,
         \mem1[5][10] , \mem1[5][9] , \mem1[5][8] , \mem1[4][15] ,
         \mem1[4][14] , \mem1[4][13] , \mem1[4][12] , \mem1[4][11] ,
         \mem1[4][10] , \mem1[4][9] , \mem1[4][8] , \mem1[3][15] ,
         \mem1[3][14] , \mem1[3][13] , \mem1[3][12] , \mem1[3][11] ,
         \mem1[3][10] , \mem1[3][9] , \mem1[3][8] , \mem1[2][15] ,
         \mem1[2][14] , \mem1[2][13] , \mem1[2][12] , \mem1[2][11] ,
         \mem1[2][10] , \mem1[2][9] , \mem1[2][8] , \mem1[1][15] ,
         \mem1[1][14] , \mem1[1][13] , \mem1[1][12] , \mem1[1][11] ,
         \mem1[1][10] , \mem1[1][9] , \mem1[1][8] , \mem1[0][15] ,
         \mem1[0][14] , \mem1[0][13] , \mem1[0][12] , \mem1[0][11] ,
         \mem1[0][10] , \mem1[0][9] , \mem1[0][8] , \mem0[255][7] ,
         \mem0[255][6] , \mem0[255][5] , \mem0[255][4] , \mem0[255][3] ,
         \mem0[255][2] , \mem0[255][1] , \mem0[255][0] , \mem0[254][7] ,
         \mem0[254][6] , \mem0[254][5] , \mem0[254][4] , \mem0[254][3] ,
         \mem0[254][2] , \mem0[254][1] , \mem0[254][0] , \mem0[253][7] ,
         \mem0[253][6] , \mem0[253][5] , \mem0[253][4] , \mem0[253][3] ,
         \mem0[253][2] , \mem0[253][1] , \mem0[253][0] , \mem0[252][7] ,
         \mem0[252][6] , \mem0[252][5] , \mem0[252][4] , \mem0[252][3] ,
         \mem0[252][2] , \mem0[252][1] , \mem0[252][0] , \mem0[251][7] ,
         \mem0[251][6] , \mem0[251][5] , \mem0[251][4] , \mem0[251][3] ,
         \mem0[251][2] , \mem0[251][1] , \mem0[251][0] , \mem0[250][7] ,
         \mem0[250][6] , \mem0[250][5] , \mem0[250][4] , \mem0[250][3] ,
         \mem0[250][2] , \mem0[250][1] , \mem0[250][0] , \mem0[249][7] ,
         \mem0[249][6] , \mem0[249][5] , \mem0[249][4] , \mem0[249][3] ,
         \mem0[249][2] , \mem0[249][1] , \mem0[249][0] , \mem0[248][7] ,
         \mem0[248][6] , \mem0[248][5] , \mem0[248][4] , \mem0[248][3] ,
         \mem0[248][2] , \mem0[248][1] , \mem0[248][0] , \mem0[247][7] ,
         \mem0[247][6] , \mem0[247][5] , \mem0[247][4] , \mem0[247][3] ,
         \mem0[247][2] , \mem0[247][1] , \mem0[247][0] , \mem0[246][7] ,
         \mem0[246][6] , \mem0[246][5] , \mem0[246][4] , \mem0[246][3] ,
         \mem0[246][2] , \mem0[246][1] , \mem0[246][0] , \mem0[245][7] ,
         \mem0[245][6] , \mem0[245][5] , \mem0[245][4] , \mem0[245][3] ,
         \mem0[245][2] , \mem0[245][1] , \mem0[245][0] , \mem0[244][7] ,
         \mem0[244][6] , \mem0[244][5] , \mem0[244][4] , \mem0[244][3] ,
         \mem0[244][2] , \mem0[244][1] , \mem0[244][0] , \mem0[243][7] ,
         \mem0[243][6] , \mem0[243][5] , \mem0[243][4] , \mem0[243][3] ,
         \mem0[243][2] , \mem0[243][1] , \mem0[243][0] , \mem0[242][7] ,
         \mem0[242][6] , \mem0[242][5] , \mem0[242][4] , \mem0[242][3] ,
         \mem0[242][2] , \mem0[242][1] , \mem0[242][0] , \mem0[241][7] ,
         \mem0[241][6] , \mem0[241][5] , \mem0[241][4] , \mem0[241][3] ,
         \mem0[241][2] , \mem0[241][1] , \mem0[241][0] , \mem0[240][7] ,
         \mem0[240][6] , \mem0[240][5] , \mem0[240][4] , \mem0[240][3] ,
         \mem0[240][2] , \mem0[240][1] , \mem0[240][0] , \mem0[239][7] ,
         \mem0[239][6] , \mem0[239][5] , \mem0[239][4] , \mem0[239][3] ,
         \mem0[239][2] , \mem0[239][1] , \mem0[239][0] , \mem0[238][7] ,
         \mem0[238][6] , \mem0[238][5] , \mem0[238][4] , \mem0[238][3] ,
         \mem0[238][2] , \mem0[238][1] , \mem0[238][0] , \mem0[237][7] ,
         \mem0[237][6] , \mem0[237][5] , \mem0[237][4] , \mem0[237][3] ,
         \mem0[237][2] , \mem0[237][1] , \mem0[237][0] , \mem0[236][7] ,
         \mem0[236][6] , \mem0[236][5] , \mem0[236][4] , \mem0[236][3] ,
         \mem0[236][2] , \mem0[236][1] , \mem0[236][0] , \mem0[235][7] ,
         \mem0[235][6] , \mem0[235][5] , \mem0[235][4] , \mem0[235][3] ,
         \mem0[235][2] , \mem0[235][1] , \mem0[235][0] , \mem0[234][7] ,
         \mem0[234][6] , \mem0[234][5] , \mem0[234][4] , \mem0[234][3] ,
         \mem0[234][2] , \mem0[234][1] , \mem0[234][0] , \mem0[233][7] ,
         \mem0[233][6] , \mem0[233][5] , \mem0[233][4] , \mem0[233][3] ,
         \mem0[233][2] , \mem0[233][1] , \mem0[233][0] , \mem0[232][7] ,
         \mem0[232][6] , \mem0[232][5] , \mem0[232][4] , \mem0[232][3] ,
         \mem0[232][2] , \mem0[232][1] , \mem0[232][0] , \mem0[231][7] ,
         \mem0[231][6] , \mem0[231][5] , \mem0[231][4] , \mem0[231][3] ,
         \mem0[231][2] , \mem0[231][1] , \mem0[231][0] , \mem0[230][7] ,
         \mem0[230][6] , \mem0[230][5] , \mem0[230][4] , \mem0[230][3] ,
         \mem0[230][2] , \mem0[230][1] , \mem0[230][0] , \mem0[229][7] ,
         \mem0[229][6] , \mem0[229][5] , \mem0[229][4] , \mem0[229][3] ,
         \mem0[229][2] , \mem0[229][1] , \mem0[229][0] , \mem0[228][7] ,
         \mem0[228][6] , \mem0[228][5] , \mem0[228][4] , \mem0[228][3] ,
         \mem0[228][2] , \mem0[228][1] , \mem0[228][0] , \mem0[227][7] ,
         \mem0[227][6] , \mem0[227][5] , \mem0[227][4] , \mem0[227][3] ,
         \mem0[227][2] , \mem0[227][1] , \mem0[227][0] , \mem0[226][7] ,
         \mem0[226][6] , \mem0[226][5] , \mem0[226][4] , \mem0[226][3] ,
         \mem0[226][2] , \mem0[226][1] , \mem0[226][0] , \mem0[225][7] ,
         \mem0[225][6] , \mem0[225][5] , \mem0[225][4] , \mem0[225][3] ,
         \mem0[225][2] , \mem0[225][1] , \mem0[225][0] , \mem0[224][7] ,
         \mem0[224][6] , \mem0[224][5] , \mem0[224][4] , \mem0[224][3] ,
         \mem0[224][2] , \mem0[224][1] , \mem0[224][0] , \mem0[223][7] ,
         \mem0[223][6] , \mem0[223][5] , \mem0[223][4] , \mem0[223][3] ,
         \mem0[223][2] , \mem0[223][1] , \mem0[223][0] , \mem0[222][7] ,
         \mem0[222][6] , \mem0[222][5] , \mem0[222][4] , \mem0[222][3] ,
         \mem0[222][2] , \mem0[222][1] , \mem0[222][0] , \mem0[221][7] ,
         \mem0[221][6] , \mem0[221][5] , \mem0[221][4] , \mem0[221][3] ,
         \mem0[221][2] , \mem0[221][1] , \mem0[221][0] , \mem0[220][7] ,
         \mem0[220][6] , \mem0[220][5] , \mem0[220][4] , \mem0[220][3] ,
         \mem0[220][2] , \mem0[220][1] , \mem0[220][0] , \mem0[219][7] ,
         \mem0[219][6] , \mem0[219][5] , \mem0[219][4] , \mem0[219][3] ,
         \mem0[219][2] , \mem0[219][1] , \mem0[219][0] , \mem0[218][7] ,
         \mem0[218][6] , \mem0[218][5] , \mem0[218][4] , \mem0[218][3] ,
         \mem0[218][2] , \mem0[218][1] , \mem0[218][0] , \mem0[217][7] ,
         \mem0[217][6] , \mem0[217][5] , \mem0[217][4] , \mem0[217][3] ,
         \mem0[217][2] , \mem0[217][1] , \mem0[217][0] , \mem0[216][7] ,
         \mem0[216][6] , \mem0[216][5] , \mem0[216][4] , \mem0[216][3] ,
         \mem0[216][2] , \mem0[216][1] , \mem0[216][0] , \mem0[215][7] ,
         \mem0[215][6] , \mem0[215][5] , \mem0[215][4] , \mem0[215][3] ,
         \mem0[215][2] , \mem0[215][1] , \mem0[215][0] , \mem0[214][7] ,
         \mem0[214][6] , \mem0[214][5] , \mem0[214][4] , \mem0[214][3] ,
         \mem0[214][2] , \mem0[214][1] , \mem0[214][0] , \mem0[213][7] ,
         \mem0[213][6] , \mem0[213][5] , \mem0[213][4] , \mem0[213][3] ,
         \mem0[213][2] , \mem0[213][1] , \mem0[213][0] , \mem0[212][7] ,
         \mem0[212][6] , \mem0[212][5] , \mem0[212][4] , \mem0[212][3] ,
         \mem0[212][2] , \mem0[212][1] , \mem0[212][0] , \mem0[211][7] ,
         \mem0[211][6] , \mem0[211][5] , \mem0[211][4] , \mem0[211][3] ,
         \mem0[211][2] , \mem0[211][1] , \mem0[211][0] , \mem0[210][7] ,
         \mem0[210][6] , \mem0[210][5] , \mem0[210][4] , \mem0[210][3] ,
         \mem0[210][2] , \mem0[210][1] , \mem0[210][0] , \mem0[209][7] ,
         \mem0[209][6] , \mem0[209][5] , \mem0[209][4] , \mem0[209][3] ,
         \mem0[209][2] , \mem0[209][1] , \mem0[209][0] , \mem0[208][7] ,
         \mem0[208][6] , \mem0[208][5] , \mem0[208][4] , \mem0[208][3] ,
         \mem0[208][2] , \mem0[208][1] , \mem0[208][0] , \mem0[207][7] ,
         \mem0[207][6] , \mem0[207][5] , \mem0[207][4] , \mem0[207][3] ,
         \mem0[207][2] , \mem0[207][1] , \mem0[207][0] , \mem0[206][7] ,
         \mem0[206][6] , \mem0[206][5] , \mem0[206][4] , \mem0[206][3] ,
         \mem0[206][2] , \mem0[206][1] , \mem0[206][0] , \mem0[205][7] ,
         \mem0[205][6] , \mem0[205][5] , \mem0[205][4] , \mem0[205][3] ,
         \mem0[205][2] , \mem0[205][1] , \mem0[205][0] , \mem0[204][7] ,
         \mem0[204][6] , \mem0[204][5] , \mem0[204][4] , \mem0[204][3] ,
         \mem0[204][2] , \mem0[204][1] , \mem0[204][0] , \mem0[203][7] ,
         \mem0[203][6] , \mem0[203][5] , \mem0[203][4] , \mem0[203][3] ,
         \mem0[203][2] , \mem0[203][1] , \mem0[203][0] , \mem0[202][7] ,
         \mem0[202][6] , \mem0[202][5] , \mem0[202][4] , \mem0[202][3] ,
         \mem0[202][2] , \mem0[202][1] , \mem0[202][0] , \mem0[201][7] ,
         \mem0[201][6] , \mem0[201][5] , \mem0[201][4] , \mem0[201][3] ,
         \mem0[201][2] , \mem0[201][1] , \mem0[201][0] , \mem0[200][7] ,
         \mem0[200][6] , \mem0[200][5] , \mem0[200][4] , \mem0[200][3] ,
         \mem0[200][2] , \mem0[200][1] , \mem0[200][0] , \mem0[199][7] ,
         \mem0[199][6] , \mem0[199][5] , \mem0[199][4] , \mem0[199][3] ,
         \mem0[199][2] , \mem0[199][1] , \mem0[199][0] , \mem0[198][7] ,
         \mem0[198][6] , \mem0[198][5] , \mem0[198][4] , \mem0[198][3] ,
         \mem0[198][2] , \mem0[198][1] , \mem0[198][0] , \mem0[197][7] ,
         \mem0[197][6] , \mem0[197][5] , \mem0[197][4] , \mem0[197][3] ,
         \mem0[197][2] , \mem0[197][1] , \mem0[197][0] , \mem0[196][7] ,
         \mem0[196][6] , \mem0[196][5] , \mem0[196][4] , \mem0[196][3] ,
         \mem0[196][2] , \mem0[196][1] , \mem0[196][0] , \mem0[195][7] ,
         \mem0[195][6] , \mem0[195][5] , \mem0[195][4] , \mem0[195][3] ,
         \mem0[195][2] , \mem0[195][1] , \mem0[195][0] , \mem0[194][7] ,
         \mem0[194][6] , \mem0[194][5] , \mem0[194][4] , \mem0[194][3] ,
         \mem0[194][2] , \mem0[194][1] , \mem0[194][0] , \mem0[193][7] ,
         \mem0[193][6] , \mem0[193][5] , \mem0[193][4] , \mem0[193][3] ,
         \mem0[193][2] , \mem0[193][1] , \mem0[193][0] , \mem0[192][7] ,
         \mem0[192][6] , \mem0[192][5] , \mem0[192][4] , \mem0[192][3] ,
         \mem0[192][2] , \mem0[192][1] , \mem0[192][0] , \mem0[191][7] ,
         \mem0[191][6] , \mem0[191][5] , \mem0[191][4] , \mem0[191][3] ,
         \mem0[191][2] , \mem0[191][1] , \mem0[191][0] , \mem0[190][7] ,
         \mem0[190][6] , \mem0[190][5] , \mem0[190][4] , \mem0[190][3] ,
         \mem0[190][2] , \mem0[190][1] , \mem0[190][0] , \mem0[189][7] ,
         \mem0[189][6] , \mem0[189][5] , \mem0[189][4] , \mem0[189][3] ,
         \mem0[189][2] , \mem0[189][1] , \mem0[189][0] , \mem0[188][7] ,
         \mem0[188][6] , \mem0[188][5] , \mem0[188][4] , \mem0[188][3] ,
         \mem0[188][2] , \mem0[188][1] , \mem0[188][0] , \mem0[187][7] ,
         \mem0[187][6] , \mem0[187][5] , \mem0[187][4] , \mem0[187][3] ,
         \mem0[187][2] , \mem0[187][1] , \mem0[187][0] , \mem0[186][7] ,
         \mem0[186][6] , \mem0[186][5] , \mem0[186][4] , \mem0[186][3] ,
         \mem0[186][2] , \mem0[186][1] , \mem0[186][0] , \mem0[185][7] ,
         \mem0[185][6] , \mem0[185][5] , \mem0[185][4] , \mem0[185][3] ,
         \mem0[185][2] , \mem0[185][1] , \mem0[185][0] , \mem0[184][7] ,
         \mem0[184][6] , \mem0[184][5] , \mem0[184][4] , \mem0[184][3] ,
         \mem0[184][2] , \mem0[184][1] , \mem0[184][0] , \mem0[183][7] ,
         \mem0[183][6] , \mem0[183][5] , \mem0[183][4] , \mem0[183][3] ,
         \mem0[183][2] , \mem0[183][1] , \mem0[183][0] , \mem0[182][7] ,
         \mem0[182][6] , \mem0[182][5] , \mem0[182][4] , \mem0[182][3] ,
         \mem0[182][2] , \mem0[182][1] , \mem0[182][0] , \mem0[181][7] ,
         \mem0[181][6] , \mem0[181][5] , \mem0[181][4] , \mem0[181][3] ,
         \mem0[181][2] , \mem0[181][1] , \mem0[181][0] , \mem0[180][7] ,
         \mem0[180][6] , \mem0[180][5] , \mem0[180][4] , \mem0[180][3] ,
         \mem0[180][2] , \mem0[180][1] , \mem0[180][0] , \mem0[179][7] ,
         \mem0[179][6] , \mem0[179][5] , \mem0[179][4] , \mem0[179][3] ,
         \mem0[179][2] , \mem0[179][1] , \mem0[179][0] , \mem0[178][7] ,
         \mem0[178][6] , \mem0[178][5] , \mem0[178][4] , \mem0[178][3] ,
         \mem0[178][2] , \mem0[178][1] , \mem0[178][0] , \mem0[177][7] ,
         \mem0[177][6] , \mem0[177][5] , \mem0[177][4] , \mem0[177][3] ,
         \mem0[177][2] , \mem0[177][1] , \mem0[177][0] , \mem0[176][7] ,
         \mem0[176][6] , \mem0[176][5] , \mem0[176][4] , \mem0[176][3] ,
         \mem0[176][2] , \mem0[176][1] , \mem0[176][0] , \mem0[175][7] ,
         \mem0[175][6] , \mem0[175][5] , \mem0[175][4] , \mem0[175][3] ,
         \mem0[175][2] , \mem0[175][1] , \mem0[175][0] , \mem0[174][7] ,
         \mem0[174][6] , \mem0[174][5] , \mem0[174][4] , \mem0[174][3] ,
         \mem0[174][2] , \mem0[174][1] , \mem0[174][0] , \mem0[173][7] ,
         \mem0[173][6] , \mem0[173][5] , \mem0[173][4] , \mem0[173][3] ,
         \mem0[173][2] , \mem0[173][1] , \mem0[173][0] , \mem0[172][7] ,
         \mem0[172][6] , \mem0[172][5] , \mem0[172][4] , \mem0[172][3] ,
         \mem0[172][2] , \mem0[172][1] , \mem0[172][0] , \mem0[171][7] ,
         \mem0[171][6] , \mem0[171][5] , \mem0[171][4] , \mem0[171][3] ,
         \mem0[171][2] , \mem0[171][1] , \mem0[171][0] , \mem0[170][7] ,
         \mem0[170][6] , \mem0[170][5] , \mem0[170][4] , \mem0[170][3] ,
         \mem0[170][2] , \mem0[170][1] , \mem0[170][0] , \mem0[169][7] ,
         \mem0[169][6] , \mem0[169][5] , \mem0[169][4] , \mem0[169][3] ,
         \mem0[169][2] , \mem0[169][1] , \mem0[169][0] , \mem0[168][7] ,
         \mem0[168][6] , \mem0[168][5] , \mem0[168][4] , \mem0[168][3] ,
         \mem0[168][2] , \mem0[168][1] , \mem0[168][0] , \mem0[167][7] ,
         \mem0[167][6] , \mem0[167][5] , \mem0[167][4] , \mem0[167][3] ,
         \mem0[167][2] , \mem0[167][1] , \mem0[167][0] , \mem0[166][7] ,
         \mem0[166][6] , \mem0[166][5] , \mem0[166][4] , \mem0[166][3] ,
         \mem0[166][2] , \mem0[166][1] , \mem0[166][0] , \mem0[165][7] ,
         \mem0[165][6] , \mem0[165][5] , \mem0[165][4] , \mem0[165][3] ,
         \mem0[165][2] , \mem0[165][1] , \mem0[165][0] , \mem0[164][7] ,
         \mem0[164][6] , \mem0[164][5] , \mem0[164][4] , \mem0[164][3] ,
         \mem0[164][2] , \mem0[164][1] , \mem0[164][0] , \mem0[163][7] ,
         \mem0[163][6] , \mem0[163][5] , \mem0[163][4] , \mem0[163][3] ,
         \mem0[163][2] , \mem0[163][1] , \mem0[163][0] , \mem0[162][7] ,
         \mem0[162][6] , \mem0[162][5] , \mem0[162][4] , \mem0[162][3] ,
         \mem0[162][2] , \mem0[162][1] , \mem0[162][0] , \mem0[161][7] ,
         \mem0[161][6] , \mem0[161][5] , \mem0[161][4] , \mem0[161][3] ,
         \mem0[161][2] , \mem0[161][1] , \mem0[161][0] , \mem0[160][7] ,
         \mem0[160][6] , \mem0[160][5] , \mem0[160][4] , \mem0[160][3] ,
         \mem0[160][2] , \mem0[160][1] , \mem0[160][0] , \mem0[159][7] ,
         \mem0[159][6] , \mem0[159][5] , \mem0[159][4] , \mem0[159][3] ,
         \mem0[159][2] , \mem0[159][1] , \mem0[159][0] , \mem0[158][7] ,
         \mem0[158][6] , \mem0[158][5] , \mem0[158][4] , \mem0[158][3] ,
         \mem0[158][2] , \mem0[158][1] , \mem0[158][0] , \mem0[157][7] ,
         \mem0[157][6] , \mem0[157][5] , \mem0[157][4] , \mem0[157][3] ,
         \mem0[157][2] , \mem0[157][1] , \mem0[157][0] , \mem0[156][7] ,
         \mem0[156][6] , \mem0[156][5] , \mem0[156][4] , \mem0[156][3] ,
         \mem0[156][2] , \mem0[156][1] , \mem0[156][0] , \mem0[155][7] ,
         \mem0[155][6] , \mem0[155][5] , \mem0[155][4] , \mem0[155][3] ,
         \mem0[155][2] , \mem0[155][1] , \mem0[155][0] , \mem0[154][7] ,
         \mem0[154][6] , \mem0[154][5] , \mem0[154][4] , \mem0[154][3] ,
         \mem0[154][2] , \mem0[154][1] , \mem0[154][0] , \mem0[153][7] ,
         \mem0[153][6] , \mem0[153][5] , \mem0[153][4] , \mem0[153][3] ,
         \mem0[153][2] , \mem0[153][1] , \mem0[153][0] , \mem0[152][7] ,
         \mem0[152][6] , \mem0[152][5] , \mem0[152][4] , \mem0[152][3] ,
         \mem0[152][2] , \mem0[152][1] , \mem0[152][0] , \mem0[151][7] ,
         \mem0[151][6] , \mem0[151][5] , \mem0[151][4] , \mem0[151][3] ,
         \mem0[151][2] , \mem0[151][1] , \mem0[151][0] , \mem0[150][7] ,
         \mem0[150][6] , \mem0[150][5] , \mem0[150][4] , \mem0[150][3] ,
         \mem0[150][2] , \mem0[150][1] , \mem0[150][0] , \mem0[149][7] ,
         \mem0[149][6] , \mem0[149][5] , \mem0[149][4] , \mem0[149][3] ,
         \mem0[149][2] , \mem0[149][1] , \mem0[149][0] , \mem0[148][7] ,
         \mem0[148][6] , \mem0[148][5] , \mem0[148][4] , \mem0[148][3] ,
         \mem0[148][2] , \mem0[148][1] , \mem0[148][0] , \mem0[147][7] ,
         \mem0[147][6] , \mem0[147][5] , \mem0[147][4] , \mem0[147][3] ,
         \mem0[147][2] , \mem0[147][1] , \mem0[147][0] , \mem0[146][7] ,
         \mem0[146][6] , \mem0[146][5] , \mem0[146][4] , \mem0[146][3] ,
         \mem0[146][2] , \mem0[146][1] , \mem0[146][0] , \mem0[145][7] ,
         \mem0[145][6] , \mem0[145][5] , \mem0[145][4] , \mem0[145][3] ,
         \mem0[145][2] , \mem0[145][1] , \mem0[145][0] , \mem0[144][7] ,
         \mem0[144][6] , \mem0[144][5] , \mem0[144][4] , \mem0[144][3] ,
         \mem0[144][2] , \mem0[144][1] , \mem0[144][0] , \mem0[143][7] ,
         \mem0[143][6] , \mem0[143][5] , \mem0[143][4] , \mem0[143][3] ,
         \mem0[143][2] , \mem0[143][1] , \mem0[143][0] , \mem0[142][7] ,
         \mem0[142][6] , \mem0[142][5] , \mem0[142][4] , \mem0[142][3] ,
         \mem0[142][2] , \mem0[142][1] , \mem0[142][0] , \mem0[141][7] ,
         \mem0[141][6] , \mem0[141][5] , \mem0[141][4] , \mem0[141][3] ,
         \mem0[141][2] , \mem0[141][1] , \mem0[141][0] , \mem0[140][7] ,
         \mem0[140][6] , \mem0[140][5] , \mem0[140][4] , \mem0[140][3] ,
         \mem0[140][2] , \mem0[140][1] , \mem0[140][0] , \mem0[139][7] ,
         \mem0[139][6] , \mem0[139][5] , \mem0[139][4] , \mem0[139][3] ,
         \mem0[139][2] , \mem0[139][1] , \mem0[139][0] , \mem0[138][7] ,
         \mem0[138][6] , \mem0[138][5] , \mem0[138][4] , \mem0[138][3] ,
         \mem0[138][2] , \mem0[138][1] , \mem0[138][0] , \mem0[137][7] ,
         \mem0[137][6] , \mem0[137][5] , \mem0[137][4] , \mem0[137][3] ,
         \mem0[137][2] , \mem0[137][1] , \mem0[137][0] , \mem0[136][7] ,
         \mem0[136][6] , \mem0[136][5] , \mem0[136][4] , \mem0[136][3] ,
         \mem0[136][2] , \mem0[136][1] , \mem0[136][0] , \mem0[135][7] ,
         \mem0[135][6] , \mem0[135][5] , \mem0[135][4] , \mem0[135][3] ,
         \mem0[135][2] , \mem0[135][1] , \mem0[135][0] , \mem0[134][7] ,
         \mem0[134][6] , \mem0[134][5] , \mem0[134][4] , \mem0[134][3] ,
         \mem0[134][2] , \mem0[134][1] , \mem0[134][0] , \mem0[133][7] ,
         \mem0[133][6] , \mem0[133][5] , \mem0[133][4] , \mem0[133][3] ,
         \mem0[133][2] , \mem0[133][1] , \mem0[133][0] , \mem0[132][7] ,
         \mem0[132][6] , \mem0[132][5] , \mem0[132][4] , \mem0[132][3] ,
         \mem0[132][2] , \mem0[132][1] , \mem0[132][0] , \mem0[131][7] ,
         \mem0[131][6] , \mem0[131][5] , \mem0[131][4] , \mem0[131][3] ,
         \mem0[131][2] , \mem0[131][1] , \mem0[131][0] , \mem0[130][7] ,
         \mem0[130][6] , \mem0[130][5] , \mem0[130][4] , \mem0[130][3] ,
         \mem0[130][2] , \mem0[130][1] , \mem0[130][0] , \mem0[129][7] ,
         \mem0[129][6] , \mem0[129][5] , \mem0[129][4] , \mem0[129][3] ,
         \mem0[129][2] , \mem0[129][1] , \mem0[129][0] , \mem0[128][7] ,
         \mem0[128][6] , \mem0[128][5] , \mem0[128][4] , \mem0[128][3] ,
         \mem0[128][2] , \mem0[128][1] , \mem0[128][0] , \mem0[127][7] ,
         \mem0[127][6] , \mem0[127][5] , \mem0[127][4] , \mem0[127][3] ,
         \mem0[127][2] , \mem0[127][1] , \mem0[127][0] , \mem0[126][7] ,
         \mem0[126][6] , \mem0[126][5] , \mem0[126][4] , \mem0[126][3] ,
         \mem0[126][2] , \mem0[126][1] , \mem0[126][0] , \mem0[125][7] ,
         \mem0[125][6] , \mem0[125][5] , \mem0[125][4] , \mem0[125][3] ,
         \mem0[125][2] , \mem0[125][1] , \mem0[125][0] , \mem0[124][7] ,
         \mem0[124][6] , \mem0[124][5] , \mem0[124][4] , \mem0[124][3] ,
         \mem0[124][2] , \mem0[124][1] , \mem0[124][0] , \mem0[123][7] ,
         \mem0[123][6] , \mem0[123][5] , \mem0[123][4] , \mem0[123][3] ,
         \mem0[123][2] , \mem0[123][1] , \mem0[123][0] , \mem0[122][7] ,
         \mem0[122][6] , \mem0[122][5] , \mem0[122][4] , \mem0[122][3] ,
         \mem0[122][2] , \mem0[122][1] , \mem0[122][0] , \mem0[121][7] ,
         \mem0[121][6] , \mem0[121][5] , \mem0[121][4] , \mem0[121][3] ,
         \mem0[121][2] , \mem0[121][1] , \mem0[121][0] , \mem0[120][7] ,
         \mem0[120][6] , \mem0[120][5] , \mem0[120][4] , \mem0[120][3] ,
         \mem0[120][2] , \mem0[120][1] , \mem0[120][0] , \mem0[119][7] ,
         \mem0[119][6] , \mem0[119][5] , \mem0[119][4] , \mem0[119][3] ,
         \mem0[119][2] , \mem0[119][1] , \mem0[119][0] , \mem0[118][7] ,
         \mem0[118][6] , \mem0[118][5] , \mem0[118][4] , \mem0[118][3] ,
         \mem0[118][2] , \mem0[118][1] , \mem0[118][0] , \mem0[117][7] ,
         \mem0[117][6] , \mem0[117][5] , \mem0[117][4] , \mem0[117][3] ,
         \mem0[117][2] , \mem0[117][1] , \mem0[117][0] , \mem0[116][7] ,
         \mem0[116][6] , \mem0[116][5] , \mem0[116][4] , \mem0[116][3] ,
         \mem0[116][2] , \mem0[116][1] , \mem0[116][0] , \mem0[115][7] ,
         \mem0[115][6] , \mem0[115][5] , \mem0[115][4] , \mem0[115][3] ,
         \mem0[115][2] , \mem0[115][1] , \mem0[115][0] , \mem0[114][7] ,
         \mem0[114][6] , \mem0[114][5] , \mem0[114][4] , \mem0[114][3] ,
         \mem0[114][2] , \mem0[114][1] , \mem0[114][0] , \mem0[113][7] ,
         \mem0[113][6] , \mem0[113][5] , \mem0[113][4] , \mem0[113][3] ,
         \mem0[113][2] , \mem0[113][1] , \mem0[113][0] , \mem0[112][7] ,
         \mem0[112][6] , \mem0[112][5] , \mem0[112][4] , \mem0[112][3] ,
         \mem0[112][2] , \mem0[112][1] , \mem0[112][0] , \mem0[111][7] ,
         \mem0[111][6] , \mem0[111][5] , \mem0[111][4] , \mem0[111][3] ,
         \mem0[111][2] , \mem0[111][1] , \mem0[111][0] , \mem0[110][7] ,
         \mem0[110][6] , \mem0[110][5] , \mem0[110][4] , \mem0[110][3] ,
         \mem0[110][2] , \mem0[110][1] , \mem0[110][0] , \mem0[109][7] ,
         \mem0[109][6] , \mem0[109][5] , \mem0[109][4] , \mem0[109][3] ,
         \mem0[109][2] , \mem0[109][1] , \mem0[109][0] , \mem0[108][7] ,
         \mem0[108][6] , \mem0[108][5] , \mem0[108][4] , \mem0[108][3] ,
         \mem0[108][2] , \mem0[108][1] , \mem0[108][0] , \mem0[107][7] ,
         \mem0[107][6] , \mem0[107][5] , \mem0[107][4] , \mem0[107][3] ,
         \mem0[107][2] , \mem0[107][1] , \mem0[107][0] , \mem0[106][7] ,
         \mem0[106][6] , \mem0[106][5] , \mem0[106][4] , \mem0[106][3] ,
         \mem0[106][2] , \mem0[106][1] , \mem0[106][0] , \mem0[105][7] ,
         \mem0[105][6] , \mem0[105][5] , \mem0[105][4] , \mem0[105][3] ,
         \mem0[105][2] , \mem0[105][1] , \mem0[105][0] , \mem0[104][7] ,
         \mem0[104][6] , \mem0[104][5] , \mem0[104][4] , \mem0[104][3] ,
         \mem0[104][2] , \mem0[104][1] , \mem0[104][0] , \mem0[103][7] ,
         \mem0[103][6] , \mem0[103][5] , \mem0[103][4] , \mem0[103][3] ,
         \mem0[103][2] , \mem0[103][1] , \mem0[103][0] , \mem0[102][7] ,
         \mem0[102][6] , \mem0[102][5] , \mem0[102][4] , \mem0[102][3] ,
         \mem0[102][2] , \mem0[102][1] , \mem0[102][0] , \mem0[101][7] ,
         \mem0[101][6] , \mem0[101][5] , \mem0[101][4] , \mem0[101][3] ,
         \mem0[101][2] , \mem0[101][1] , \mem0[101][0] , \mem0[100][7] ,
         \mem0[100][6] , \mem0[100][5] , \mem0[100][4] , \mem0[100][3] ,
         \mem0[100][2] , \mem0[100][1] , \mem0[100][0] , \mem0[99][7] ,
         \mem0[99][6] , \mem0[99][5] , \mem0[99][4] , \mem0[99][3] ,
         \mem0[99][2] , \mem0[99][1] , \mem0[99][0] , \mem0[98][7] ,
         \mem0[98][6] , \mem0[98][5] , \mem0[98][4] , \mem0[98][3] ,
         \mem0[98][2] , \mem0[98][1] , \mem0[98][0] , \mem0[97][7] ,
         \mem0[97][6] , \mem0[97][5] , \mem0[97][4] , \mem0[97][3] ,
         \mem0[97][2] , \mem0[97][1] , \mem0[97][0] , \mem0[96][7] ,
         \mem0[96][6] , \mem0[96][5] , \mem0[96][4] , \mem0[96][3] ,
         \mem0[96][2] , \mem0[96][1] , \mem0[96][0] , \mem0[95][7] ,
         \mem0[95][6] , \mem0[95][5] , \mem0[95][4] , \mem0[95][3] ,
         \mem0[95][2] , \mem0[95][1] , \mem0[95][0] , \mem0[94][7] ,
         \mem0[94][6] , \mem0[94][5] , \mem0[94][4] , \mem0[94][3] ,
         \mem0[94][2] , \mem0[94][1] , \mem0[94][0] , \mem0[93][7] ,
         \mem0[93][6] , \mem0[93][5] , \mem0[93][4] , \mem0[93][3] ,
         \mem0[93][2] , \mem0[93][1] , \mem0[93][0] , \mem0[92][7] ,
         \mem0[92][6] , \mem0[92][5] , \mem0[92][4] , \mem0[92][3] ,
         \mem0[92][2] , \mem0[92][1] , \mem0[92][0] , \mem0[91][7] ,
         \mem0[91][6] , \mem0[91][5] , \mem0[91][4] , \mem0[91][3] ,
         \mem0[91][2] , \mem0[91][1] , \mem0[91][0] , \mem0[90][7] ,
         \mem0[90][6] , \mem0[90][5] , \mem0[90][4] , \mem0[90][3] ,
         \mem0[90][2] , \mem0[90][1] , \mem0[90][0] , \mem0[89][7] ,
         \mem0[89][6] , \mem0[89][5] , \mem0[89][4] , \mem0[89][3] ,
         \mem0[89][2] , \mem0[89][1] , \mem0[89][0] , \mem0[88][7] ,
         \mem0[88][6] , \mem0[88][5] , \mem0[88][4] , \mem0[88][3] ,
         \mem0[88][2] , \mem0[88][1] , \mem0[88][0] , \mem0[87][7] ,
         \mem0[87][6] , \mem0[87][5] , \mem0[87][4] , \mem0[87][3] ,
         \mem0[87][2] , \mem0[87][1] , \mem0[87][0] , \mem0[86][7] ,
         \mem0[86][6] , \mem0[86][5] , \mem0[86][4] , \mem0[86][3] ,
         \mem0[86][2] , \mem0[86][1] , \mem0[86][0] , \mem0[85][7] ,
         \mem0[85][6] , \mem0[85][5] , \mem0[85][4] , \mem0[85][3] ,
         \mem0[85][2] , \mem0[85][1] , \mem0[85][0] , \mem0[84][7] ,
         \mem0[84][6] , \mem0[84][5] , \mem0[84][4] , \mem0[84][3] ,
         \mem0[84][2] , \mem0[84][1] , \mem0[84][0] , \mem0[83][7] ,
         \mem0[83][6] , \mem0[83][5] , \mem0[83][4] , \mem0[83][3] ,
         \mem0[83][2] , \mem0[83][1] , \mem0[83][0] , \mem0[82][7] ,
         \mem0[82][6] , \mem0[82][5] , \mem0[82][4] , \mem0[82][3] ,
         \mem0[82][2] , \mem0[82][1] , \mem0[82][0] , \mem0[81][7] ,
         \mem0[81][6] , \mem0[81][5] , \mem0[81][4] , \mem0[81][3] ,
         \mem0[81][2] , \mem0[81][1] , \mem0[81][0] , \mem0[80][7] ,
         \mem0[80][6] , \mem0[80][5] , \mem0[80][4] , \mem0[80][3] ,
         \mem0[80][2] , \mem0[80][1] , \mem0[80][0] , \mem0[79][7] ,
         \mem0[79][6] , \mem0[79][5] , \mem0[79][4] , \mem0[79][3] ,
         \mem0[79][2] , \mem0[79][1] , \mem0[79][0] , \mem0[78][7] ,
         \mem0[78][6] , \mem0[78][5] , \mem0[78][4] , \mem0[78][3] ,
         \mem0[78][2] , \mem0[78][1] , \mem0[78][0] , \mem0[77][7] ,
         \mem0[77][6] , \mem0[77][5] , \mem0[77][4] , \mem0[77][3] ,
         \mem0[77][2] , \mem0[77][1] , \mem0[77][0] , \mem0[76][7] ,
         \mem0[76][6] , \mem0[76][5] , \mem0[76][4] , \mem0[76][3] ,
         \mem0[76][2] , \mem0[76][1] , \mem0[76][0] , \mem0[75][7] ,
         \mem0[75][6] , \mem0[75][5] , \mem0[75][4] , \mem0[75][3] ,
         \mem0[75][2] , \mem0[75][1] , \mem0[75][0] , \mem0[74][7] ,
         \mem0[74][6] , \mem0[74][5] , \mem0[74][4] , \mem0[74][3] ,
         \mem0[74][2] , \mem0[74][1] , \mem0[74][0] , \mem0[73][7] ,
         \mem0[73][6] , \mem0[73][5] , \mem0[73][4] , \mem0[73][3] ,
         \mem0[73][2] , \mem0[73][1] , \mem0[73][0] , \mem0[72][7] ,
         \mem0[72][6] , \mem0[72][5] , \mem0[72][4] , \mem0[72][3] ,
         \mem0[72][2] , \mem0[72][1] , \mem0[72][0] , \mem0[71][7] ,
         \mem0[71][6] , \mem0[71][5] , \mem0[71][4] , \mem0[71][3] ,
         \mem0[71][2] , \mem0[71][1] , \mem0[71][0] , \mem0[70][7] ,
         \mem0[70][6] , \mem0[70][5] , \mem0[70][4] , \mem0[70][3] ,
         \mem0[70][2] , \mem0[70][1] , \mem0[70][0] , \mem0[69][7] ,
         \mem0[69][6] , \mem0[69][5] , \mem0[69][4] , \mem0[69][3] ,
         \mem0[69][2] , \mem0[69][1] , \mem0[69][0] , \mem0[68][7] ,
         \mem0[68][6] , \mem0[68][5] , \mem0[68][4] , \mem0[68][3] ,
         \mem0[68][2] , \mem0[68][1] , \mem0[68][0] , \mem0[67][7] ,
         \mem0[67][6] , \mem0[67][5] , \mem0[67][4] , \mem0[67][3] ,
         \mem0[67][2] , \mem0[67][1] , \mem0[67][0] , \mem0[66][7] ,
         \mem0[66][6] , \mem0[66][5] , \mem0[66][4] , \mem0[66][3] ,
         \mem0[66][2] , \mem0[66][1] , \mem0[66][0] , \mem0[65][7] ,
         \mem0[65][6] , \mem0[65][5] , \mem0[65][4] , \mem0[65][3] ,
         \mem0[65][2] , \mem0[65][1] , \mem0[65][0] , \mem0[64][7] ,
         \mem0[64][6] , \mem0[64][5] , \mem0[64][4] , \mem0[64][3] ,
         \mem0[64][2] , \mem0[64][1] , \mem0[64][0] , \mem0[63][7] ,
         \mem0[63][6] , \mem0[63][5] , \mem0[63][4] , \mem0[63][3] ,
         \mem0[63][2] , \mem0[63][1] , \mem0[63][0] , \mem0[62][7] ,
         \mem0[62][6] , \mem0[62][5] , \mem0[62][4] , \mem0[62][3] ,
         \mem0[62][2] , \mem0[62][1] , \mem0[62][0] , \mem0[61][7] ,
         \mem0[61][6] , \mem0[61][5] , \mem0[61][4] , \mem0[61][3] ,
         \mem0[61][2] , \mem0[61][1] , \mem0[61][0] , \mem0[60][7] ,
         \mem0[60][6] , \mem0[60][5] , \mem0[60][4] , \mem0[60][3] ,
         \mem0[60][2] , \mem0[60][1] , \mem0[60][0] , \mem0[59][7] ,
         \mem0[59][6] , \mem0[59][5] , \mem0[59][4] , \mem0[59][3] ,
         \mem0[59][2] , \mem0[59][1] , \mem0[59][0] , \mem0[58][7] ,
         \mem0[58][6] , \mem0[58][5] , \mem0[58][4] , \mem0[58][3] ,
         \mem0[58][2] , \mem0[58][1] , \mem0[58][0] , \mem0[57][7] ,
         \mem0[57][6] , \mem0[57][5] , \mem0[57][4] , \mem0[57][3] ,
         \mem0[57][2] , \mem0[57][1] , \mem0[57][0] , \mem0[56][7] ,
         \mem0[56][6] , \mem0[56][5] , \mem0[56][4] , \mem0[56][3] ,
         \mem0[56][2] , \mem0[56][1] , \mem0[56][0] , \mem0[55][7] ,
         \mem0[55][6] , \mem0[55][5] , \mem0[55][4] , \mem0[55][3] ,
         \mem0[55][2] , \mem0[55][1] , \mem0[55][0] , \mem0[54][7] ,
         \mem0[54][6] , \mem0[54][5] , \mem0[54][4] , \mem0[54][3] ,
         \mem0[54][2] , \mem0[54][1] , \mem0[54][0] , \mem0[53][7] ,
         \mem0[53][6] , \mem0[53][5] , \mem0[53][4] , \mem0[53][3] ,
         \mem0[53][2] , \mem0[53][1] , \mem0[53][0] , \mem0[52][7] ,
         \mem0[52][6] , \mem0[52][5] , \mem0[52][4] , \mem0[52][3] ,
         \mem0[52][2] , \mem0[52][1] , \mem0[52][0] , \mem0[51][7] ,
         \mem0[51][6] , \mem0[51][5] , \mem0[51][4] , \mem0[51][3] ,
         \mem0[51][2] , \mem0[51][1] , \mem0[51][0] , \mem0[50][7] ,
         \mem0[50][6] , \mem0[50][5] , \mem0[50][4] , \mem0[50][3] ,
         \mem0[50][2] , \mem0[50][1] , \mem0[50][0] , \mem0[49][7] ,
         \mem0[49][6] , \mem0[49][5] , \mem0[49][4] , \mem0[49][3] ,
         \mem0[49][2] , \mem0[49][1] , \mem0[49][0] , \mem0[48][7] ,
         \mem0[48][6] , \mem0[48][5] , \mem0[48][4] , \mem0[48][3] ,
         \mem0[48][2] , \mem0[48][1] , \mem0[48][0] , \mem0[47][7] ,
         \mem0[47][6] , \mem0[47][5] , \mem0[47][4] , \mem0[47][3] ,
         \mem0[47][2] , \mem0[47][1] , \mem0[47][0] , \mem0[46][7] ,
         \mem0[46][6] , \mem0[46][5] , \mem0[46][4] , \mem0[46][3] ,
         \mem0[46][2] , \mem0[46][1] , \mem0[46][0] , \mem0[45][7] ,
         \mem0[45][6] , \mem0[45][5] , \mem0[45][4] , \mem0[45][3] ,
         \mem0[45][2] , \mem0[45][1] , \mem0[45][0] , \mem0[44][7] ,
         \mem0[44][6] , \mem0[44][5] , \mem0[44][4] , \mem0[44][3] ,
         \mem0[44][2] , \mem0[44][1] , \mem0[44][0] , \mem0[43][7] ,
         \mem0[43][6] , \mem0[43][5] , \mem0[43][4] , \mem0[43][3] ,
         \mem0[43][2] , \mem0[43][1] , \mem0[43][0] , \mem0[42][7] ,
         \mem0[42][6] , \mem0[42][5] , \mem0[42][4] , \mem0[42][3] ,
         \mem0[42][2] , \mem0[42][1] , \mem0[42][0] , \mem0[41][7] ,
         \mem0[41][6] , \mem0[41][5] , \mem0[41][4] , \mem0[41][3] ,
         \mem0[41][2] , \mem0[41][1] , \mem0[41][0] , \mem0[40][7] ,
         \mem0[40][6] , \mem0[40][5] , \mem0[40][4] , \mem0[40][3] ,
         \mem0[40][2] , \mem0[40][1] , \mem0[40][0] , \mem0[39][7] ,
         \mem0[39][6] , \mem0[39][5] , \mem0[39][4] , \mem0[39][3] ,
         \mem0[39][2] , \mem0[39][1] , \mem0[39][0] , \mem0[38][7] ,
         \mem0[38][6] , \mem0[38][5] , \mem0[38][4] , \mem0[38][3] ,
         \mem0[38][2] , \mem0[38][1] , \mem0[38][0] , \mem0[37][7] ,
         \mem0[37][6] , \mem0[37][5] , \mem0[37][4] , \mem0[37][3] ,
         \mem0[37][2] , \mem0[37][1] , \mem0[37][0] , \mem0[36][7] ,
         \mem0[36][6] , \mem0[36][5] , \mem0[36][4] , \mem0[36][3] ,
         \mem0[36][2] , \mem0[36][1] , \mem0[36][0] , \mem0[35][7] ,
         \mem0[35][6] , \mem0[35][5] , \mem0[35][4] , \mem0[35][3] ,
         \mem0[35][2] , \mem0[35][1] , \mem0[35][0] , \mem0[34][7] ,
         \mem0[34][6] , \mem0[34][5] , \mem0[34][4] , \mem0[34][3] ,
         \mem0[34][2] , \mem0[34][1] , \mem0[34][0] , \mem0[33][7] ,
         \mem0[33][6] , \mem0[33][5] , \mem0[33][4] , \mem0[33][3] ,
         \mem0[33][2] , \mem0[33][1] , \mem0[33][0] , \mem0[32][7] ,
         \mem0[32][6] , \mem0[32][5] , \mem0[32][4] , \mem0[32][3] ,
         \mem0[32][2] , \mem0[32][1] , \mem0[32][0] , \mem0[31][7] ,
         \mem0[31][6] , \mem0[31][5] , \mem0[31][4] , \mem0[31][3] ,
         \mem0[31][2] , \mem0[31][1] , \mem0[31][0] , \mem0[30][7] ,
         \mem0[30][6] , \mem0[30][5] , \mem0[30][4] , \mem0[30][3] ,
         \mem0[30][2] , \mem0[30][1] , \mem0[30][0] , \mem0[29][7] ,
         \mem0[29][6] , \mem0[29][5] , \mem0[29][4] , \mem0[29][3] ,
         \mem0[29][2] , \mem0[29][1] , \mem0[29][0] , \mem0[28][7] ,
         \mem0[28][6] , \mem0[28][5] , \mem0[28][4] , \mem0[28][3] ,
         \mem0[28][2] , \mem0[28][1] , \mem0[28][0] , \mem0[27][7] ,
         \mem0[27][6] , \mem0[27][5] , \mem0[27][4] , \mem0[27][3] ,
         \mem0[27][2] , \mem0[27][1] , \mem0[27][0] , \mem0[26][7] ,
         \mem0[26][6] , \mem0[26][5] , \mem0[26][4] , \mem0[26][3] ,
         \mem0[26][2] , \mem0[26][1] , \mem0[26][0] , \mem0[25][7] ,
         \mem0[25][6] , \mem0[25][5] , \mem0[25][4] , \mem0[25][3] ,
         \mem0[25][2] , \mem0[25][1] , \mem0[25][0] , \mem0[24][7] ,
         \mem0[24][6] , \mem0[24][5] , \mem0[24][4] , \mem0[24][3] ,
         \mem0[24][2] , \mem0[24][1] , \mem0[24][0] , \mem0[23][7] ,
         \mem0[23][6] , \mem0[23][5] , \mem0[23][4] , \mem0[23][3] ,
         \mem0[23][2] , \mem0[23][1] , \mem0[23][0] , \mem0[22][7] ,
         \mem0[22][6] , \mem0[22][5] , \mem0[22][4] , \mem0[22][3] ,
         \mem0[22][2] , \mem0[22][1] , \mem0[22][0] , \mem0[21][7] ,
         \mem0[21][6] , \mem0[21][5] , \mem0[21][4] , \mem0[21][3] ,
         \mem0[21][2] , \mem0[21][1] , \mem0[21][0] , \mem0[20][7] ,
         \mem0[20][6] , \mem0[20][5] , \mem0[20][4] , \mem0[20][3] ,
         \mem0[20][2] , \mem0[20][1] , \mem0[20][0] , \mem0[19][7] ,
         \mem0[19][6] , \mem0[19][5] , \mem0[19][4] , \mem0[19][3] ,
         \mem0[19][2] , \mem0[19][1] , \mem0[19][0] , \mem0[18][7] ,
         \mem0[18][6] , \mem0[18][5] , \mem0[18][4] , \mem0[18][3] ,
         \mem0[18][2] , \mem0[18][1] , \mem0[18][0] , \mem0[17][7] ,
         \mem0[17][6] , \mem0[17][5] , \mem0[17][4] , \mem0[17][3] ,
         \mem0[17][2] , \mem0[17][1] , \mem0[17][0] , \mem0[16][7] ,
         \mem0[16][6] , \mem0[16][5] , \mem0[16][4] , \mem0[16][3] ,
         \mem0[16][2] , \mem0[16][1] , \mem0[16][0] , \mem0[15][7] ,
         \mem0[15][6] , \mem0[15][5] , \mem0[15][4] , \mem0[15][3] ,
         \mem0[15][2] , \mem0[15][1] , \mem0[15][0] , \mem0[14][7] ,
         \mem0[14][6] , \mem0[14][5] , \mem0[14][4] , \mem0[14][3] ,
         \mem0[14][2] , \mem0[14][1] , \mem0[14][0] , \mem0[13][7] ,
         \mem0[13][6] , \mem0[13][5] , \mem0[13][4] , \mem0[13][3] ,
         \mem0[13][2] , \mem0[13][1] , \mem0[13][0] , \mem0[12][7] ,
         \mem0[12][6] , \mem0[12][5] , \mem0[12][4] , \mem0[12][3] ,
         \mem0[12][2] , \mem0[12][1] , \mem0[12][0] , \mem0[11][7] ,
         \mem0[11][6] , \mem0[11][5] , \mem0[11][4] , \mem0[11][3] ,
         \mem0[11][2] , \mem0[11][1] , \mem0[11][0] , \mem0[10][7] ,
         \mem0[10][6] , \mem0[10][5] , \mem0[10][4] , \mem0[10][3] ,
         \mem0[10][2] , \mem0[10][1] , \mem0[10][0] , \mem0[9][7] ,
         \mem0[9][6] , \mem0[9][5] , \mem0[9][4] , \mem0[9][3] , \mem0[9][2] ,
         \mem0[9][1] , \mem0[9][0] , \mem0[8][7] , \mem0[8][6] , \mem0[8][5] ,
         \mem0[8][4] , \mem0[8][3] , \mem0[8][2] , \mem0[8][1] , \mem0[8][0] ,
         \mem0[7][7] , \mem0[7][6] , \mem0[7][5] , \mem0[7][4] , \mem0[7][3] ,
         \mem0[7][2] , \mem0[7][1] , \mem0[7][0] , \mem0[6][7] , \mem0[6][6] ,
         \mem0[6][5] , \mem0[6][4] , \mem0[6][3] , \mem0[6][2] , \mem0[6][1] ,
         \mem0[6][0] , \mem0[5][7] , \mem0[5][6] , \mem0[5][5] , \mem0[5][4] ,
         \mem0[5][3] , \mem0[5][2] , \mem0[5][1] , \mem0[5][0] , \mem0[4][7] ,
         \mem0[4][6] , \mem0[4][5] , \mem0[4][4] , \mem0[4][3] , \mem0[4][2] ,
         \mem0[4][1] , \mem0[4][0] , \mem0[3][7] , \mem0[3][6] , \mem0[3][5] ,
         \mem0[3][4] , \mem0[3][3] , \mem0[3][2] , \mem0[3][1] , \mem0[3][0] ,
         \mem0[2][7] , \mem0[2][6] , \mem0[2][5] , \mem0[2][4] , \mem0[2][3] ,
         \mem0[2][2] , \mem0[2][1] , \mem0[2][0] , \mem0[1][7] , \mem0[1][6] ,
         \mem0[1][5] , \mem0[1][4] , \mem0[1][3] , \mem0[1][2] , \mem0[1][1] ,
         \mem0[1][0] , \mem0[0][7] , \mem0[0][6] , \mem0[0][5] , \mem0[0][4] ,
         \mem0[0][3] , \mem0[0][2] , \mem0[0][1] , \mem0[0][0] , n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n10397, n10399, n10401, n10403, n10405, n10407, n10409, n10411,
         n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419,
         n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427,
         n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435,
         n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443,
         n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451,
         n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459,
         n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467,
         n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475,
         n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483,
         n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491,
         n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499,
         n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507,
         n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515,
         n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523,
         n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531,
         n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539,
         n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547,
         n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555,
         n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563,
         n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571,
         n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579,
         n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587,
         n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595,
         n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603,
         n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611,
         n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619,
         n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627,
         n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635,
         n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643,
         n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651,
         n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659,
         n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667,
         n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675,
         n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683,
         n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691,
         n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699,
         n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707,
         n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715,
         n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723,
         n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731,
         n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739,
         n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747,
         n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755,
         n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763,
         n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771,
         n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779,
         n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787,
         n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795,
         n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803,
         n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811,
         n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819,
         n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827,
         n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835,
         n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843,
         n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851,
         n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859,
         n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867,
         n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875,
         n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883,
         n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891,
         n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899,
         n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907,
         n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915,
         n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923,
         n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931,
         n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939,
         n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947,
         n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955,
         n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963,
         n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971,
         n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979,
         n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987,
         n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995,
         n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003,
         n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011,
         n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019,
         n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027,
         n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035,
         n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043,
         n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051,
         n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059,
         n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067,
         n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075,
         n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083,
         n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091,
         n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099,
         n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107,
         n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115,
         n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123,
         n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131,
         n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139,
         n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147,
         n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155,
         n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163,
         n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171,
         n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179,
         n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187,
         n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195,
         n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203,
         n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211,
         n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219,
         n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227,
         n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235,
         n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243,
         n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251,
         n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259,
         n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267,
         n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275,
         n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283,
         n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291,
         n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299,
         n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307,
         n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315,
         n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323,
         n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331,
         n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339,
         n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347,
         n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355,
         n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363,
         n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371,
         n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379,
         n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387,
         n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395,
         n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403,
         n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411,
         n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419,
         n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427,
         n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435,
         n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443,
         n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451,
         n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459,
         n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467,
         n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475,
         n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483,
         n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491,
         n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499,
         n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507,
         n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515,
         n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523,
         n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531,
         n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539,
         n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547,
         n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555,
         n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563,
         n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571,
         n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579,
         n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587,
         n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595,
         n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603,
         n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611,
         n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619,
         n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627,
         n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635,
         n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643,
         n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651,
         n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659,
         n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667,
         n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675,
         n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683,
         n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691,
         n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699,
         n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707,
         n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715,
         n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723,
         n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731,
         n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739,
         n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747,
         n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755,
         n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763,
         n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771,
         n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779,
         n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787,
         n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795,
         n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803,
         n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811,
         n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819,
         n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827,
         n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835,
         n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843,
         n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851,
         n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859,
         n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867,
         n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875,
         n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883,
         n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891,
         n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899,
         n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907,
         n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915,
         n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923,
         n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931,
         n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939,
         n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947,
         n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955,
         n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963,
         n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971,
         n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979,
         n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987,
         n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995,
         n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003,
         n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011,
         n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019,
         n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027,
         n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035,
         n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043,
         n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051,
         n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059,
         n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067,
         n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075,
         n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083,
         n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091,
         n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099,
         n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107,
         n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115,
         n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123,
         n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131,
         n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139,
         n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147,
         n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155,
         n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163,
         n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171,
         n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179,
         n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187,
         n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195,
         n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203,
         n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211,
         n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219,
         n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227,
         n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235,
         n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243,
         n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251,
         n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259,
         n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267,
         n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275,
         n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283,
         n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291,
         n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299,
         n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307,
         n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315,
         n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323,
         n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331,
         n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339,
         n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347,
         n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355,
         n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363,
         n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371,
         n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379,
         n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387,
         n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395,
         n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403,
         n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411,
         n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419,
         n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427,
         n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435,
         n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443,
         n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451,
         n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459,
         n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467,
         n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475,
         n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483,
         n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491,
         n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499,
         n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507,
         n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515,
         n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523,
         n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531,
         n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539,
         n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547,
         n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555,
         n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563,
         n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571,
         n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579,
         n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587,
         n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595,
         n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603,
         n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611,
         n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619,
         n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627,
         n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635,
         n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643,
         n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651,
         n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659,
         n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667,
         n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675,
         n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683,
         n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691,
         n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699,
         n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707,
         n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715,
         n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723,
         n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731,
         n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739,
         n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747,
         n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755,
         n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763,
         n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771,
         n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779,
         n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787,
         n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795,
         n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803,
         n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811,
         n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819,
         n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827,
         n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835,
         n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843,
         n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851,
         n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859,
         n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867,
         n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875,
         n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883,
         n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891,
         n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899,
         n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907,
         n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915,
         n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923,
         n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931,
         n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939,
         n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947,
         n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955,
         n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963,
         n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971,
         n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979,
         n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987,
         n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995,
         n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003,
         n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011,
         n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019,
         n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027,
         n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035,
         n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043,
         n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051,
         n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059,
         n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067,
         n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075,
         n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083,
         n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091,
         n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099,
         n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107,
         n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115,
         n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123,
         n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131,
         n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139,
         n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147,
         n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155,
         n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163,
         n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171,
         n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179,
         n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187,
         n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195,
         n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203,
         n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211,
         n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219,
         n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227,
         n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235,
         n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243,
         n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251,
         n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259,
         n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267,
         n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275,
         n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283,
         n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291,
         n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299,
         n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307,
         n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315,
         n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323,
         n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331,
         n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339,
         n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347,
         n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355,
         n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363,
         n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371,
         n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379,
         n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387,
         n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395,
         n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403,
         n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411,
         n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419,
         n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427,
         n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435,
         n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443,
         n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451,
         n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459,
         n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467,
         n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475,
         n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483,
         n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491,
         n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499,
         n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507,
         n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515,
         n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523,
         n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531,
         n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539,
         n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547,
         n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555,
         n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563,
         n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571,
         n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579,
         n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587,
         n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595,
         n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603,
         n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611,
         n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619,
         n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627,
         n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635,
         n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643,
         n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651,
         n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659,
         n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667,
         n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675,
         n13676, n13677, n13678, n13679, n13680, n13681, n13682, n13683,
         n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691,
         n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699,
         n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707,
         n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715,
         n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723,
         n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731,
         n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739,
         n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747,
         n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755,
         n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763,
         n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771,
         n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779,
         n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787,
         n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795,
         n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803,
         n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811,
         n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819,
         n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827,
         n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835,
         n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843,
         n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851,
         n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859,
         n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867,
         n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875,
         n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883,
         n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891,
         n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899,
         n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907,
         n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915,
         n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923,
         n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931,
         n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939,
         n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947,
         n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955,
         n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963,
         n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971,
         n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979,
         n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987,
         n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995,
         n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003,
         n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011,
         n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019,
         n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027,
         n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035,
         n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043,
         n14044, n14045, n14046, n14047, n14048, n14049, n14050, n14051,
         n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059,
         n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067,
         n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075,
         n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083,
         n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091,
         n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099,
         n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107,
         n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115,
         n14116, n14117, n14118, n14119, n14120, n14121, n14122, n14123,
         n14124, n14125, n14126, n14127, n14128, n14129, n14130, n14131,
         n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139,
         n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14147,
         n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155,
         n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163,
         n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171,
         n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179,
         n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187,
         n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195,
         n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203,
         n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211,
         n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219,
         n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227,
         n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235,
         n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243,
         n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251,
         n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259,
         n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267,
         n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275,
         n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283,
         n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291,
         n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299,
         n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307,
         n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315,
         n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323,
         n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331,
         n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339,
         n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347,
         n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355,
         n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363,
         n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371,
         n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379,
         n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387,
         n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395,
         n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403,
         n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411,
         n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419,
         n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427,
         n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435,
         n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443,
         n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451,
         n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459,
         n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467,
         n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475,
         n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483,
         n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491,
         n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499,
         n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507,
         n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515,
         n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523,
         n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531,
         n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539,
         n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547,
         n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555,
         n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563,
         n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571,
         n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579,
         n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587,
         n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595,
         n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603,
         n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611,
         n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619,
         n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627,
         n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635,
         n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643,
         n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651,
         n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659,
         n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667,
         n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675,
         n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683,
         n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691,
         n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699,
         n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707,
         n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715,
         n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723,
         n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731,
         n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739,
         n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747,
         n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755,
         n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763,
         n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771,
         n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779,
         n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787,
         n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795,
         n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803,
         n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811,
         n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819,
         n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827,
         n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835,
         n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843,
         n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851,
         n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859,
         n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867,
         n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875,
         n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883,
         n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891,
         n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899,
         n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907,
         n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915,
         n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923,
         n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931,
         n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939,
         n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947,
         n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955,
         n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963,
         n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971,
         n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979,
         n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987,
         n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995,
         n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003,
         n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011,
         n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019,
         n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027,
         n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035,
         n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043,
         n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051,
         n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059,
         n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067,
         n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075,
         n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083,
         n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091,
         n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099,
         n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107,
         n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115,
         n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123,
         n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131,
         n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139,
         n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147,
         n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155,
         n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163,
         n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171,
         n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179,
         n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187,
         n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195,
         n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203,
         n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211,
         n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219,
         n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227,
         n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235,
         n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243,
         n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251,
         n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259,
         n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267,
         n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275,
         n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283,
         n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291,
         n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299,
         n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307,
         n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315,
         n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323,
         n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331,
         n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339,
         n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347,
         n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355,
         n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363,
         n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371,
         n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379,
         n15380, n15381, n15382, n15383, n15384, n15385, n15386, n15387,
         n15388, n15389, n15390, n15391, n15392, n15393, n15394, n15395,
         n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403,
         n15404, n15405, n15406, n15407, n15408, n15409, n15410, n15411,
         n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419,
         n15420, n15421, n15422, n15423, n15424, n15425, n15426, n15427,
         n15428, n15429, n15430, n15431, n15432, n15433, n15434, n15435,
         n15436, n15437, n15438, n15439, n15440, n15441, n15442, n15443,
         n15444, n15445, n15446, n15447, n15448, n15449, n15450, n15451,
         n15452, n15453, n15454, n15455, n15456, n15457, n15458, n15459,
         n15460, n15461, n15462, n15463, n15464, n15465, n15466, n15467,
         n15468, n15469, n15470, n15471, n15472, n15473, n15474, n15475,
         n15476, n15477, n15478, n15479, n15480, n15481, n15482, n15483,
         n15484, n15485, n15486, n15487, n15488, n15489, n15490, n15491,
         n15492, n15493, n15494, n15495, n15496, n15497, n15498, n15499,
         n15500, n15501, n15502, n15503, n15504, n15505, n15506, n15507,
         n15508, n15509, n15510, n15511, n15512, n15513, n15514, n15515,
         n15516, n15517, n15518, n15519, n15520, n15521, n15522, n15523,
         n15524, n15525, n15526, n15527, n15528, n15529, n15530, n15531,
         n15532, n15533, n15534, n15535, n15536, n15537, n15538, n15539,
         n15540, n15541, n15542, n15543, n15544, n15545, n15546, n15547,
         n15548, n15549, n15550, n15551, n15552, n15553, n15554, n15555,
         n15556, n15557, n15558, n15559, n15560, n15561, n15562, n15563,
         n15564, n15565, n15566, n15567, n15568, n15569, n15570, n15571,
         n15572, n15573, n15574, n15575, n15576, n15577, n15578, n15579,
         n15580, n15581, n15582, n15583, n15584, n15585, n15586, n15587,
         n15588, n15589, n15590, n15591, n15592, n15593, n15594, n15595,
         n15596, n15597, n15598, n15599, n15600, n15601, n15602, n15603,
         n15604, n15605, n15606, n15607, n15608, n15609, n15610, n15611,
         n15612, n15613, n15614, n15615, n15616, n15617, n15618, n15619,
         n15620, n15621, n15622, n15623, n15624, n15625, n15626, n15627,
         n15628, n15629, n15630, n15631, n15632, n15633, n15634, n15635,
         n15636, n15637, n15638, n15639, n15640, n15641, n15642, n15643,
         n15644, n15645, n15646, n15647, n15648, n15649, n15650, n15651,
         n15652, n15653, n15654, n15655, n15656, n15657, n15658, n15659,
         n15660, n15661, n15662, n15663, n15664, n15665, n15666, n15667,
         n15668, n15669, n15670, n15671, n15672, n15673, n15674, n15675,
         n15676, n15677, n15678, n15679, n15680, n15681, n15682, n15683,
         n15684, n15685, n15686, n15687, n15688, n15689, n15690, n15691,
         n15692, n15693, n15694, n15695, n15696, n15697, n15698, n15699,
         n15700, n15701, n15702, n15703, n15704, n15705, n15706, n15707,
         n15708, n15709, n15710, n15711, n15712, n15713, n15714, n15715,
         n15716, n15717, n15718, n15719, n15720, n15721, n15722, n15723,
         n15724, n15725, n15726, n15727, n15728, n15729, n15730, n15731,
         n15732, n15733, n15734, n15735, n15736, n15737, n15738, n15739,
         n15740, n15741, n15742, n15743, n15744, n15745, n15746, n15747,
         n15748, n15749, n15750, n15751, n15752, n15753, n15754, n15755,
         n15756, n15757, n15758, n15759, n15760, n15761, n15762, n15763,
         n15764, n15765, n15766, n15767, n15768, n15769, n15770, n15771,
         n15772, n15773, n15774, n15775, n15776, n15777, n15778, n15779,
         n15780, n15781, n15782, n15783, n15784, n15785, n15786, n15787,
         n15788, n15789, n15790, n15791, n15792, n15793, n15794, n15795,
         n15796, n15797, n15798, n15799, n15800, n15801, n15802, n15803,
         n15804, n15805, n15806, n15807, n15808, n15809, n15810, n15811,
         n15812, n15813, n15814, n15815, n15816, n15817, n15818, n15819,
         n15820, n15821, n15822, n15823, n15824, n15825, n15826, n15827,
         n15828, n15829, n15830, n15831, n15832, n15833, n15834, n15835,
         n15836, n15837, n15838, n15839, n15840, n15841, n15842, n15843,
         n15844, n15845, n15846, n15847, n15848, n15849, n15850, n15851,
         n15852, n15853, n15854, n15855, n15856, n15857, n15858, n15859,
         n15860, n15861, n15862, n15863, n15864, n15865, n15866, n15867,
         n15868, n15869, n15870, n15871, n15872, n15873, n15874, n15875,
         n15876, n15877, n15878, n15879, n15880, n15881, n15882, n15883,
         n15884, n15885, n15886, n15887, n15888, n15889, n15890, n15891,
         n15892, n15893, n15894, n15895, n15896, n15897, n15898, n15899,
         n15900, n15901, n15902, n15903, n15904, n15905, n15906, n15907,
         n15908, n15909, n15910, n15911, n15912, n15913, n15914, n15915,
         n15916, n15917, n15918, n15919, n15920, n15921, n15922, n15923,
         n15924, n15925, n15926, n15927, n15928, n15929, n15930, n15931,
         n15932, n15933, n15934, n15935, n15936, n15937, n15938, n15939,
         n15940, n15941, n15942, n15943, n15944, n15945, n15946, n15947,
         n15948, n15949, n15950, n15951, n15952, n15953, n15954, n15955,
         n15956, n15957, n15958, n15959, n15960, n15961, n15962, n15963,
         n15964, n15965, n15966, n15967, n15968, n15969, n15970, n15971,
         n15972, n15973, n15974, n15975, n15976, n15977, n15978, n15979,
         n15980, n15981, n15982, n15983, n15984, n15985, n15986, n15987,
         n15988, n15989, n15990, n15991, n15992, n15993, n15994, n15995,
         n15996, n15997, n15998, n15999, n16000, n16001, n16002, n16003,
         n16004, n16005, n16006, n16007, n16008, n16009, n16010, n16011,
         n16012, n16013, n16014, n16015, n16016, n16017, n16018, n16019,
         n16020, n16021, n16022, n16023, n16024, n16025, n16026, n16027,
         n16028, n16029, n16030, n16031, n16032, n16033, n16034, n16035,
         n16036, n16037, n16038, n16039, n16040, n16041, n16042, n16043,
         n16044, n16045, n16046, n16047, n16048, n16049, n16050, n16051,
         n16052, n16053, n16054, n16055, n16056, n16057, n16058, n16059,
         n16060, n16061, n16062, n16063, n16064, n16065, n16066, n16067,
         n16068, n16069, n16070, n16071, n16072, n16073, n16074, n16075,
         n16076, n16077, n16078, n16079, n16080, n16081, n16082, n16083,
         n16084, n16085, n16086, n16087, n16088, n16089, n16090, n16091,
         n16092, n16093, n16094, n16095, n16096, n16097, n16098, n16099,
         n16100, n16101, n16102, n16103, n16104, n16105, n16106, n16107,
         n16108, n16109, n16110, n16111, n16112, n16113, n16114, n16115,
         n16116, n16117, n16118, n16119, n16120, n16121, n16122, n16123,
         n16124, n16125, n16126, n16127, n16128, n16129, n16130, n16131,
         n16132, n16133, n16134, n16135, n16136, n16137, n16138, n16139,
         n16140, n16141, n16142, n16143, n16144, n16145, n16146, n16147,
         n16148, n16149, n16150, n16151, n16152, n16153, n16154, n16155,
         n16156, n16157, n16158, n16159, n16160, n16161, n16162, n16163,
         n16164, n16165, n16166, n16167, n16168, n16169, n16170, n16171,
         n16172, n16173, n16174, n16175, n16176, n16177, n16178, n16179,
         n16180, n16181, n16182, n16183, n16184, n16185, n16186, n16187,
         n16188, n16189, n16190, n16191, n16192, n16193, n16194, n16195,
         n16196, n16197, n16198, n16199, n16200, n16201, n16202, n16203,
         n16204, n16205, n16206, n16207, n16208, n16209, n16210, n16211,
         n16212, n16213, n16214, n16215, n16216, n16217, n16218, n16219,
         n16220, n16221, n16222, n16223, n16224, n16225, n16226, n16227,
         n16228, n16229, n16230, n16231, n16232, n16233, n16234, n16235,
         n16236, n16237, n16238, n16239, n16240, n16241, n16242, n16243,
         n16244, n16245, n16246, n16247, n16248, n16249, n16250, n16251,
         n16252, n16253, n16254, n16255, n16256, n16257, n16258, n16259,
         n16260, n16261, n16262, n16263, n16264, n16265, n16266, n16267,
         n16268, n16269, n16270, n16271, n16272, n16273, n16274, n16275,
         n16276, n16277, n16278, n16279, n16280, n16281, n16282, n16283,
         n16284, n16285, n16286, n16287, n16288, n16289, n16290, n16291,
         n16292, n16293, n16294, n16295, n16296, n16297, n16298, n16299,
         n16300, n16301, n16302, n16303, n16304, n16305, n16306, n16307,
         n16308, n16309, n16310, n16311, n16312, n16313, n16314, n16315,
         n16316, n16317, n16318, n16319, n16320, n16321, n16322, n16323,
         n16324, n16325, n16326, n16327, n16328, n16329, n16330, n16331,
         n16332, n16333, n16334, n16335, n16336, n16337, n16338, n16339,
         n16340, n16341, n16342, n16343, n16344, n16345, n16346, n16347,
         n16348, n16349, n16350, n16351, n16352, n16353, n16354, n16355,
         n16356, n16357, n16358, n16359, n16360, n16361, n16362, n16363,
         n16364, n16365, n16366, n16367, n16368, n16369, n16370, n16371,
         n16372, n16373, n16374, n16375, n16376, n16377, n16378, n16379,
         n16380, n16381, n16382, n16383, n16384, n16385, n16386, n16387,
         n16388, n16389, n16390, n16391, n16392, n16393, n16394, n16395,
         n16396, n16397, n16398, n16399, n16400, n16401, n16402, n16403,
         n16404, n16405, n16406, n16407, n16408, n16409, n16410, n16411,
         n16412, n16413, n16414, n16415, n16416, n16417, n16418, n16419,
         n16420, n16421, n16422, n16423, n16424, n16425, n16426, n16427,
         n16428, n16429, n16430, n16431, n16432, n16433, n16434, n16435,
         n16436, n16437, n16438, n16439, n16440, n16441, n16442, n16443,
         n16444, n16445, n16446, n16447, n16448, n16449, n16450, n16451,
         n16452, n16453, n16454, n16455, n16456, n16457, n16458, n16459,
         n16460, n16461, n16462, n16463, n16464, n16465, n16466, n16467,
         n16468, n16469, n16470, n16471, n16472, n16473, n16474, n16475,
         n16476, n16477, n16478, n16479, n16480, n16481, n16482, n16483,
         n16484, n16485, n16486, n16487, n16488, n16489, n16490, n16491,
         n16492, n16493, n16494, n16495, n16496, n16497, n16498, n16499,
         n16500, n16501, n16502, n16503, n16504, n16505, n16506, n16507,
         n16508, n16509, n16510, n16511, n16512, n16513, n16514, n16515,
         n16516, n16517, n16518, n16519, n16520, n16521, n16522, n16523,
         n16524, n16525, n16526, n16527, n16528, n16529, n16530, n16531,
         n16532, n16533, n16534, n16535, n16536, n16537, n16538, n16539,
         n16540, n16541, n16542, n16543, n16544, n16545, n16546, n16547,
         n16548, n16549, n16550, n16551, n16552, n16553, n16554, n16555,
         n16556, n16557, n16558, n16559, n16560, n16561, n16562, n16563,
         n16564, n16565, n16566, n16567, n16568, n16569, n16570, n16571,
         n16572, n16573, n16574, n16575, n16576, n16577, n16578, n16579,
         n16580, n16581, n16582, n16583, n16584, n16585, n16586, n16587,
         n16588, n16589, n16590, n16591, n16592, n16593, n16594, n16595,
         n16596, n16597, n16598, n16599, n16600, n16601, n16602, n16603,
         n16604, n16605, n16606, n16607, n16608, n16609, n16610, n16611,
         n16612, n16613, n16614, n16615, n16616, n16617, n16618, n16619,
         n16620, n16621, n16622, n16623, n16624, n16625, n16626, n16627,
         n16628, n16629, n16630, n16631, n16632, n16633, n16634, n16635,
         n16636, n16637, n16638, n16639, n16640, n16641, n16642, n16643,
         n16644, n16645, n16646, n16647, n16648, n16649, n16650, n16651,
         n16652, n16653, n16654, n16655, n16656, n16657, n16658, n16659,
         n16660, n16661, n16662, n16663, n16664, n16665, n16666, n16667,
         n16668, n16669, n16670, n16671, n16672, n16673, n16674, n16675,
         n16676, n16677, n16678, n16679, n16680, n16681, n16682, n16683,
         n16684, n16685, n16686, n16687, n16688, n16689, n16690, n16691,
         n16692, n16693, n16694, n16695, n16696, n16697, n16698, n16699,
         n16700, n16701, n16702, n16703, n16704, n16705, n16706, n16707,
         n16708, n16709, n16710, n16711, n16712, n16713, n16714, n16715,
         n16716, n16717, n16718, n16719, n16720, n16721, n16722, n16723,
         n16724, n16725, n16726, n16727, n16728, n16729, n16730, n16731,
         n16732, n16733, n16734, n16735, n16736, n16737, n16738, n16739,
         n16740, n16741, n16742, n16743, n16744, n16745, n16746, n16747,
         n16748, n16749, n16750, n16751, n16752, n16753, n16754, n16755,
         n16756, n16757, n16758, n16759, n16760, n16761, n16762, n16763,
         n16764, n16765, n16766, n16767, n16768, n16769, n16770, n16771,
         n16772, n16773, n16774, n16775, n16776, n16777, n16778, n16779,
         n16780, n16781, n16782, n16783, n16784, n16785, n16786, n16787,
         n16788, n16789, n16790, n16791, n16792, n16793, n16794, n16795,
         n16796, n16797, n16798, n16799, n16800, n16801, n16802, n16803,
         n16804, n16805, n16806, n16807, n16808, n16809, n16810, n16811,
         n16812, n16813, n16814, n16815, n16816, n16817, n16818, n16819,
         n16820, n16821, n16822, n16823, n16824, n16825, n16826, n16827,
         n16828, n16829, n16830, n16831, n16832, n16833, n16834, n16835,
         n16836, n16837, n16838, n16839, n16840, n16841, n16842, n16843,
         n16844, n16845, n16846, n16847, n16848, n16849, n16850, n16851,
         n16852, n16853, n16854, n16855, n16856, n16857, n16858, n16859,
         n16860, n16861, n16862, n16863, n16864, n16865, n16866, n16867,
         n16868, n16869, n16870, n16871, n16872, n16873, n16874, n16875,
         n16876, n16877, n16878, n16879, n16880, n16881, n16882, n16883,
         n16884, n16885, n16886, n16887, n16888, n16889, n16890, n16891,
         n16892, n16893, n16894, n16895, n16896, n16897, n16898, n16899,
         n16900, n16901, n16902, n16903, n16904, n16905, n16906, n16907,
         n16908, n16909, n16910, n16911, n16912, n16913, n16914, n16915,
         n16916, n16917, n16918, n16919, n16920, n16921, n16922, n16923,
         n16924, n16925, n16926, n16927, n16928, n16929, n16930, n16931,
         n16932, n16933, n16934, n16935, n16936, n16937, n16938, n16939,
         n16940, n16941, n16942, n16943, n16944, n16945, n16946, n16947,
         n16948, n16949, n16950, n16951, n16952, n16953, n16954, n16955,
         n16956, n16957, n16958, n16959, n16960, n16961, n16962, n16963,
         n16964, n16965, n16966, n16967, n16968, n16969, n16970, n16971,
         n16972, n16973, n16974, n16975, n16976, n16977, n16978, n16979,
         n16980, n16981, n16982, n16983, n16984, n16985, n16986, n16987,
         n16988, n16989, n16990, n16991, n16992, n16993, n16994, n16995,
         n16996, n16997, n16998, n16999, n17000, n17001, n17002, n17003,
         n17004, n17005, n17006, n17007, n17008, n17009, n17010, n17011,
         n17012, n17013, n17014, n17015, n17016, n17017, n17018, n17019,
         n17020, n17021, n17022, n17023, n17024, n17025, n17026, n17027,
         n17028, n17029, n17030, n17031, n17032, n17033, n17034, n17035,
         n17036, n17037, n17038, n17039, n17040, n17041, n17042, n17043,
         n17044, n17045, n17046, n17047, n17048, n17049, n17050, n17051,
         n17052, n17053, n17054, n17055, n17056, n17057, n17058, n17059,
         n17060, n17061, n17062, n17063, n17064, n17065, n17066, n17067,
         n17068, n17069, n17070, n17071, n17072, n17073, n17074, n17075,
         n17076, n17077, n17078, n17079, n17080, n17081, n17082, n17083,
         n17084, n17085, n17086, n17087, n17088, n17089, n17090, n17091,
         n17092, n17093, n17094, n17095, n17096, n17097, n17098, n17099,
         n17100, n17101, n17102, n17103, n17104, n17105, n17106, n17107,
         n17108, n17109, n17110, n17111, n17112, n17113, n17114, n17115,
         n17116, n17117, n17118, n17119, n17120, n17121, n17122, n17123,
         n17124, n17125, n17126, n17127, n17128, n17129, n17130, n17131,
         n17132, n17133, n17134, n17135, n17136, n17137, n17138, n17139,
         n17140, n17141, n17142, n17143, n17144, n17145, n17146, n17147,
         n17148, n17149, n17150, n17151, n17152, n17153, n17154, n17155,
         n17156, n17157, n17158, n17159, n17160, n17161, n17162, n17163,
         n17164, n17165, n17166, n17167, n17168, n17169, n17170, n17171,
         n17172, n17173, n17174, n17175, n17176, n17177, n17178, n17179,
         n17180, n17181, n17182, n17183, n17184, n17185, n17186, n17187,
         n17188, n17189, n17190, n17191, n17192, n17193, n17194, n17195,
         n17196, n17197, n17198, n17199, n17200, n17201, n17202, n17203,
         n17204, n17205, n17206, n17207, n17208, n17209, n17210, n17211,
         n17212, n17213, n17214, n17215, n17216, n17217, n17218, n17219,
         n17220, n17221, n17222, n17223, n17224, n17225, n17226, n17227,
         n17228, n17229, n17230, n17231, n17232, n17233, n17234, n17235,
         n17236, n17237, n17238, n17239, n17240, n17241, n17242, n17243,
         n17244, n17245, n17246, n17247, n17248, n17249, n17250, n17251,
         n17252, n17253, n17254, n17255, n17256, n17257, n17258, n17259,
         n17260, n17261, n17262, n17263, n17264, n17265, n17266, n17267,
         n17268, n17269, n17270, n17271, n17272, n17273, n17274, n17275,
         n17276, n17277, n17278, n17279, n17280, n17281, n17282, n17283,
         n17284, n17285, n17286, n17287, n17288, n17289, n17290, n17291,
         n17292, n17293, n17294, n17295, n17296, n17297, n17298, n17299,
         n17300, n17301, n17302, n17303, n17304, n17305, n17306, n17307,
         n17308, n17309, n17310, n17311, n17312, n17313, n17314, n17315,
         n17316, n17317, n17318, n17319, n17320, n17321, n17322, n17323,
         n17324, n17325, n17326, n17327, n17328, n17329, n17330, n17331,
         n17332, n17333, n17334, n17335, n17336, n17337, n17338, n17339,
         n17340, n17341, n17342, n17343, n17344, n17345, n17346, n17347,
         n17348, n17349, n17350, n17351, n17352, n17353, n17354, n17355,
         n17356, n17357, n17358, n17359, n17360, n17361, n17362, n17363,
         n17364, n17365, n17366, n17367, n17368, n17369, n17370, n17371,
         n17372, n17373, n17374, n17375, n17376, n17377, n17378, n17379,
         n17380, n17381, n17382, n17383, n17384, n17385, n17386, n17387,
         n17388, n17389, n17390, n17391, n17392, n17393, n17394, n17395,
         n17396, n17397, n17398, n17399, n17400, n17401, n17402, n17403,
         n17404, n17405, n17406, n17407, n17408, n17409, n17410, n17411,
         n17412, n17413, n17414, n17415, n17416, n17417, n17418, n17419,
         n17420, n17421, n17422, n17423, n17424, n17425, n17426, n17427,
         n17428, n17429, n17430, n17431, n17432, n17433, n17434, n17435,
         n17436, n17437, n17438, n17439, n17440, n17441, n17442, n17443,
         n17444, n17445, n17446, n17447, n17448, n17449, n17450, n17451,
         n17452, n17453, n17454, n17455, n17456, n17457, n17458, n17459,
         n17460, n17461, n17462, n17463, n17464, n17465, n17466, n17467,
         n17468, n17469, n17470, n17471, n17472, n17473, n17474, n17475,
         n17476, n17477, n17478, n17479, n17480, n17481, n17482, n17483,
         n17484, n17485, n17486, n17487, n17488, n17489, n17490, n17491,
         n17492, n17493, n17494, n17495, n17496, n17497, n17498, n17499,
         n17500, n17501, n17502, n17503, n17504, n17505, n17506, n17507,
         n17508, n17509, n17510, n17511, n17512, n17513, n17514, n17515,
         n17516, n17517, n17518, n17519, n17520, n17521, n17522, n17523,
         n17524, n17525, n17526, n17527, n17528, n17529, n17530, n17531,
         n17532, n17533, n17534, n17535, n17536, n17537, n17538, n17539,
         n17540, n17541, n17542, n17543, n17544, n17545, n17546, n17547,
         n17548, n17549, n17550, n17551, n17552, n17553, n17554, n17555,
         n17556, n17557, n17558, n17559, n17560, n17561, n17562, n17563,
         n17564, n17565, n17566, n17567, n17568, n17569, n17570, n17571,
         n17572, n17573, n17574, n17575, n17576, n17577, n17578, n17579,
         n17580, n17581, n17582, n17583, n17584, n17585, n17586, n17587,
         n17588, n17589, n17590, n17591, n17592, n17593, n17594, n17595,
         n17596, n17597, n17598, n17599, n17600, n17601, n17602, n17603,
         n17604, n17605, n17606, n17607, n17608, n17609, n17610, n17611,
         n17612, n17613, n17614, n17615, n17616, n17617, n17618, n17619,
         n17620, n17621, n17622, n17623, n17624, n17625, n17626, n17627,
         n17628, n17629, n17630, n17631, n17632, n17633, n17634, n17635,
         n17636, n17637, n17638, n17639, n17640, n17641, n17642, n17643,
         n17644, n17645, n17646, n17647, n17648, n17649, n17650, n17651,
         n17652, n17653, n17654, n17655, n17656, n17657, n17658, n17659,
         n17660, n17661, n17662, n17663, n17664, n17665, n17666, n17667,
         n17668, n17669, n17670, n17671, n17672, n17673, n17674, n17675,
         n17676, n17677, n17678, n17679, n17680, n17681, n17682, n17683,
         n17684, n17685, n17686, n17687, n17688, n17689, n17690, n17691,
         n17692, n17693, n17694, n17695, n17696, n17697, n17698, n17699,
         n17700, n17701, n17702, n17703, n17704, n17705, n17706, n17707,
         n17708, n17709, n17710, n17711, n17712, n17713, n17714, n17715,
         n17716, n17717, n17718, n17719, n17720, n17721, n17722, n17723,
         n17724, n17725, n17726, n17727, n17728, n17729, n17730, n17731,
         n17732, n17733, n17734, n17735, n17736, n17737, n17738, n17739,
         n17740, n17741, n17742, n17743, n17744, n17745, n17746, n17747,
         n17748, n17749, n17750, n17751, n17752, n17753, n17754, n17755,
         n17756, n17757, n17758, n17759, n17760, n17761, n17762, n17763,
         n17764, n17765, n17766, n17767, n17768, n17769, n17770, n17771,
         n17772, n17773, n17774, n17775, n17776, n17777, n17778, n17779,
         n17780, n17781, n17782, n17783, n17784, n17785, n17786, n17787,
         n17788, n17789, n17790, n17791, n17792, n17793, n17794, n17795,
         n17796, n17797, n17798, n17799, n17800, n17801, n17802, n17803,
         n17804, n17805, n17806, n17807, n17808, n17809, n17810, n17811,
         n17812, n17813, n17814, n17815, n17816, n17817, n17818, n17819,
         n17820, n17821, n17822, n17823, n17824, n17825, n17826, n17827,
         n17828, n17829, n17830, n17831, n17832, n17833, n17834, n17835,
         n17836, n17837, n17838, n17839, n17840, n17841, n17842, n17843,
         n17844, n17845, n17846, n17847, n17848, n17849, n17850, n17851,
         n17852, n17853, n17854, n17855, n17856, n17857, n17858, n17859,
         n17860, n17861, n17862, n17863, n17864, n17865, n17866, n17867,
         n17868, n17869, n17870, n17871, n17872, n17873, n17874, n17875,
         n17876, n17877, n17878, n17879, n17880, n17881, n17882, n17883,
         n17884, n17885, n17886, n17887, n17888, n17889, n17890, n17891,
         n17892, n17893, n17894, n17895, n17896, n17897, n17898, n17899,
         n17900, n17901, n17902, n17903, n17904, n17905, n17906, n17907,
         n17908, n17909, n17910, n17911, n17912, n17913, n17914, n17915,
         n17916, n17917, n17918, n17919, n17920, n17921, n17922, n17923,
         n17924, n17925, n17926, n17927, n17928, n17929, n17930, n17931,
         n17932, n17933, n17934, n17935, n17936, n17937, n17938, n17939,
         n17940, n17941, n17942, n17943, n17944, n17945, n17946, n17947,
         n17948, n17949, n17950, n17951, n17952, n17953, n17954, n17955,
         n17956, n17957, n17958, n17959, n17960, n17961, n17962, n17963,
         n17964, n17965, n17966, n17967, n17968, n17969, n17970, n17971,
         n17972, n17973, n17974, n17975, n17976, n17977, n17978, n17979,
         n17980, n17981, n17982, n17983, n17984, n17985, n17986, n17987,
         n17988, n17989, n17990, n17991, n17992, n17993, n17994, n17995,
         n17996, n17997, n17998, n17999, n18000, n18001, n18002, n18003,
         n18004, n18005, n18006, n18007, n18008, n18009, n18010, n18011,
         n18012, n18013, n18014, n18015, n18016, n18017, n18018, n18019,
         n18020, n18021, n18022, n18023, n18024, n18025, n18026, n18027,
         n18028, n18029, n18030, n18031, n18032, n18033, n18034, n18035,
         n18036, n18037, n18038, n18039, n18040, n18041, n18042, n18043,
         n18044, n18045, n18046, n18047, n18048, n18049, n18050, n18051,
         n18052, n18053, n18054, n18055, n18056, n18057, n18058, n18059,
         n18060, n18061, n18062, n18063, n18064, n18065, n18066, n18067,
         n18068, n18069, n18070, n18071, n18072, n18073, n18074, n18075,
         n18076, n18077, n18078, n18079, n18080, n18081, n18082, n18083,
         n18084, n18085, n18086, n18087, n18088, n18089, n18090, n18091,
         n18092, n18093, n18094, n18095, n18096, n18097, n18098, n18099,
         n18100, n18101, n18102, n18103, n18104, n18105, n18106, n18107,
         n18108, n18109, n18110, n18111, n18112, n18113, n18114, n18115,
         n18116, n18117, n18118, n18119, n18120, n18121, n18122, n18123,
         n18124, n18125, n18126, n18127, n18128, n18129, n18130, n18131,
         n18132, n18133, n18134, n18135, n18136, n18137, n18138, n18139,
         n18140, n18141, n18142, n18143, n18144, n18145, n18146, n18147,
         n18148, n18149, n18150, n18151, n18152, n18153, n18154, n18155,
         n18156, n18157, n18158, n18159, n18160, n18161, n18162, n18163,
         n18164, n18165, n18166, n18167, n18168, n18169, n18170, n18171,
         n18172, n18173, n18174, n18175, n18176, n18177, n18178, n18179,
         n18180, n18181, n18182, n18183, n18184, n18185, n18186, n18187,
         n18188, n18189, n18190, n18191, n18192, n18193, n18194, n18195,
         n18196, n18197, n18198, n18199, n18200, n18201, n18202, n18203,
         n18204, n18205, n18206, n18207, n18208, n18209, n18210, n18211,
         n18212, n18213, n18214, n18215, n18216, n18217, n18218, n18219,
         n18220, n18221, n18222, n18223, n18224, n18225, n18226, n18227,
         n18228, n18229, n18230, n18231, n18232, n18233, n18234, n18235,
         n18236, n18237, n18238, n18239, n18240, n18241, n18242, n18243,
         n18244, n18245, n18246, n18247, n18248, n18249, n18250, n18251,
         n18252, n18253, n18254, n18255, n18256, n18257, n18258, n18259,
         n18260, n18261, n18262, n18263, n18264, n18265, n18266, n18267,
         n18268, n18269, n18270, n18271, n18272, n18273, n18274, n18275,
         n18276, n18277, n18278, n18279, n18280, n18281, n18282, n18283,
         n18284, n18285, n18286, n18287, n18288, n18289, n18290, n18291,
         n18292, n18293, n18294, n18295, n18296, n18297, n18298, n18299,
         n18300, n18301, n18302, n18303, n18304, n18305, n18306, n18307,
         n18308, n18309, n18310, n18311, n18312, n18313, n18314, n18315,
         n18316, n18317, n18318, n18319, n18320, n18321, n18322, n18323,
         n18324, n18325, n18326, n18327, n18328, n18329, n18330, n18331,
         n18332, n18333, n18334, n18335, n18336, n18337, n18338, n18339,
         n18340, n18341, n18342, n18343, n18344, n18345, n18346, n18347,
         n18348, n18349, n18350, n18351, n18352, n18353, n18354, n18355,
         n18356, n18357, n18358, n18359, n18360, n18361, n18362, n18363,
         n18364, n18365, n18366, n18367, n18368, n18369, n18370, n18371,
         n18372, n18373, n18374, n18375, n18376, n18377, n18378, n18379,
         n18380, n18381, n18382, n18383, n18384, n18385, n18386, n18387,
         n18388, n18389, n18390, n18391, n18392, n18393, n18394, n18395,
         n18396, n18397, n18398, n18399, n18400, n18401, n18402, n18403,
         n18404, n18405, n18406, n18407, n18408, n18409, n18410, n18411,
         n18412, n18413, n18414, n18415, n18416, n18417, n18418, n18419,
         n18420, n18421, n18422, n18423, n18424, n18425, n18426, n18427,
         n18428, n18429, n18430, n18431, n18432, n18433, n18434, n18435,
         n18436, n18437, n18438, n18439, n18440, n18441, n18442, n18443,
         n18444, n18445, n18446, n18447, n18448, n18449, n18450, n18451,
         n18452, n18453, n18454, n18455, n18456, n18457, n18458, n18459,
         n18460, n18461, n18462, n18463, n18464, n18465, n18466, n18467,
         n18468, n18469, n18470, n18471, n18472, n18473, n18474, n18475,
         n18476, n18477, n18478, n18479, n18480, n18481, n18482, n18483,
         n18484, n18485, n18486, n18487, n18488, n18489, n18490, n18491,
         n18492, n18493, n18494, n18495, n18496, n18497, n18498, n18499,
         n18500, n18501, n18502, n18503, n18504, n18505, n18506, n18507,
         n18508, n18509, n18510, n18511, n18512, n18513, n18514, n18515,
         n18516, n18517, n18518, n18519, n18520, n18521, n18522, n18523,
         n18524, n18525, n18526, n18527, n18528, n18529, n18530, n18531,
         n18532, n18533, n18534, n18535, n18536, n18537, n18538, n18539,
         n18540, n18541, n18542, n18543, n18544, n18545, n18546, n18547,
         n18548, n18549, n18550, n18551, n18552, n18553, n18554, n18555,
         n18556, n18557, n18558, n18559, n18560, n18561, n18562, n18563,
         n18564, n18565, n18566, n18567, n18568, n18569, n18570, n18571,
         n18572, n18573, n18574, n18575, n18576, n18577, n18578, n18579,
         n18580, n18581, n18582, n18583, n18584, n18585, n18586, n18587,
         n18588, n18589, n18590, n18591, n18592, n18593, n18594, n18595,
         n18596, n18597, n18598, n18599, n18600, n18601, n18602, n18603,
         n21496, n21497, n21510, n23553, n23554, n23555, n23556, n23557,
         n23558, n23559, n23560, n23561, n23562, n23563, n23564, n23565,
         n23566, n23567, n23568, n23569, n23570, n23571, n23572, n23573,
         n23574, n23575, n23576, n23577, n23578, n23579, n23580, n23581,
         n23582, n23583, n23584, n23585, n23586, n23587, n23588, n23589,
         n23590, n23591, n23592, n23593, n23594, n23595, n23596, n23597,
         n23598, n23599, n23600, n23601, n23602, n23603, n23604, n23605,
         n23606, n23607, n23608, n23609, n23610, n23611, n23612, n23613,
         n23614, n23615, n23616, n23617, n23618, n23619, n23620, n23621,
         n23622, n23623, n23624, n23625, n23626, n23627, n23628, n23629,
         n23630, n23631, n23632, n23633, n23634, n23635, n23636, n23637,
         n23638, n23639, n23640, n23641, n23642, n23643, n23644, n23645,
         n23646, n23647, n23648, n23649, n23650, n23651, n23652, n23653,
         n23654, n23655, n23656, n23657, n23658, n23659, n23660, n23661,
         n23662, n23663, n23664, n23665, n23666, n23667, n23668, n23669,
         n23670, n23671, n23672, n23673, n23674, n23675, n23676, n23677,
         n23678, n23679, n23680, n23681, n23682, n23683, n23684, n23685,
         n23686, n23687, n23688, n23689, n23690, n23691, n23692, n23693,
         n23694, n23695, n23696, n23697, n23698, n23699, n23700, n23701,
         n23702, n23703, n23704, n23705, n23706, n23707, n23708, n23709,
         n23710, n23711, n23712, n23713, n23714, n23715, n23716, n23717,
         n23718, n23719, n23720, n23721, n23722, n23723, n23724, n23725,
         n23726, n23727, n23728, n23729, n23730, n23731, n23732, n23733,
         n23734, n23735, n23736, n23737, n23738, n23739, n23740, n23741,
         n23742, n23743, n23744, n23745, n23746, n23747, n23748, n23749,
         n23750, n23751, n23752, n23753, n23754, n23755, n23756, n23757,
         n23758, n23759, n23760, n23761, n23762, n23763, n23764, n23765,
         n23766, n23767, n23768, n23769, n23770, n23771, n23772, n23773,
         n23774, n23775, n23776, n23777, n23778, n23779, n23780, n23781,
         n23782, n23783, n23784, n23785, n23786, n23787, n23788, n23789,
         n23790, n23791, n23792, n23793, n23794, n23795, n23796, n23797,
         n23798, n23799, n23800, n23801, n23802, n23803, n23804, n23805,
         n23806, n23807, n23808, n23809, n23810, n23811, n23812, n23813,
         n23814, n23815, n23816, n23817, n23818, n23819, n23820, n23821,
         n23822, n23823, n23824, n23825, n23826, n23827, n23828, n23829,
         n23830, n23831, n23832, n23833, n23834, n23835, n23836, n23837,
         n23838, n23839, n23840, n23841, n23842, n23843, n23844, n23845,
         n23846, n23847, n23848, n23849, n23850, n23851, n23852, n23853,
         n23854, n23855, n23856, n23857, n23858, n23859, n23860, n23861,
         n23862, n23863, n23864, n23865, n23866, n23867, n23868, n23869,
         n23870, n23871, n23872, n23873, n23874, n23875, n23876, n23877,
         n23878, n23879, n23880, n23881, n23882, n23883, n23884, n23885,
         n23886, n23887, n23888, n23889, n23890, n23891, n23892, n23893,
         n23894, n23895, n23896, n23897, n23898, n23899, n23900, n23901,
         n23902, n23903, n23904, n23905, n23906, n23907, n23908, n23909,
         n23910, n23911, n23912, n23913, n23914, n23915, n23916, n23917,
         n23918, n23919, n23920, n23921, n23922, n23923, n23924, n23925,
         n23926, n23927, n23928, n23929, n23930, n23931, n23932, n23933,
         n23934, n23935, n23936, n23937, n23938, n23939, n23940, n23941,
         n23942, n23943, n23944, n23945, n23946, n23947, n23948, n23949,
         n23950, n23951, n23952, n23953, n23954, n23955, n23956, n23957,
         n23958, n23959, n23960, n23961, n23962, n23963, n23964, n23965,
         n23966, n23967, n23968, n23969, n23970, n23971, n23972, n23973,
         n23974, n23975, n23976, n23977, n23978, n23979, n23980, n23981,
         n23982, n23983, n23984, n23985, n23986, n23987, n23988, n23989,
         n23990, n23991, n23992, n23993, n23994, n23995, n23996, n23997,
         n23998, n23999, n24000, n24001, n24002, n24003, n24004, n24005,
         n24006, n24007, n24008, n24009, n24010, n24011, n24012, n24013,
         n24014, n24015, n24016, n24017, n24018, n24019, n24020, n24021,
         n24022, n24023, n24024, n24025, n24026, n24027, n24028, n24029,
         n24030, n24031, n24032, n24033, n24034, n24035, n24036, n24037,
         n24038, n24039, n24040, n24041, n24042, n24043, n24044, n24045,
         n24046, n24047, n24048, n24049, n24050, n24051, n24052, n24053,
         n24054, n24055, n24056, n24057, n24058, n24059, n24060, n24061,
         n24062, n24063, n24064, n24065, n24066, n24067, n24068, n24069,
         n24070, n24071, n24072, n24073, n24074, n24075, n24076, n24077,
         n24078, n24079, n24080, n24081, n24082, n24083, n24084, n24085,
         n24086, n24087, n24088, n24089, n24090, n24091, n24092, n24093,
         n24094, n24095, n24096, n24097, n24098, n24099, n24100, n24101,
         n24102, n24103, n24104, n24105, n24106, n24107, n24108, n24109,
         n24110, n24111, n24112, n24113, n24114, n24115, n24116, n24117,
         n24118, n24119, n24120, n24121, n24122, n24123, n24124, n24125,
         n24126, n24127, n24128, n24129, n24130, n24131, n24132, n24133,
         n24134, n24135, n24136, n24137, n24138, n24139, n24140, n24141,
         n24142, n24143, n24144, n24145, n24146, n24147, n24148, n24149,
         n24150, n24151, n24152, n24153, n24154, n24155, n24156, n24157,
         n24158, n24159, n24160, n24161, n24162, n24163, n24164, n24165,
         n24166, n24167, n24168, n24169, n24170, n24171, n24172, n24173,
         n24174, n24175, n24176, n24177, n24178, n24179, n24180, n24181,
         n24182, n24183, n24184, n24185, n24186, n24187, n24188, n24189,
         n24190, n24191, n24192, n24193, n24194, n24195, n24196, n24197,
         n24198, n24199, n24200, n24201, n24202, n24203, n24204, n24205,
         n24206, n24207, n24208, n24209, n24210, n24211, n24212, n24213,
         n24214, n24215, n24216, n24217, n24218, n24219, n24220, n24221,
         n24222, n24223, n24224, n24225, n24226, n24227, n24228, n24229,
         n24230, n24231, n24232, n24233, n24234, n24235, n24236, n24237,
         n24238, n24239, n24240, n24241, n24242, n24243, n24244, n24245,
         n24246, n24247, n24248, n24249, n24250, n24251, n24252, n24253,
         n24254, n24255, n24256, n24257, n24258, n24259, n24260, n24261,
         n24262, n24263, n24264, n24265, n24266, n24267, n24268, n24269,
         n24270, n24271, n24272, n24273, n24274, n24275, n24276, n24277,
         n24278, n24279, n24280, n24281, n24282, n24283, n24284, n24285,
         n24286, n24287, n24288, n24289, n24290, n24291, n24292, n24293,
         n24294, n24295, n24296, n24297, n24298, n24299, n24300, n24301,
         n24302, n24303, n24304, n24305, n24306, n24307, n24308, n24309,
         n24310, n24311, n24312, n24313, n24314, n24315, n24316, n24317,
         n24318, n24319, n24320, n24321, n24322, n24323, n24324, n24325,
         n24326, n24327, n24328, n24329, n24330, n24331, n24332, n24333,
         n24334, n24335, n24336, n24337, n24338, n24339, n24340, n24341,
         n24342, n24343, n24344, n24345, n24346, n24347, n24348, n24349,
         n24350, n24351, n24352, n24353, n24354, n24355, n24356, n24357,
         n24358, n24359, n24360, n24361, n24362, n24363, n24364, n24365,
         n24366, n24367, n24368, n24369, n24370, n24371, n24372, n24373,
         n24374, n24375, n24376, n24377, n24378, n24379, n24380, n24381,
         n24382, n24383, n24384, n24385, n24386, n24387, n24388, n24389,
         n24390, n24391, n24392, n24393, n24394, n24395, n24396, n24397,
         n24398, n24399, n24400, n24401, n24402, n24403, n24404, n24405,
         n24406, n24407, n24408, n24409, n24410, n24411, n24412, n24413,
         n24414, n24415, n24416, n24417, n24418, n24419, n24420, n24421,
         n24422, n24423, n24424, n24425, n24426, n24427, n24428, n24429,
         n24430, n24431, n24432, n24433, n24434, n24435, n24436, n24437,
         n24438, n24439, n24440, n24441, n24442, n24443, n24444, n24445,
         n24446, n24447, n24448, n24449, n24450, n24451, n24452, n24453,
         n24454, n24455, n24456, n24457, n24458, n24459, n24460, n24461,
         n24462, n24463, n24464, n24465, n24466, n24467, n24468, n24469,
         n24470, n24471, n24472, n24473, n24474, n24475, n24476, n24477,
         n24478, n24479, n24480, n24481, n24482, n24483, n24484, n24485,
         n24486, n24487, n24488, n24489, n24490, n24491, n24492, n24493,
         n24494, n24495, n24496, n24497, n24498, n24499, n24500, n24501,
         n24502, n24503, n24504, n24505, n24506, n24507, n24508, n24509,
         n24510, n24511, n24512, n24513, n24514, n24515, n24516, n24517,
         n24518, n24519, n24520, n24521, n24522, n24523, n24524, n24525,
         n24526, n24527, n24528, n24529, n24530, n24531, n24532, n24533,
         n24534, n24535, n24536, n24537, n24538, n24539, n24540, n24541,
         n24542, n24543, n24544, n24545, n24546, n24547, n24548, n24549,
         n24550, n24551, n24552, n24553, n24554, n24555, n24556, n24557,
         n24558, n24559, n24560, n24561, n24562, n24563, n24564, n24565,
         n24566, n24567, n24568, n24569, n24570, n24571, n24572, n24573,
         n24574, n24575, n24576, n24577, n24578, n24579, n24580, n24581,
         n24582, n24583, n24584, n24585, n24586, n24587, n24588, n24589,
         n24590, n24591, n24592, n24593, n24594, n24595, n24596, n24597,
         n24598, n24599, n24600, n24601, n24602, n24603, n24604, n24605,
         n24606, n24607, n24608, n24609, n24610, n24611, n24612, n24613,
         n24614, n24615, n24616, n24617, n24618, n24619, n24620, n24621,
         n24622, n24623, n24624, n24625, n24626, n24627, n24628, n24629,
         n24630, n24631, n24632, n24633, n24634, n24635, n24636, n24637,
         n24638, n24639, n24640, n24641, n24642, n24643, n24644, n24645,
         n24646, n24647, n24648, n24649, n24650, n24651, n24652, n24653,
         n24654, n24655, n24656, n24657, n24658, n24659, n24660, n24661,
         n24662, n24663, n24664, n24665, n24666, n24667, n24668, n24669,
         n24670, n24671, n24672, n24673, n24674, n24675, n24676, n24677,
         n24678, n24679, n24680, n24681, n24682, n24683, n24684, n24685,
         n24686, n24687, n24688, n24689, n24690, n24691, n24692, n24693,
         n24694, n24695, n24696, n24697, n24698, n24699, n24700, n24701,
         n24702, n24703, n24704, n24705, n24706, n24707, n24708, n24709,
         n24710, n24711, n24712, n24713, n24714, n24715, n24716, n24717,
         n24718, n24719, n24720, n24721, n24722, n24723, n24724, n24725,
         n24726, n24727, n24728, n24729, n24730, n24731, n24732, n24733,
         n24734, n24735, n24736, n24737, n24738, n24739, n24740, n24741,
         n24742, n24743, n24744, n24745, n24746, n24747, n24748, n24749,
         n24750, n24751, n24752, n24753, n24754, n24755, n24756, n24757,
         n24758, n24759, n24760, n24761, n24762, n24763, n24764, n24765,
         n24766, n24767, n24768, n24769, n24770, n24771, n24772, n24773,
         n24774, n24775, n24776, n24777, n24778, n24779, n24780, n24781,
         n24782, n24783, n24784, n24785, n24786, n24787, n24788, n24789,
         n24790, n24791, n24792, n24793, n24794, n24795, n24796, n24797,
         n24798, n24799, n24800, n24801, n24802, n24803, n24804, n24805,
         n24806, n24807, n24808, n24809, n24810, n24811, n24812, n24813,
         n24814, n24815, n24816, n24817, n24818, n24819, n24820, n24821,
         n24822, n24823, n24824, n24825, n24826, n24827, n24828, n24829,
         n24830, n24831, n24832, n24833, n24834, n24835, n24836, n24837,
         n24838, n24839, n24840, n24841, n24842, n24843, n24844, n24845,
         n24846, n24847, n24848, n24849, n24850, n24851, n24852, n24853,
         n24854, n24855, n24856, n24857, n24858, n24859, n24860, n24861,
         n24862, n24863, n24864, n24865, n24866, n24867, n24868, n24869,
         n24870, n24871, n24872, n24873, n24874, n24875, n24876, n24877,
         n24878, n24879, n24880, n24881, n24882, n24883, n24884, n24885,
         n24886, n24887, n24888, n24889, n24890, n24891, n24892, n24893,
         n24894, n24895, n24896, n24897, n24898, n24899, n24900, n24901,
         n24902, n24903, n24904, n24905, n24906, n24907, n24908, n24909,
         n24910, n24911, n24912, n24913, n24914, n24915, n24916, n24917,
         n24918, n24919, n24920, n24921, n24922, n24923, n24924, n24925,
         n24926, n24927, n24928, n24929, n24930, n24931, n24932, n24933,
         n24934, n24935, n24936, n24937, n24938, n24939, n24940, n24941,
         n24942, n24943, n24944, n24945, n24946, n24947, n24948, n24949,
         n24950, n24951, n24952, n24953, n24954, n24955, n24956, n24957,
         n24958, n24959, n24960, n24961, n24962, n24963, n24964, n24965,
         n24966, n24967, n24968, n24969, n24970, n24971, n24972, n24973,
         n24974, n24975, n24976, n24977, n24978, n24979, n24980, n24981,
         n24982, n24983, n24984, n24985, n24986, n24987, n24988, n24989,
         n24990, n24991, n24992, n24993, n24994, n24995, n24996, n24997,
         n24998, n24999, n25000, n25001, n25002, n25003, n25004, n25005,
         n25006, n25007, n25008, n25009, n25010, n25011, n25012, n25013,
         n25014, n25015, n25016, n25017, n25018, n25019, n25020, n25021,
         n25022, n25023, n25024, n25025, n25026, n25027, n25028, n25029,
         n25030, n25031, n25032, n25033, n25034, n25035, n25036, n25037,
         n25038, n25039, n25040, n25041, n25042, n25043, n25044, n25045,
         n25046, n25047, n25048, n25049, n25050, n25051, n25052, n25053,
         n25054, n25055, n25056, n25057, n25058, n25059, n25060, n25061,
         n25062, n25063, n25064, n25065, n25066, n25067, n25068, n25069,
         n25070, n25071, n25072, n25073, n25074, n25075, n25076, n25077,
         n25078, n25079, n25080, n25081, n25082, n25083, n25084, n25085,
         n25086, n25087, n25088, n25089, n25090, n25091, n25092, n25093,
         n25094, n25095, n25096, n25097, n25098, n25099, n25100, n25101,
         n25102, n25103, n25104, n25105, n25106, n25107, n25108, n25109,
         n25110, n25111, n25112, n25113, n25114, n25115, n25116, n25117,
         n25118, n25119, n25120, n25121, n25122, n25123, n25124, n25125,
         n25126, n25127, n25128, n25129, n25130, n25131, n25132, n25133,
         n25134, n25135, n25136, n25137, n25138, n25139, n25140, n25141,
         n25142, n25143, n25144, n25145, n25146, n25147, n25148, n25149,
         n25150, n25151, n25152, n25153, n25154, n25155, n25156, n25157,
         n25158, n25159, n25160, n25161, n25162, n25163, n25164, n25165,
         n25166, n25167, n25168, n25169, n25170, n25171, n25172, n25173,
         n25174, n25175, n25176, n25177, n25178, n25179, n25180, n25181,
         n25182, n25183, n25184, n25185, n25186, n25187, n25188, n25189,
         n25190, n25191, n25192, n25193, n25194, n25195, n25196, n25197,
         n25198, n25199, n25200, n25201, n25202, n25203, n25204, n25205,
         n25206, n25207, n25208, n25209, n25210, n25211, n25212, n25213,
         n25214, n25215, n25216, n25217, n25218, n25219, n25220, n25221,
         n25222, n25223, n25224, n25225, n25226, n25227, n25228, n25229,
         n25230, n25231, n25232, n25233, n25234, n25235, n25236, n25237,
         n25238, n25239, n25240, n25241, n25242, n25243, n25244, n25245,
         n25246, n25247, n25248, n25249, n25250, n25251, n25252, n25253,
         n25254, n25255, n25256, n25257, n25258, n25259, n25260, n25261,
         n25262, n25263, n25264, n25265, n25266, n25267, n25268, n25269,
         n25270, n25271, n25272, n25273, n25274, n25275, n25276, n25277,
         n25278, n25279, n25280, n25281, n25282, n25283, n25284, n25285,
         n25286, n25287, n25288, n25289, n25290, n25291, n25292, n25293,
         n25294, n25295, n25296, n25297, n25298, n25299, n25300, n25301,
         n25302, n25303, n25304, n25305, n25306, n25307, n25308, n25309,
         n25310, n25311, n25312, n25313, n25314, n25315, n25316, n25317,
         n25318, n25319, n25320, n25321, n25322, n25323, n25324, n25325,
         n25326, n25327, n25328, n25329, n25330, n25331, n25332, n25333,
         n25334, n25335, n25336, n25337, n25338, n25339, n25340, n25341,
         n25342, n25343, n25344, n25345, n25346, n25347, n25348, n25349,
         n25350, n25351, n25352, n25353, n25354, n25355, n25356, n25357,
         n25358, n25359, n25360, n25361, n25362, n25363, n25364, n25365,
         n25366, n25367, n25368, n25369, n25370, n25371, n25372, n25373,
         n25374, n25375, n25376, n25377, n25378, n25379, n25380, n25381,
         n25382, n25383, n25384, n25385, n25386, n25387, n25388, n25389,
         n25390, n25391, n25392, n25393, n25394, n25395, n25396, n25397,
         n25398, n25399, n25400, n25401, n25402, n25403, n25404, n25405,
         n25406, n25407, n25408, n25409, n25410, n25411, n25412, n25413,
         n25414, n25415, n25416, n25417, n25418, n25419, n25420, n25421,
         n25422, n25423, n25424, n25425, n25426, n25427, n25428, n25429,
         n25430, n25431, n25432, n25433, n25434, n25435, n25436, n25437,
         n25438, n25439, n25440, n25441, n25442, n25443, n25444, n25445,
         n25446, n25447, n25448, n25449, n25450, n25451, n25452, n25453,
         n25454, n25455, n25456, n25457, n25458, n25459, n25460, n25461,
         n25462, n25463, n25464, n25465, n25466, n25467, n25468, n25469,
         n25470, n25471, n25472, n25473, n25474, n25475, n25476, n25477,
         n25478, n25479, n25480, n25481, n25482, n25483, n25484, n25485,
         n25486, n25487, n25488, n25489, n25490, n25491, n25492, n25493,
         n25494, n25495, n25496, n25497, n25498, n25499, n25500, n25501,
         n25502, n25503, n25504, n25505, n25506, n25507, n25508, n25509,
         n25510, n25511, n25512, n25513, n25514, n25515, n25516, n25517,
         n25518, n25519, n25520, n25521, n25522, n25523, n25524, n25525,
         n25526, n25527, n25528, n25529, n25530, n25531, n25532, n25533,
         n25534, n25535, n25536, n25537, n25538, n25539, n25540, n25541,
         n25542, n25543, n25544, n25545, n25546, n25547, n25548, n25549,
         n25550, n25551, n25552, n25553, n25554, n25555, n25556, n25557,
         n25558, n25559, n25560, n25561, n25562, n25563, n25564, n25565,
         n25566, n25567, n25568, n25569, n25570, n25571, n25572, n25573,
         n25574, n25575, n25576, n25577, n25578, n25579, n25580, n25581,
         n25582, n25583, n25584, n25585, n25586, n25587, n25588, n25589,
         n25590, n25591, n25592, n25593, n25594, n25595, n25596, n25597,
         n25598, n25599, n25600, n25601, n25602, n25603, n25604, n25605,
         n25606, n25607, n25608, n25609, n25610, n25611, n25612, n25613,
         n25614, n25615, n25616, n25617, n25618, n25619, n25620, n25621,
         n25622, n25623, n25624, n25625, n25626, n25627, n25628, n25629,
         n25630, n25631, n25632, n25633, n25634, n25635, n25636, n25637,
         n25638, n25639, n25640, n25641, n25642, n25643, n25644, n25645,
         n25646, n25647, n25648, n25649, n25650, n25651, n25652, n25653,
         n25654, n25655, n25656, n25657, n25658, n25659, n25660, n25661,
         n25662, n25663, n25664, n25665, n25666, n25667, n25668, n25669,
         n25670, n25671, n25672, n25673, n25674, n25675, n25676, n25677,
         n25678, n25679, n25680, n25681, n25682, n25683, n25684, n25685,
         n25686, n25687, n25688, n25689, n25690, n25691, n25692, n25693,
         n25694, n25695, n25696, n25697, n25698, n25699, n25700, n25701,
         n25702, n25703, n25704, n25705, n25706, n25707, n25708, n25709,
         n25710, n25711, n25712, n25713, n25714, n25715, n25716, n25717,
         n25718, n25719, n25720, n25721, n25722, n25723, n25724, n25725,
         n25726, n25727, n25728, n25729, n25730, n25731, n25732, n25733,
         n25734, n25735, n25736, n25737, n25738, n25739, n25740, n25741,
         n25742, n25743, n25744, n25745, n25746, n25747, n25748, n25749,
         n25750, n25751, n25752, n25753, n25754, n25755, n25756, n25757,
         n25758, n25759, n25760, n25761, n25762, n25763, n25764, n25765,
         n25766, n25767, n25768, n25769, n25770, n25771, n25772, n25773,
         n25774, n25775, n25776, n25777, n25778, n25779, n25780, n25781,
         n25782, n25783, n25784, n25785, n25786, n25787, n25788, n25789,
         n25790, n25791, n25792, n25793, n25794, n25795, n25796, n25797,
         n25798, n25799, n25800, n25801, n25802, n25803, n25804, n25805,
         n25806, n25807, n25808, n25809, n25810, n25811, n25812, n25813,
         n25814, n25815, n25816, n25817, n25818, n25819, n25820, n25821,
         n25822, n25823, n25824, n25825, n25826, n25827, n25828, n25829,
         n25830, n25831, n25832, n25833, n25834, n25835, n25836, n25837,
         n25838, n25839, n25840, n25841, n25842, n25843, n25844, n25845,
         n25846, n25847, n25848, n25849, n25850, n25851, n25852, n25853,
         n25854, n25855, n25856, n25857, n25858, n25859, n25860, n25861,
         n25862, n25863, n25864, n25865, n25866, n25867, n25868, n25869,
         n25870, n25871, n25872, n25873, n25874, n25875, n25876, n25877,
         n25878, n25879, n25880, n25881, n25882, n25883, n25884, n25885,
         n25886, n25887, n25888, n25889, n25890, n25891, n25892, n25893,
         n25894, n25895, n25896, n25897, n25898, n25899, n25900, n25901,
         n25902, n25903, n25904, n25905, n25906, n25907, n25908, n25909,
         n25910, n25911, n25912, n25913, n25914, n25915, n25916, n25917,
         n25918, n25919, n25920, n25921, n25922, n25923, n25924, n25925,
         n25926, n25927, n25928, n25929, n25930, n25931, n25932, n25933,
         n25934, n25935, n25936, n25937, n25938, n25939, n25940, n25941,
         n25942, n25943, n25944, n25945, n25946, n25947, n25948, n25949,
         n25950, n25951, n25952, n25953, n25954, n25955, n25956, n25957,
         n25958, n25959, n25960, n25961, n25962, n25963, n25964, n25965,
         n25966, n25967, n25968, n25969, n25970, n25971, n25972, n25973,
         n25974, n25975, n25976, n25977, n25978, n25979, n25980, n25981,
         n25982, n25983, n25984, n25985, n25986, n25987, n25988, n25989,
         n25990, n25991, n25992, n25993, n25994, n25995, n25996, n25997,
         n25998, n25999, n26000, n26001, n26002, n26003, n26004, n26005,
         n26006, n26007, n26008, n26009, n26010, n26011, n26012, n26013,
         n26014, n26015, n26016, n26017, n26018, n26019, n26020, n26021,
         n26022, n26023, n26024, n26025, n26026, n26027, n26028, n26029,
         n26030, n26031, n26032, n26033, n26034, n26035, n26036, n26037,
         n26038, n26039, n26040, n26041, n26042, n26043, n26044, n26045,
         n26046, n26047, n26048, n26049, n26050, n26051, n26052, n26053,
         n26054, n26055, n26056, n26057, n26058, n26059, n26060, n26061,
         n26062, n26063, n26064, n26065, n26066, n26067, n26068, n26069,
         n26070, n26071, n26072, n26073, n26074, n26075, n26076, n26077,
         n26078, n26079, n26080, n26081, n26082, n26083, n26084, n26085,
         n26086, n26087, n26088, n26089, n26090, n26091, n26092, n26093,
         n26094, n26095, n26096, n26097, n26098, n26099, n26100, n26101,
         n26102, n26103, n26104, n26105, n26106, n26107, n26108, n26109,
         n26110, n26111, n26112, n26113, n26114, n26115, n26116, n26117,
         n26118, n26119, n26120, n26121, n26122, n26123, n26124, n26125,
         n26126, n26127, n26128, n26129, n26130, n26131, n26132, n26133,
         n26134, n26135, n26136, n26137, n26138, n26139, n26140, n26141,
         n26142, n26143, n26144, n26145, n26146, n26147, n26148, n26149,
         n26150, n26151, n26152, n26153, n26154, n26155, n26156, n26157,
         n26158, n26159, n26160, n26161, n26162, n26163, n26164, n26165,
         n26166, n26167, n26168, n26169, n26170, n26171, n26172, n26173,
         n26174, n26175, n26176, n26177, n26178, n26179, n26180, n26181,
         n26182, n26183, n26184, n26185, n26186, n26187, n26188, n26189,
         n26190, n26191, n26192, n26193, n26194, n26195, n26196, n26197,
         n26198, n26199, n26200, n26201, n26202, n26203, n26204, n26205,
         n26206, n26207, n26208, n26209, n26210, n26211, n26212, n26213,
         n26214, n26215, n26216, n26217, n26218, n26219, n26220, n26221,
         n26222, n26223, n26224, n26225, n26226, n26227, n26228, n26229,
         n26230, n26231, n26232, n26233, n26234, n26235, n26236, n26237,
         n26238, n26239, n26240, n26241, n26242, n26243, n26244, n26245,
         n26246, n26247, n26248, n26249, n26250, n26251, n26252, n26253,
         n26254, n26255, n26256, n26257, n26258, n26259, n26260, n26261,
         n26262, n26263, n26264, n26265, n26266, n26267, n26268, n26269,
         n26270, n26271, n26272, n26273, n26274, n26275, n26276, n26277,
         n26278, n26279, n26280, n26281, n26282, n26283, n26284, n26285,
         n26286, n26287, n26288, n26289, n26290, n26291, n26292, n26293,
         n26294, n26295, n26296, n26297, n26298, n26299, n26300, n26301,
         n26302, n26303, n26304, n26305, n26306, n26307, n26308, n26309,
         n26310, n26311, n26312, n26313, n26314, n26315, n26316, n26317,
         n26318, n26319, n26320, n26321, n26322, n26323, n26324, n26325,
         n26326, n26327, n26328, n26329, n26330, n26331, n26332, n26333,
         n26334, n26335, n26336, n26337, n26338, n26339, n26340, n26341,
         n26342, n26343, n26344, n26345, n26346, n26347, n26348, n26349,
         n26350, n26351, n26352, n26353, n26354, n26355, n26356, n26357,
         n26358, n26359, n26360, n26361, n26362, n26363, n26364, n26365,
         n26366, n26367, n26368, n26369, n26370, n26371, n26372, n26373,
         n26374, n26375, n26376, n26377, n26378, n26379, n26380, n26381,
         n26382, n26383, n26384, n26385, n26386, n26387, n26388, n26389,
         n26390, n26391, n26392, n26393, n26394, n26395, n26396, n26397,
         n26398, n26399, n26400, n26401, n26402, n26403, n26404, n26405,
         n26406, n26407, n26408, n26409, n26410, n26411, n26412, n26413,
         n26414, n26415, n26416, n26417, n26418, n26419, n26420, n26421,
         n26422, n26423, n26424, n26425, n26426, n26427, n26428, n26429,
         n26430, n26431, n26432, n26433, n26434, n26435, n26436, n26437,
         n26438, n26439, n26440, n26441, n26442, n26443, n26444, n26445,
         n26446, n26447, n26448, n26449, n26450, n26451, n26452, n26453,
         n26454, n26455, n26456, n26457, n26458, n26459, n26460, n26461,
         n26462, n26463, n26464, n26465, n26466, n26467, n26468, n26469,
         n26470, n26471, n26472, n26473, n26474, n26475, n26476, n26477,
         n26478, n26479, n26480, n26481, n26482, n26483, n26484, n26485,
         n26486, n26487, n26488, n26489, n26490, n26491, n26492, n26493,
         n26494, n26495, n26496, n26497, n26498, n26499, n26500, n26501,
         n26502, n26503, n26504, n26505, n26506, n26507, n26508, n26509,
         n26510, n26511, n26512, n26513, n26514, n26515, n26516, n26517,
         n26518, n26519, n26520, n26521, n26522, n26523, n26524, n26525,
         n26526, n26527, n26528, n26529, n26530, n26531, n26532, n26533,
         n26534, n26535, n26536, n26537, n26538, n26539, n26540, n26541,
         n26542, n26543, n26544, n26545, n26546, n26547, n26548, n26549,
         n26550, n26551, n26552, n26553, n26554, n26555, n26556, n26557,
         n26558, n26559, n26560, n26561, n26562, n26563, n26564, n26565,
         n26566, n26567, n26568, n26569, n26570, n26571, n26572, n26573,
         n26574, n26575, n26576, n26577, n26578, n26579, n26580, n26581,
         n26582, n26583, n26584, n26585, n26586, n26587, n26588, n26589,
         n26590, n26591, n26592, n26593, n26594, n26595, n26596, n26597,
         n26598, n26599, n26600, n26601, n26602, n26603, n26604, n26605,
         n26606, n26607, n26608, n26609, n26610, n26611, n26612, n26613,
         n26614, n26615, n26616, n26617, n26618, n26619, n26620, n26621,
         n26622, n26623, n26624, n26625, n26626, n26627, n26628, n26629,
         n26630, n26631, n26632, n26633, n26634, n26635, n26636, n26637,
         n26638, n26639, n26640, n26641, n26642, n26643, n26644, n26645,
         n26646, n26647, n26648, n26649, n26650, n26651, n26652, n26653,
         n26654, n26655, n26656, n26657, n26658, n26659, n26660, n26661,
         n26662, n26663, n26664, n26665, n26666, n26667, n26668, n26669,
         n26670, n26671, n26672, n26673, n26674, n26675, n26676, n26677,
         n26678, n26679, n26680, n26681, n26682, n26683, n26684, n26685,
         n26686, n26687, n26688, n26689, n26690, n26691, n26692, n26693,
         n26694, n26695, n26696, n26697, n26698, n26699, n26700, n26701,
         n26702, n26703, n26704, n26705, n26706, n26707, n26708, n26709,
         n26710, n26711, n26712, n26713, n26714, n26715, n26716, n26717,
         n26718, n26719, n26720, n26721, n26722, n26723, n26724, n26725,
         n26726, n26727, n26728, n26729, n26730, n26731, n26732, n26733,
         n26734, n26735, n26736, n26737, n26738, n26739, n26740, n26741,
         n26742, n26743, n26744, n26745, n26746, n26747, n26748, n26749,
         n26750, n26751, n26752, n26753, n26754, n26755, n26756, n26757,
         n26758, n26759, n26760, n26761, n26762, n26763, n26764, n26765,
         n26766, n26767, n26768, n26769, n26770, n26771, n26772, n26773,
         n26774, n26775, n26776, n26777, n26778, n26779, n26780, n26781,
         n26782, n26783, n26784, n26785, n26786, n26787, n26788, n26789,
         n26790, n26791, n26792, n26793, n26794, n26795, n26796, n26797,
         n26798, n26799, n26800, n26801, n26802, n26803, n26804, n26805,
         n26806, n26807, n26808, n26809, n26810, n26811, n26812, n26813,
         n26814, n26815, n26816, n26817, n26818, n26819, n26820, n26821,
         n26822, n26823, n26824, n26825, n26826, n26827, n26828, n26829,
         n26830, n26831, n26832, n26833, n26834, n26835, n26836, n26837,
         n26838, n26839, n26840, n26841, n26842, n26843, n26844, n26845,
         n26846, n26847, n26848, n26849, n26850, n26851, n26852, n26853,
         n26854, n26855, n26856, n26857, n26858, n26859, n26860, n26861,
         n26862, n26863, n26864, n26865, n26866, n26867, n26868, n26869,
         n26870, n26871, n26872, n26873, n26874, n26875, n26876, n26877,
         n26878, n26879, n26880, n26881, n26882, n26883, n26884, n26885,
         n26886, n26887, n26888, n26889, n26890, n26891, n26892, n26893,
         n26894, n26895, n26896, n26897, n26898, n26899, n26900, n26901,
         n26902, n26903, n26904, n26905, n26906, n26907, n26908, n26909,
         n26910, n26911, n26912, n26913, n26914, n26915, n26916, n26917,
         n26918, n26919, n26920, n26921, n26922, n26923, n26924, n26925,
         n26926, n26927, n26928, n26929, n26930, n26931, n26932, n26933,
         n26934, n26935, n26936, n26937, n26938, n26939, n26940, n26941,
         n26942, n26943, n26944, n26945, n26946, n26947, n26948, n26949,
         n26950, n26951, n26952, n26953, n26954, n26955, n26956, n26957,
         n26958, n26959, n26960, n26961, n26962, n26963, n26964, n26965,
         n26966, n26967, n26968, n26969, n26970, n26971, n26972, n26973,
         n26974, n26975, n26976, n26977, n26978, n26979, n26980, n26981,
         n26982, n26983, n26984, n26985, n26986, n26987, n26988, n26989,
         n26990, n26991, n26992, n26993, n26994, n26995, n26996, n26997,
         n26998, n26999, n27000, n27001, n27002, n27003, n27004, n27005,
         n27006, n27007, n27008, n27009, n27010, n27011, n27012, n27013,
         n27014, n27015, n27016, n27017, n27018, n27019, n27020, n27021,
         n27022, n27023, n27024, n27025, n27026, n27027, n27028, n27029,
         n27030, n27031, n27032, n27033, n27034, n27035, n27036, n27037,
         n27038, n27039, n27040, n27041, n27042, n27043, n27044, n27045,
         n27046, n27047, n27048, n27049, n27050, n27051, n27052, n27053,
         n27054, n27055, n27056, n27057, n27058, n27059, n27060, n27061,
         n27062, n27063, n27064, n27065, n27066, n27067, n27068, n27069,
         n27070, n27071, n27072, n27073, n27074, n27075, n27076, n27077,
         n27078, n27079, n27080, n27081, n27082, n27083, n27084, n27085,
         n27086, n27087, n27088, n27089, n27090, n27091, n27092, n27093,
         n27094, n27095, n27096, n27097, n27098, n27099, n27100, n27101,
         n27102, n27103, n27104, n27105, n27106, n27107, n27108, n27109,
         n27110, n27111, n27112, n27113, n27114, n27115, n27116, n27117,
         n27118, n27119, n27120, n27121, n27122, n27123, n27124, n27125,
         n27126, n27127, n27128, n27129, n27130, n27131, n27132, n27133,
         n27134, n27135, n27136, n27137, n27138, n27139, n27140, n27141,
         n27142, n27143, n27144, n27145, n27146, n27147, n27148, n27149,
         n27150, n27151, n27152, n27153, n27154, n27155, n27156, n27157,
         n27158, n27159, n27160, n27161, n27162, n27163, n27164, n27165,
         n27166, n27167, n27168, n27169, n27170, n27171, n27172, n27173,
         n27174, n27175, n27176, n27177, n27178, n27179, n27180, n27181,
         n27182, n27183, n27184, n27185, n27186, n27187, n27188, n27189,
         n27190, n27191, n27192, n27193, n27194, n27195, n27196, n27197,
         n27198, n27199, n27200, n27201, n27202, n27203, n27204, n27205,
         n27206, n27207, n27208, n27209, n27210, n27211, n27212, n27213,
         n27214, n27215, n27216, n27217, n27218, n27219, n27220, n27221,
         n27222, n27223, n27224, n27225, n27226, n27227, n27228, n27229,
         n27230, n27231, n27232, n27233, n27234, n27235, n27236, n27237,
         n27238, n27239, n27240, n27241, n27242, n27243, n27244, n27245,
         n27246, n27247, n27248, n27249, n27250, n27251, n27252, n27253,
         n27254, n27255, n27256, n27257, n27258, n27259, n27260, n27261,
         n27262, n27263, n27264, n27265, n27266, n27267, n27268, n27269,
         n27270, n27271, n27272, n27273, n27274, n27275, n27276, n27277,
         n27278, n27279, n27280, n27281, n27282, n27283, n27284, n27285,
         n27286, n27287, n27288, n27289, n27290, n27291, n27292, n27293,
         n27294, n27295, n27296, n27297, n27298, n27299, n27300, n27301,
         n27302, n27303, n27304, n27305, n27306, n27307, n27308, n27309,
         n27310, n27311, n27312, n27313, n27314, n27315, n27316, n27317,
         n27318, n27319, n27320, n27321, n27322, n27323, n27324, n27325,
         n27326, n27327, n27328, n27329, n27330, n27331, n27332, n27333,
         n27334, n27335, n27336, n27337, n27338, n27339, n27340, n27341,
         n27342, n27343, n27344, n27345, n27346, n27347, n27348, n27349,
         n27350, n27351, n27352, n27353, n27354, n27355, n27356, n27357,
         n27358, n27359, n27360, n27361, n27362, n27363, n27364, n27365,
         n27366, n27367, n27368, n27369, n27370, n27371, n27372, n27373,
         n27374, n27375, n27376, n27377, n27378, n27379, n27380, n27381,
         n27382, n27383, n27384, n27385, n27386, n27387, n27388, n27389,
         n27390, n27391, n27392, n27393, n27394, n27395, n27396, n27397,
         n27398, n27399, n27400, n27401, n27402, n27403, n27404, n27405,
         n27406, n27407, n27408, n27409, n27410, n27411, n27412, n27413,
         n27414, n27415, n27416, n27417, n27418, n27419, n27420, n27421,
         n27422, n27423, n27424, n27425, n27426, n27427, n27428, n27429,
         n27430, n27431, n27432, n27433, n27434, n27435, n27436, n27437,
         n27438, n27439, n27440, n27441, n27442, n27443, n27444, n27445,
         n27446, n27447, n27448, n27449, n27450, n27451, n27452, n27453,
         n27454, n27455, n27456, n27457, n27458, n27459, n27460, n27461,
         n27462, n27463, n27464, n27465, n27466, n27467, n27468, n27469,
         n27470, n27471, n27472, n27473, n27474, n27475, n27476, n27477,
         n27478, n27479, n27480, n27481, n27482, n27483, n27484, n27485,
         n27486, n27487, n27488, n27489, n27490, n27491, n27492, n27493,
         n27494, n27495, n27496, n27497, n27498, n27499, n27500, n27501,
         n27502, n27503, n27504, n27505, n27506, n27507, n27508, n27509,
         n27510, n27511, n27512, n27513, n27514, n27515, n27516, n27517,
         n27518, n27519, n27520, n27521, n27522, n27523, n27524, n27525,
         n27526, n27527, n27528, n27529, n27530, n27531, n27532, n27533,
         n27534, n27535, n27536, n27537, n27538, n27539, n27540, n27541,
         n27542, n27543, n27544, n27545, n27546, n27547, n27548, n27549,
         n27550, n27551, n27552, n27553, n27554, n27555, n27556, n27557,
         n27558, n27559, n27560, n27561, n27562, n27563, n27564, n27565,
         n27566, n27567, n27568, n27569, n27570, n27571, n27572, n27573,
         n27574, n27575, n27576, n27577, n27578, n27579, n27580, n27581,
         n27582, n27583, n27584, n27585, n27586, n27587, n27588, n27589,
         n27590, n27591, n27592, n27593, n27594, n27595, n27596, n27597,
         n27598, n27599, n27600, n27601, n27602, n27603, n27604, n27605,
         n27606, n27607, n27608, n27609, n27610, n27611, n27612, n27613,
         n27614, n27615, n27616, n27617, n27618, n27619, n27620, n27621,
         n27622, n27623, n27624, n27625, n27626, n27627, n27628, n27629,
         n27630, n27631, n27632, n27633, n27634, n27635, n27636, n27637,
         n27638, n27639, n27640, n27641, n27642, n27643, n27644, n27645,
         n27646, n27647, n27648, n27649, n27650, n27651, n27652, n27653,
         n27654, n27655, n27656, n27657, n27658, n27659, n27660, n27661,
         n27662, n27663, n27664, n27665, n27666, n27667, n27668, n27669,
         n27670, n27671, n27672, n27673, n27674, n27675, n27676, n27677,
         n27678, n27679, n27680, n27681, n27682, n27683, n27684, n27685,
         n27686, n27687, n27688, n27689, n27690, n27691, n27692, n27693,
         n27694, n27695, n27696, n27697, n27698, n27699, n27700, n27701,
         n27702, n27703, n27704, n27705, n27706, n27707, n27708, n27709,
         n27710, n27711, n27712, n27713, n27714, n27715, n27716, n27717,
         n27718, n27719, n27720, n27721, n27722, n27723, n27724, n27725,
         n27726, n27727, n27728, n27729, n27730, n27731, n27732, n27733,
         n27734, n27735, n27736, n27737, n27738, n27739, n27740, n27741,
         n27742, n27743, n27744, n27745, n27746, n27747, n27748, n27749,
         n27750, n27751, n27752, n27753, n27754, n27755, n27756, n27757,
         n27758, n27759, n27760, n27761, n27762, n27763, n27764, n27765,
         n27766, n27767, n27768, n27769, n27770, n27771, n27772, n27773,
         n27774, n27775, n27776, n27777, n27778, n27779, n27780, n27781,
         n27782, n27783, n27784, n27785, n27786, n27787, n27788, n27789,
         n27790, n27791, n27792, n27793, n27794, n27795, n27796, n27797,
         n27798, n27799, n27800, n27801, n27802, n27803, n27804, n27805,
         n27806, n27807, n27808, n27809, n27810, n27811, n27812, n27813,
         n27814, n27815, n27816, n27817, n27818, n27819, n27820, n27821,
         n27822, n27823, n27824, n27825, n27826, n27827, n27828, n27829,
         n27830, n27831, n27832, n27833, n27834, n27835, n27836, n27837,
         n27838, n27839, n27840, n27841, n27842, n27843, n27844, n27845,
         n27846, n27847, n27848, n27849, n27850, n27851, n27852, n27853,
         n27854, n27855, n27856, n27857, n27858, n27859, n27860, n27861,
         n27862, n27863, n27864, n27865, n27866, n27867, n27868, n27869,
         n27870, n27871, n27872, n27873, n27874, n27875, n27876, n27877,
         n27878, n27879, n27880, n27881, n27882, n27883, n27884, n27885,
         n27886, n27887, n27888, n27889, n27890, n27891, n27892, n27893,
         n27894, n27895, n27896, n27897, n27898, n27899, n27900, n27901,
         n27902, n27903, n27904, n27905, n27906, n27907, n27908, n27909,
         n27910, n27911, n27912, n27913, n27914, n27915, n27916, n27917,
         n27918, n27919, n27920, n27921, n27922, n27923, n27924, n27925,
         n27926, n27927, n27928, n27929, n27930, n27931, n27932, n27933,
         n27934, n27935, n27936, n27937, n27938, n27939, n27940, n27941,
         n27942, n27943, n27944, n27945, n27946, n27947, n27948, n27949,
         n27950, n27951, n27952, n27953, n27954, n27955, n27956, n27957,
         n27958, n27959, n27960, n27961, n27962, n27963, n27964, n27965,
         n27966, n27967, n27968, n27969, n27970, n27971, n27972, n27973,
         n27974, n27975, n27976, n27977, n27978, n27979, n27980, n27981,
         n27982, n27983, n27984, n27985, n27986, n27987, n27988, n27989,
         n27990, n27991, n27992, n27993, n27994, n27995, n27996, n27997,
         n27998, n27999, n28000, n28001, n28002, n28003, n28004, n28005,
         n28006, n28007, n28008, n28009, n28010, n28011, n28012, n28013,
         n28014, n28015, n28016, n28017, n28018, n28019, n28020, n28021,
         n28022, n28023, n28024, n28025, n28026, n28027, n28028, n28029,
         n28030, n28031, n28032, n28033, n28034, n28035, n28036, n28037,
         n28038, n28039, n28040, n28041, n28042, n28043, n28044, n28045,
         n28046, n28047, n28048, n28049, n28050, n28051, n28052, n28053,
         n28054, n28055, n28056, n28057, n28058, n28059, n28060, n28061,
         n28062, n28063, n28064, n28065, n28066, n28067, n28068, n28069,
         n28070, n28071, n28072, n28073, n28074, n28075, n28076, n28077,
         n28078, n28079, n28080, n28081, n28082, n28083, n28084, n28085,
         n28086, n28087, n28088, n28089, n28090, n28091, n28092, n28093,
         n28094, n28095, n28096, n28097, n28098, n28099, n28100, n28101,
         n28102, n28103, n28104, n28105, n28106, n28107, n28108, n28109,
         n28110, n28111, n28112, n28113, n28114, n28115, n28116, n28117,
         n28118, n28119, n28120, n28121, n28122, n28123, n28124, n28125,
         n28126, n28127, n28128, n28129, n28130, n28131, n28132, n28133,
         n28134, n28135, n28136, n28137, n28138, n28139, n28140, n28141,
         n28142, n28143, n28144, n28145, n28146, n28147, n28148, n28149,
         n28150, n28151, n28152, n28153, n28154, n28155, n28156, n28157,
         n28158, n28159, n28160, n28161, n28162, n28163, n28164, n28165,
         n28166, n28167, n28168, n28169, n28170, n28171, n28172, n28173,
         n28174, n28175, n28176, n28177, n28178, n28179, n28180, n28181,
         n28182, n28183, n28184, n28185, n28186, n28187, n28188, n28189,
         n28190, n28191, n28192, n28193, n28194, n28195, n28196, n28197,
         n28198, n28199, n28200, n28201, n28202, n28203, n28204, n28205,
         n28206, n28207, n28208, n28209, n28210, n28211, n28212, n28213,
         n28214, n28215, n28216, n28217, n28218, n28219, n28220, n28221,
         n28222, n28223, n28224, n28225, n28226, n28227, n28228, n28229,
         n28230, n28231, n28232, n28233, n28234, n28235, n28236, n28237,
         n28238, n28239, n28240, n28241, n28242, n28243, n28244, n28245,
         n28246, n28247, n28248, n28249, n28250, n28251, n28252, n28253,
         n28254, n28255, n28256, n28257, n28258, n28259, n28260, n28261,
         n28262, n28263, n28264, n28265, n28266, n28267, n28268, n28269,
         n28270, n28271, n28272, n28273, n28274, n28275, n28276, n28277,
         n28278, n28279, n28280, n28281, n28282, n28283, n28284, n28285,
         n28286, n28287, n28288, n28289, n28290, n28291, n28292, n28293,
         n28294, n28295, n28296, n28297, n28298, n28299, n28300, n28301,
         n28302, n28303, n28304, n28305, n28306, n28307, n28308, n28309,
         n28310, n28311, n28312, n28313, n28314, n28315, n28316, n28317,
         n28318, n28319, n28320, n28321, n28322, n28323, n28324, n28325,
         n28326, n28327, n28328, n28329, n28330, n28331, n28332, n28333,
         n28334, n28335, n28336, n28337, n28338, n28339, n28340, n28341,
         n28342, n28343, n28344, n28345, n28346, n28347, n28348, n28349,
         n28350, n28351, n28352, n28353, n28354, n28355, n28356, n28357,
         n28358, n28359, n28360, n28361, n28362, n28363, n28364, n28365,
         n28366, n28367, n28368, n28369, n28370, n28371, n28372, n28373,
         n28374, n28375, n28376, n28377, n28378, n28379, n28380, n28381,
         n28382, n28383, n28384, n28385, n28386, n28387, n28388, n28389,
         n28390, n28391, n28392, n28393, n28394, n28395, n28396, n28397,
         n28398, n28399, n28400, n28401, n28402, n28403, n28404, n28405,
         n28406, n28407, n28408, n28409, n28410, n28411, n28412, n28413,
         n28414, n28415, n28416, n28417, n28418, n28419, n28420, n28421,
         n28422, n28423, n28424, n28425, n28426, n28427, n28428, n28429,
         n28430, n28431, n28432, n28433, n28434, n28435, n28436, n28437,
         n28438, n28439, n28440, n28441, n28442, n28443, n28444, n28445,
         n28446, n28447, n28448, n28449, n28450, n28451, n28452, n28453,
         n28454, n28455, n28456, n28457, n28458, n28459, n28460, n28461,
         n28462, n28463, n28464, n28465, n28466, n28467, n28468, n28469,
         n28470, n28471, n28472, n28473, n28474, n28475, n28476, n28477,
         n28478, n28479, n28480, n28481, n28482, n28483, n28484, n28485,
         n28486, n28487, n28488, n28489, n28490, n28491, n28492, n28493,
         n28494, n28495, n28496, n28497, n28498, n28499, n28500, n28501,
         n28502, n28503, n28504, n28505, n28506, n28507, n28508, n28509,
         n28510, n28511, n28512, n28513, n28514, n28515, n28516, n28517,
         n28518, n28519, n28520, n28521, n28522, n28523, n28524, n28525,
         n28526, n28527, n28528, n28529, n28530, n28531, n28532, n28533,
         n28534, n28535, n28536, n28537, n28538, n28539, n28540, n28541,
         n28542, n28543, n28544, n28545, n28546, n28547, n28548, n28549,
         n28550, n28551, n28552, n28553, n28554, n28555, n28556, n28557,
         n28558, n28559, n28560, n28561, n28562, n28563, n28564, n28565,
         n28566, n28567, n28568, n28569, n28570, n28571, n28572, n28573,
         n28574, n28575, n28576, n28577, n28578, n28579, n28580, n28581,
         n28582, n28583, n28584, n28585, n28586, n28587, n28588, n28589,
         n28590, n28591, n28592, n28593, n28594, n28595, n28596, n28597,
         n28598, n28599, n28600, n28601, n28602, n28603, n28604, n28605,
         n28606, n28607, n28608, n28609, n28610, n28611, n28612, n28613,
         n28614, n28615, n28616, n28617, n28618, n28619, n28620, n28621,
         n28622, n28623, n28624, n28625, n28626, n28627, n28628, n28629,
         n28630, n28631, n28632, n28633, n28634, n28635, n28636, n28637,
         n28638, n28639, n28640, n28641, n28642, n28643, n28644, n28645,
         n28646, n28647, n28648, n28649, n28650, n28651, n28652, n28653,
         n28654, n28655, n28656, n28657, n28658, n28659, n28660, n28661,
         n28662, n28663, n28664, n28665, n28666, n28667, n28668, n28669,
         n28670, n28671, n28672, n28673, n28674, n28675, n28676, n28677,
         n28678, n28679, n28680, n28681, n28682, n28683, n28684, n28685,
         n28686, n28687, n28688, n28689, n28690, n28691, n28692, n28693,
         n28694, n28695, n28696, n28697, n28698, n28699, n28700, n28701,
         n28702, n28703, n28704, n28705, n28706, n28707, n28708, n28709,
         n28710, n28711, n28712, n28713, n28714, n28715, n28716, n28717,
         n28718, n28719, n28720, n28721, n28722, n28723, n28724, n28725,
         n28726, n28727, n28728, n28729, n28730, n28731, n28732, n28733,
         n28734, n28735, n28736, n28737, n28738, n28739, n28740, n28741,
         n28742, n28743, n28744, n28745, n28746, n28747, n28748, n28749,
         n28750, n28751, n28752, n28753, n28754, n28755, n28756, n28757,
         n28758, n28759, n28760, n28761, n28762, n28763, n28764, n28765,
         n28766, n28767, n28768, n28769, n28770, n28771, n28772, n28773,
         n28774, n28775, n28776, n28777, n28778, n28779, n28780, n28781,
         n28782, n28783, n28784, n28785, n28786, n28787, n28788, n28789,
         n28790, n28791, n28792, n28793, n28794, n28795, n28796, n28797,
         n28798, n28799, n28800, n28801, n28802, n28803, n28804, n28805,
         n28806, n28807, n28808, n28809, n28810, n28811, n28812, n28813,
         n28814, n28815, n28816, n28817, n28818, n28819, n28820, n28821,
         n28822, n28823, n28824, n28825, n28826, n28827, n28828, n28829,
         n28830, n28831, n28832, n28833, n28834, n28835, n28836, n28837,
         n28838, n28839, n28840, n28841, n28842, n28843, n28844, n28845,
         n28846, n28847, n28848, n28849, n28850, n28851, n28852, n28853,
         n28854, n28855, n28856, n28857, n28858, n28859, n28860, n28861,
         n28862, n28863, n28864, n28865, n28866, n28867, n28868, n28869,
         n28870, n28871, n28872, n28873, n28874, n28875, n28876, n28877,
         n28878, n28879, n28880, n28881, n28882, n28883, n28884, n28885,
         n28886, n28887, n28888, n28889, n28890, n28891, n28892, n28893,
         n28894, n28895, n28896, n28897, n28898, n28899, n28900, n28901,
         n28902, n28903, n28904, n28905, n28906, n28907, n28908, n28909,
         n28910, n28911, n28912, n28913, n28914, n28915, n28916, n28917,
         n28918, n28919, n28920, n28921, n28922, n28923, n28924, n28925,
         n28926, n28927, n28928, n28929, n28930, n28931, n28932, n28933,
         n28934, n28935, n28936, n28937, n28938, n28939, n28940, n28941,
         n28942, n28943, n28944, n28945, n28946, n28947, n28948, n28949,
         n28950, n28951, n28952, n28953, n28954, n28955, n28956, n28957,
         n28958, n28959, n28960, n28961, n28962, n28963, n28964, n28965,
         n28966, n28967, n28968, n28969, n28970, n28971, n28972, n28973,
         n28974, n28975, n28976, n28977, n28978, n28979, n28980, n28981,
         n28982, n28983, n28984, n28985, n28986, n28987, n28988, n28989,
         n28990, n28991, n28992, n28993, n28994, n28995, n28996, n28997,
         n28998, n28999, n29000, n29001, n29002, n29003, n29004, n29005,
         n29006, n29007, n29008, n29009, n29010, n29011, n29012, n29013,
         n29014, n29015, n29016, n29017, n29018, n29019, n29020, n29021,
         n29022, n29023, n29024, n29025, n29026, n29027, n29028, n29029,
         n29030, n29031, n29032, n29033, n29034, n29035, n29036, n29037,
         n29038, n29039, n29040, n29041, n29042, n29043, n29044, n29045,
         n29046, n29047, n29048, n29049, n29050, n29051, n29052, n29053,
         n29054, n29055, n29056, n29057, n29058, n29059, n29060, n29061,
         n29062, n29063, n29064, n29065, n29066, n29067, n29068, n29069,
         n29070, n29071, n29072, n29073, n29074, n29075, n29076, n29077,
         n29078, n29079, n29080, n29081, n29082, n29083, n29084, n29085,
         n29086, n29087, n29088, n29089, n29090, n29091, n29092, n29093,
         n29094, n29095, n29096, n29097, n29098, n29099, n29100, n29101,
         n29102, n29103, n29104, n29105, n29106, n29107, n29108, n29109,
         n29110, n29111, n29112, n29113, n29114, n29115, n29116, n29117,
         n29118, n29119, n29120, n29121, n29122, n29123, n29124, n29125,
         n29126, n29127, n29128, n29129, n29130, n29131, n29132, n29133,
         n29134, n29135, n29136, n29137, n29138, n29139, n29140, n29141,
         n29142, n29143, n29144, n29145, n29146, n29147, n29148, n29149,
         n29150, n29151, n29152, n29153, n29154, n29155, n29156, n29157,
         n29158, n29159, n29160, n29161, n29162, n29163, n29164, n29165,
         n29166, n29167, n29168, n29169, n29170, n29171, n29172, n29173,
         n29174, n29175, n29176, n29177, n29178, n29179, n29180, n29181,
         n29182, n29183, n29184, n29185, n29186, n29187, n29188, n29189,
         n29190, n29191, n29192, n29193, n29194, n29195, n29196, n29197,
         n29198, n29199, n29200, n29201, n29202, n29203, n29204, n29205,
         n29206, n29207, n29208, n29209, n29210, n29211, n29212, n29213,
         n29214, n29215, n29216, n29217, n29218, n29219, n29220, n29221,
         n29222, n29223, n29224, n29225, n29226, n29227, n29228, n29229,
         n29230, n29231, n29232, n29233, n29234, n29235, n29236, n29237,
         n29238, n29239, n29240, n29241, n29242, n29243, n29244, n29245,
         n29246, n29247, n29248, n29249, n29250, n29251, n29252, n29253,
         n29254, n29255, n29256, n29257, n29258, n29259, n29260, n29261,
         n29262, n29263, n29264, n29265, n29266, n29267, n29268, n29269,
         n29270, n29271, n29272, n29273, n29274, n29275, n29276, n29277,
         n29278, n29279, n29280, n29281, n29282, n29283, n29284, n29285,
         n29286, n29287, n29288, n29289, n29290, n29291, n29292, n29293,
         n29294, n29295, n29296, n29297, n29298, n29299, n29300, n29301,
         n29302, n29303, n29304, n29305, n29306, n29307, n29308, n29309,
         n29310, n29311, n29312, n29313, n29314, n29315, n29316, n29317,
         n29318, n29319, n29320, n29321, n29322, n29323, n29324, n29325,
         n29326, n29327, n29328, n29329, n29330, n29331, n29332, n29333,
         n29334, n29335, n29336, n29337, n29338, n29339, n29340, n29341,
         n29342, n29343, n29344, n29345, n29346, n29347, n29348, n29349,
         n29350, n29351, n29352, n29353, n29354, n29355, n29356, n29357,
         n29358, n29359, n29360, n29361, n29362, n29363, n29364, n29365,
         n29366, n29367, n29368, n29369, n29370, n29371, n29372, n29373,
         n29374, n29375, n29376, n29377, n29378, n29379, n29380, n29381,
         n29382, n29383, n29384, n29385, n29386, n29387, n29388, n29389,
         n29390, n29391, n29392, n29393, n29394, n29395, n29396, n29397,
         n29398, n29399, n29400, n29401, n29402, n29403, n29404, n29405,
         n29406, n29407, n29408, n29409, n29410, n29411, n29412, n29413,
         n29414, n29415, n29416, n29417, n29418, n29419, n29420, n29421,
         n29422, n29423, n29424, n29425, n29426, n29427, n29428, n29429,
         n29430, n29431, n29432, n29433, n29434, n29435, n29436, n29437,
         n29438, n29439, n29440, n29441, n29442, n29443, n29444, n29445,
         n29446, n29447, n29448, n29449, n29450, n29451, n29452, n29453,
         n29454, n29455, n29456, n29457, n29458, n29459, n29460, n29461,
         n29462, n29463, n29464, n29465, n29466, n29467, n29468, n29469,
         n29470, n29471, n29472, n29473, n29474, n29475, n29476, n29477,
         n29478, n29479, n29480, n29481, n29482, n29483, n29484, n29485,
         n29486, n29487, n29488, n29489, n29490, n29491, n29492, n29493,
         n29494, n29495, n29496, n29497, n29498, n29499, n29500, n29501,
         n29502, n29503, n29504, n29505, n29506, n29507, n29508, n29509,
         n29510, n29511, n29512, n29513, n29514, n29515, n29516, n29517,
         n29518, n29519, n29520, n29521, n29522, n29523, n29524, n29525,
         n29526, n29527, n29528, n29529, n29530, n29531, n29532, n29533,
         n29534, n29535, n29536, n29537, n29538, n29539, n29540, n29541,
         n29542, n29543, n29544, n29545, n29546, n29547, n29548, n29549,
         n29550, n29551, n29552, n29553, n29554, n29555, n29556, n29557,
         n29558, n29559, n29560, n29561, n29562, n29563, n29564, n29565,
         n29566, n29567, n29568, n29569, n29570, n29571, n29572, n29573,
         n29574, n29575, n29576, n29577, n29578, n29579, n29580, n29581,
         n29582, n29583, n29584, n29585, n29586, n29587, n29588, n29589,
         n29590, n29591, n29592, n29593, n29594, n29595, n29596, n29597,
         n29598, n29599, n29600, n29601, n29602, n29603, n29604, n29605,
         n29606, n29607, n29608, n29609, n29610, n29611, n29612, n29613,
         n29614, n29615, n29616, n29617, n29618, n29619, n29620, n29621,
         n29622, n29623, n29624, n29625, n29626, n29627, n29628, n29629,
         n29630, n29631, n29632, n29633, n29634, n29635, n29636, n29637,
         n29638, n29639, n29640, n29641, n29642, n29643, n29644, n29645,
         n29646, n29647, n29648, n29649, n29650, n29651, n29652, n29653,
         n29654, n29655, n29656, n29657, n29658, n29659, n29660, n29661,
         n29662, n29663, n29664, n29665, n29666, n29667, n29668, n29669,
         n29670, n29671, n29672, n29673, n29674, n29675, n29676, n29677,
         n29678, n29679, n29680, n29681, n29682, n29683, n29684, n29685,
         n29686, n29687, n29688, n29689, n29690, n29691, n29692, n29693,
         n29694, n29695, n29696, n29697, n29698, n29699, n29700, n29701,
         n29702, n29703, n29704, n29705, n29706, n29707, n29708, n29709,
         n29710, n29711, n29712, n29713, n29714, n29715, n29716, n29717,
         n29718, n29719, n29720, n29721, n29722, n29723, n29724, n29725,
         n29726, n29727, n29728, n29729, n29730, n29731, n29732, n29733,
         n29734, n29735, n29736, n29737, n29738, n29739, n29740, n29741,
         n29742, n29743, n29744, n29745, n29746, n29747, n29748, n29749,
         n29750, n29751, n29752, n29753, n29754, n29755, n29756, n29757,
         n29758, n29759, n29760, n29761, n29762, n29763, n29764, n29765,
         n29766, n29767, n29768, n29769, n29770, n29771, n29772, n29773,
         n29774, n29775, n29776, n29777, n29778, n29779, n29780, n29781,
         n29782, n29783, n29784, n29785, n29786, n29787, n29788, n29789,
         n29790, n29791, n29792, n29793, n29794, n29795, n29796, n29797,
         n29798, n29799, n29800, n29801, n29802, n29803, n29804, n29805,
         n29806, n29807, n29808, n29809, n29810, n29811, n29812, n29813,
         n29814, n29815, n29816, n29817, n29818, n29819, n29820, n29821,
         n29822, n29823, n29824, n29825, n29826, n29827, n29828, n29829,
         n29830, n29831, n29832, n29833, n29834, n29835, n29836, n29837,
         n29838, n29839, n29840, n29841, n29842, n29843, n29844, n29845,
         n29846, n29847, n29848, n29849, n29850, n29851, n29852, n29853,
         n29854, n29855, n29856, n29857, n29858, n29859, n29860, n29861,
         n29862, n29863, n29864, n29865, n29866, n29867, n29868, n29869,
         n29870, n29871, n29872, n29873, n29874, n29875, n29876, n29877,
         n29878, n29879, n29880, n29881, n29882, n29883, n29884, n29885,
         n29886, n29887, n29888, n29889, n29890, n29891, n29892, n29893,
         n29894, n29895, n29896, n29897, n29898, n29899, n29900, n29901,
         n29902, n29903, n29904, n29905, n29906, n29907, n29908, n29909,
         n29910, n29911, n29912, n29913, n29914, n29915, n29916, n29917,
         n29918, n29919, n29920, n29921, n29922, n29923, n29924, n29925,
         n29926, n29927, n29928, n29929, n29930, n29931, n29932, n29933,
         n29934, n29935, n29936, n29937, n29938, n29939, n29940, n29941,
         n29942, n29943, n29944, n29945, n29946, n29947, n29948, n29949,
         n29950, n29951, n29952, n29953, n29954, n29955, n29956, n29957,
         n29958, n29959, n29960, n29961, n29962, n29963, n29964, n29965,
         n29966, n29967, n29968, n29969, n29970, n29971, n29972, n29973,
         n29974, n29975, n29976, n29977, n29978, n29979, n29980, n29981,
         n29982, n29983, n29984, n29985, n29986, n29987, n29988, n29989,
         n29990, n29991, n29992, n29993, n29994, n29995, n29996, n29997,
         n29998, n29999, n30000, n30001, n30002, n30003, n30004, n30005,
         n30006, n30007, n30008, n30009, n30010, n30011, n30012, n30013,
         n30014, n30015, n30016, n30017, n30018, n30019, n30020, n30021,
         n30022, n30023, n30024, n30025, n30026, n30027, n30028, n30029,
         n30030, n30031, n30032, n30033, n30034, n30035, n30036, n30037,
         n30038, n30039, n30040, n30041, n30042, n30043, n30044, n30045,
         n30046, n30047, n30048, n30049, n30050, n30051, n30052, n30053,
         n30054, n30055, n30056, n30057, n30058, n30059, n30060, n30061,
         n30062, n30063, n30064, n30065, n30066, n30067, n30068, n30069,
         n30070, n30071, n30072, n30073, n30074, n30075, n30076, n30077,
         n30078, n30079, n30080, n30081, n30082, n30083, n30084, n30085,
         n30086, n30087, n30088, n30089, n30090, n30091, n30092, n30093,
         n30094, n30095, n30096, n30097, n30098, n30099, n30100, n30101,
         n30102, n30103, n30104, n30105, n30106, n30107, n30108, n30109,
         n30110, n30111, n30112, n30113, n30114, n30115, n30116, n30117,
         n30118, n30119, n30120, n30121, n30122, n30123, n30124, n30125,
         n30126, n30127, n30128, n30129, n30130, n30131, n30132, n30133,
         n30134, n30135, n30136, n30137, n30138, n30139, n30140, n30141,
         n30142, n30143, n30144, n30145, n30146, n30147, n30148, n30149,
         n30150, n30151, n30152, n30153, n30154, n30155, n30156, n30157,
         n30158, n30159, n30160, n30161, n30162, n30163, n30164, n30165,
         n30166, n30167, n30168, n30169, n30170, n30171, n30172, n30173,
         n30174, n30175, n30176, n30177, n30178, n30179, n30180, n30181,
         n30182, n30183, n30184, n30185, n30186, n30187, n30188, n30189,
         n30190, n30191, n30192, n30193, n30194, n30195, n30196, n30197,
         n30198, n30199, n30200, n30201, n30202, n30203, n30204, n30205,
         n30206, n30207, n30208, n30209, n30210, n30211, n30212, n30213,
         n30214, n30215, n30216, n30217, n30218, n30219, n30220, n30221,
         n30222, n30223, n30224, n30225, n30226, n30227, n30228, n30229,
         n30230, n30231, n30232, n30233, n30234, n30235, n30236, n30237,
         n30238, n30239, n30240, n30241, n30242, n30243, n30244, n30245,
         n30246, n30247, n30248, n30249, n30250, n30251, n30252, n30253,
         n30254, n30255, n30256, n30257, n30258, n30259, n30260, n30261,
         n30262, n30263, n30264, n30265, n30266, n30267, n30268, n30269,
         n30270, n30271, n30272, n30273, n30274, n30275, n30276, n30277,
         n30278, n30279, n30280, n30281, n30282, n30283, n30284, n30285,
         n30286, n30287, n30288, n30289, n30290, n30291, n30292, n30293,
         n30294, n30295, n30296, n30297, n30298, n30299, n30300, n30301,
         n30302, n30303, n30304, n30305, n30306, n30307, n30308, n30309,
         n30310, n30311, n30312, n30313, n30314, n30315, n30316, n30317,
         n30318, n30319, n30320, n30321, n30322, n30323, n30324, n30325,
         n30326, n30327, n30328, n30329, n30330, n30331, n30332, n30333,
         n30334, n30335, n30336, n30337, n30338, n30339, n30340, n30341,
         n30342, n30343, n30344, n30345, n30346, n30347, n30348, n30349,
         n30350, n30351, n30352, n30353, n30354, n30355, n30356, n30357,
         n30358, n30359, n30360, n30361, n30362, n30363, n30364, n30365,
         n30366, n30367, n30368, n30369, n30370, n30371, n30372, n30373,
         n30374, n30375, n30376, n30377, n30378, n30379, n30380, n30381,
         n30382, n30383, n30384, n30385, n30386, n30387, n30388, n30389,
         n30390, n30391, n30392, n30393, n30394, n30395, n30396, n30397,
         n30398, n30399, n30400, n30401, n30402, n30403, n30404, n30405,
         n30406, n30407, n30408, n30409, n30410, n30411, n30412, n30413,
         n30414, n30415, n30416, n30417, n30418, n30419, n30420, n30421,
         n30422, n30423, n30424, n30425, n30426, n30427, n30428, n30429,
         n30430, n30431, n30432, n30433, n30434, n30435, n30436, n30437,
         n30438, n30439, n30440, n30441, n30442, n30443, n30444, n30445,
         n30446, n30447, n30448, n30449, n30450, n30451, n30452, n30453,
         n30454, n30455, n30456, n30457, n30458, n30459, n30460, n30461,
         n30462, n30463, n30464, n30465, n30466, n30467, n30468, n30469,
         n30470, n30471, n30472, n30473, n30474, n30475, n30476, n30477,
         n30478, n30479, n30480, n30481, n30482, n30483, n30484, n30485,
         n30486, n30487, n30488, n30489, n30490, n30491, n30492, n30493,
         n30494, n30495, n30496, n30497, n30498, n30499, n30500, n30501,
         n30502, n30503, n30504, n30505, n30506, n30507, n30508, n30509,
         n30510, n30511, n30512, n30513, n30514, n30515, n30516, n30517,
         n30518, n30519, n30520, n30521, n30522, n30523, n30524, n30525,
         n30526, n30527, n30528, n30529, n30530, n30531, n30532, n30533,
         n30534, n30535, n30536, n30537, n30538, n30539, n30540, n30541,
         n30542, n30543, n30544, n30545, n30546, n30547, n30548, n30549,
         n30550, n30551, n30552, n30553, n30554, n30555, n30556, n30557,
         n30558, n30559, n30560, n30561, n30562, n30563, n30564, n30565,
         n30566, n30567, n30568, n30569, n30570, n30571, n30572, n30573,
         n30574, n30575, n30576, n30577, n30578, n30579, n30580, n30581,
         n30582, n30583, n30584, n30585, n30586, n30587, n30588, n30589,
         n30590, n30591, n30592, n30593, n30594, n30595, n30596, n30597,
         n30598, n30599, n30600, n30601, n30602, n30603, n30604, n30605,
         n30606, n30607, n30608, n30609, n30610, n30611, n30612, n30613,
         n30614, n30615, n30616, n30617, n30618, n30619, n30620, n30621,
         n30622, n30623, n30624, n30625, n30626, n30627, n30628, n30629,
         n30630, n30631, n30632, n30633, n30634, n30635, n30636, n30637,
         n30638, n30639, n30640, n30641, n30642, n30643, n30644, n30645,
         n30646, n30647, n30648, n30649, n30650, n30651, n30652, n30653,
         n30654, n30655, n30656, n30657, n30658, n30659, n30660, n30661,
         n30662, n30663, n30664, n30665, n30666, n30667, n30668, n30669,
         n30670, n30671, n30672, n30673, n30674, n30675, n30676, n30677,
         n30678, n30679, n30680, n30681, n30682, n30683, n30684, n30685,
         n30686, n30687, n30688, n30689, n30690, n30691, n30692, n30693,
         n30694, n30695, n30696, n30697, n30698, n30699, n30700, n30701,
         n30702, n30703, n30704, n30705, n30706, n30707, n30708, n30709,
         n30710, n30711, n30712, n30713, n30714, n30715, n30716, n30717,
         n30718, n30719, n30720, n30721, n30722, n30723, n30724, n30725,
         n30726, n30727, n30728, n30729, n30730, n30731, n30732, n30733,
         n30734, n30735, n30736, n30737, n30738, n30739, n30740, n30741,
         n30742, n30743, n30744, n30745, n30746, n30747, n30748, n30749,
         n30750, n30751, n30752, n30753, n30754, n30755, n30756, n30757,
         n30758, n30759, n30760, n30761, n30762, n30763, n30764, n30765,
         n30766, n30767, n30768, n30769, n30770, n30771, n30772, n30773,
         n30774, n30775, n30776, n30777, n30778, n30779, n30780, n30781,
         n30782, n30783, n30784, n30785, n30786, n30787, n30788, n30789,
         n30790, n30791, n30792, n30793, n30794, n30795, n30796, n30797,
         n30798, n30799, n30800, n30801, n30802, n30803, n30804, n30805,
         n30806, n30807, n30808, n30809, n30810, n30811, n30812, n30813,
         n30814, n30815, n30816, n30817, n30818, n30819, n30820, n30821,
         n30822, n30823, n30824, n30825, n30826, n30827, n30828, n30829,
         n30830, n30831, n30832, n30833, n30834, n30835, n30836, n30837,
         n30838, n30839, n30840, n30841, n30842, n30843, n30844, n30845,
         n30846, n30847, n30848, n30849, n30850, n30851, n30852, n30853,
         n30854, n30855, n30856, n30857, n30858, n30859, n30860, n30861,
         n30862, n30863, n30864, n30865, n30866, n30867, n30868, n30869,
         n30870, n30871, n30872, n30873, n30874, n30875, n30876, n30877,
         n30878, n30879, n30880, n30881, n30882, n30883, n30884, n30885,
         n30886, n30887, n30888, n30889, n30890, n30891, n30892, n30893,
         n30894, n30895, n30896, n30897, n30898, n30899, n30900, n30901,
         n30902, n30903, n30904, n30905, n30906, n30907, n30908, n30909,
         n30910, n30911, n30912, n30913, n30914, n30915, n30916, n30917,
         n30918, n30919, n30920, n30921, n30922, n30923, n30924, n30925,
         n30926, n30927, n30928, n30929, n30930, n30931, n30932, n30933,
         n30934, n30935, n30936, n30937, n30938, n30939, n30940, n30941,
         n30942, n30943, n30944, n30945, n30946, n30947, n30948, n30949,
         n30950, n30951, n30952, n30953, n30954, n30955, n30956, n30957,
         n30958, n30959, n30960, n30961, n30962, n30963, n30964, n30965,
         n30966, n30967, n30968, n30969, n30970, n30971, n30972, n30973,
         n30974, n30975, n30976, n30977, n30978, n30979, n30980, n30981,
         n30982, n30983, n30984, n30985, n30986, n30987, n30988, n30989,
         n30990, n30991, n30992, n30993, n30994, n30995, n30996, n30997,
         n30998, n30999, n31000, n31001, n31002, n31003, n31004, n31005,
         n31006, n31007, n31008, n31009, n31010, n31011, n31012, n31013,
         n31014, n31015, n31016, n31017, n31018, n31019, n31020, n31021,
         n31022, n31023, n31024, n31025, n31026, n31027, n31028, n31029,
         n31030, n31031, n31032, n31033, n31034, n31035, n31036, n31037,
         n31038, n31039, n31040, n31041, n31042, n31043, n31044, n31045,
         n31046, n31047, n31048, n31049, n31050, n31051, n31052, n31053,
         n31054, n31055, n31056, n31057, n31058, n31059, n31060, n31061,
         n31062, n31063, n31064, n31065, n31066, n31067, n31068, n31069,
         n31070, n31071, n31072, n31073, n31074, n31075, n31076, n31077,
         n31078, n31079, n31080, n31081, n31082, n31083, n31084, n31085,
         n31086, n31087, n31088, n31089, n31090, n31091, n31092, n31093,
         n31094, n31095, n31096, n31097, n31098, n31099, n31100, n31101,
         n31102, n31103, n31104, n31105, n31106, n31107, n31108, n31109,
         n31110, n31111, n31112, n31113, n31114, n31115, n31116, n31117,
         n31118, n31119, n31120, n31121, n31122, n31123, n31124, n31125,
         n31126, n31127, n31128, n31129, n31130, n31131, n31132, n31133,
         n31134, n31135, n31136, n31137, n31138, n31139, n31140, n31141,
         n31142, n31143, n31144, n31145, n31146, n31147, n31148, n31149,
         n31150, n31151, n31152, n31153, n31154, n31155, n31156, n31157,
         n31158, n31159, n31160, n31161, n31162, n31163, n31164, n31165,
         n31166, n31167, n31168, n31169, n31170, n31171, n31172, n31173,
         n31174, n31175, n31176, n31177, n31178, n31179, n31180, n31181,
         n31182, n31183, n31184, n31185, n31186, n31187, n31188, n31189,
         n31190, n31191, n31192, n31193, n31194, n31195, n31196, n31197,
         n31198, n31199, n31200, n31201, n31202, n31203, n31204, n31205,
         n31206, n31207, n31208, n31209, n31210, n31211, n31212, n31213,
         n31214, n31215, n31216, n31217, n31218, n31219, n31220, n31221,
         n31222, n31223, n31224, n31225, n31226, n31227, n31228, n31229,
         n31230, n31231, n31232, n31233, n31234, n31235, n31236, n31237,
         n31238, n31239, n31240, n31241, n31242, n31243, n31244, n31245,
         n31246, n31247, n31248, n31249, n31250, n31251, n31252, n31253,
         n31254, n31255, n31256, n31257, n31258, n31259, n31260, n31261,
         n31262, n31263, n31264, n31265, n31266, n31267, n31268, n31269,
         n31270, n31271, n31272, n31273, n31274, n31275, n31276, n31277,
         n31278, n31279, n31280, n31281, n31282, n31283, n31284, n31285,
         n31286, n31287, n31288, n31289, n31290, n31291, n31292, n31293,
         n31294, n31295, n31296, n31297, n31298, n31299, n31300, n31301,
         n31302, n31303, n31304, n31305, n31306, n31307, n31308, n31309,
         n31310, n31311, n31312, n31313, n31314, n31315, n31316, n31317,
         n31318, n31319, n31320, n31321, n31322, n31323, n31324, n31325,
         n31326, n31327, n31328, n31329, n31330, n31331, n31332, n31333,
         n31334, n31335, n31336, n31337, n31338, n31339, n31340, n31341,
         n31342, n31343, n31344, n31345, n31346, n31347, n31348, n31349,
         n31350, n31351, n31352, n31353, n31354, n31355, n31356, n31357,
         n31358, n31359, n31360, n31361, n31362, n31363, n31364, n31365,
         n31366, n31367, n31368, n31369, n31370, n31371, n31372, n31373,
         n31374, n31375, n31376, n31377, n31378, n31379, n31380, n31381,
         n31382, n31383, n31384, n31385, n31386, n31387, n31388, n31389,
         n31390, n31391, n31392, n31393, n31394, n31395, n31396, n31397,
         n31398, n31399, n31400, n31401, n31402, n31403, n31404, n31405,
         n31406, n31407, n31408, n31409, n31410, n31411, n31412, n31413,
         n31414, n31415, n31416, n31417, n31418, n31419, n31420, n31421,
         n31422, n31423, n31424, n31425, n31426, n31427, n31428, n31429,
         n31430, n31431, n31432, n31433, n31434, n31435, n31436, n31437,
         n31438, n31439, n31440, n31441, n31442, n31443, n31444, n31445,
         n31446, n31447, n31448, n31449, n31450, n31451, n31452, n31453,
         n31454, n31455, n31456, n31457, n31458, n31459, n31460, n31461,
         n31462, n31463, n31464, n31465, n31466, n31467, n31468, n31469,
         n31470, n31471, n31472, n31473, n31474, n31475, n31476, n31477,
         n31478, n31479, n31480, n31481, n31482, n31483, n31484, n31485,
         n31486, n31487, n31488, n31489, n31490, n31491, n31492, n31493,
         n31494, n31495, n31496, n31497, n31498, n31499, n31500, n31501,
         n31502, n31503, n31504, n31505, n31506, n31507, n31508, n31509,
         n31510, n31511, n31512, n31513, n31514, n31515, n31516, n31517,
         n31518, n31519, n31520, n31521, n31522, n31523, n31524, n31525,
         n31526, n31527, n31528, n31529, n31530, n31531, n31532, n31533,
         n31534, n31535, n31536, n31537, n31538, n31539, n31540, n31541,
         n31542, n31543, n31544, n31545, n31546, n31547, n31548, n31549,
         n31550, n31551, n31552, n31553, n31554, n31555, n31556, n31557,
         n31558, n31559, n31560, n31561, n31562, n31563, n31564, n31565,
         n31566, n31567, n31568, n31569, n31570, n31571, n31572, n31573,
         n31574, n31575, n31576, n31577, n31578, n31579, n31580, n31581,
         n31582, n31583, n31584, n31585, n31586, n31587, n31588, n31589,
         n31590, n31591, n31592, n31593, n31594, n31595, n31596, n31597,
         n31598, n31599, n31600, n31601, n31602, n31603, n31604, n31605,
         n31606, n31607, n31608, n31609, n31610, n31611, n31612, n31613,
         n31614, n31615, n31616, n31617, n31618, n31619, n31620, n31621,
         n31622, n31623, n31624, n31625, n31626, n31627, n31628, n31629,
         n31630, n31631, n31632, n31633, n31634, n31635, n31636, n31637,
         n31638, n31639, n31640, n31641, n31642, n31643, n31644, n31645,
         n31646, n31647, n31648, n31649, n31650, n31651, n31652, n31653,
         n31654, n31655, n31656, n31657, n31658, n31659, n31660, n31661,
         n31662, n31663, n31664, n31665, n31666, n31667, n31668, n31669,
         n31670, n31671, n31672, n31673, n31674, n31675, n31676, n31677,
         n31678, n31679, n31680, n31681, n31682, n31683, n31684, n31685,
         n31686, n31687, n31688, n31689, n31690, n31691, n31692, n31693,
         n31694, n31695, n31696, n31697, n31698, n31699, n31700, n31701,
         n31702, n31703, n31704, n31705, n31706, n31707, n31708, n31709,
         n31710, n31711, n31712, n31713, n31714, n31715, n31716, n31717,
         n31718, n31719, n31720, n31721, n31722, n31723, n31724, n31725,
         n31726, n31727, n31728, n31729, n31730, n31731, n31732, n31733,
         n31734, n31735, n31736, n31737, n31738, n31739, n31740, n31741,
         n31742, n31743, n31744, n31745, n31746, n31747, n31748, n31749,
         n31750, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
         n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
         n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
         n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
         n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
         n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
         n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
         n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
         n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
         n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471,
         n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
         n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491,
         n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501,
         n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
         n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
         n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531,
         n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541,
         n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551,
         n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561,
         n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571,
         n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581,
         n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591,
         n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
         n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611,
         n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
         n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
         n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
         n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651,
         n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661,
         n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671,
         n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
         n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691,
         n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701,
         n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711,
         n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721,
         n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731,
         n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741,
         n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751,
         n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761,
         n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771,
         n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
         n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791,
         n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801,
         n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811,
         n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821,
         n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831,
         n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841,
         n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851,
         n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861,
         n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871,
         n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881,
         n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891,
         n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901,
         n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911,
         n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921,
         n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931,
         n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941,
         n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951,
         n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961,
         n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971,
         n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981,
         n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991,
         n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001,
         n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011,
         n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021,
         n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031,
         n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041,
         n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051,
         n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061,
         n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071,
         n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081,
         n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091,
         n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101,
         n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111,
         n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121,
         n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131,
         n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141,
         n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
         n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
         n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2194,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
         n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
         n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
         n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
         n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
         n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
         n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
         n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
         n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
         n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
         n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
         n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
         n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
         n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
         n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
         n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
         n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
         n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
         n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
         n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
         n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
         n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653,
         n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
         n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
         n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
         n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693,
         n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
         n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
         n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723,
         n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733,
         n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743,
         n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
         n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
         n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773,
         n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
         n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
         n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
         n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
         n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
         n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
         n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843,
         n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
         n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
         n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
         n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883,
         n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
         n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
         n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
         n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923,
         n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933,
         n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
         n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953,
         n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
         n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973,
         n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
         n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
         n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
         n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013,
         n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023,
         n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033,
         n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
         n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
         n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
         n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
         n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
         n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
         n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
         n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
         n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
         n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
         n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
         n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
         n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
         n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
         n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
         n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
         n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
         n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
         n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
         n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
         n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
         n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
         n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
         n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
         n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
         n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
         n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
         n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
         n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
         n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
         n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
         n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
         n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
         n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
         n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
         n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
         n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
         n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843,
         n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853,
         n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863,
         n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
         n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
         n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
         n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
         n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
         n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
         n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933,
         n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943,
         n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953,
         n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963,
         n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973,
         n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983,
         n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993,
         n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003,
         n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013,
         n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023,
         n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033,
         n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043,
         n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053,
         n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063,
         n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073,
         n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083,
         n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
         n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103,
         n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113,
         n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123,
         n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133,
         n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143,
         n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153,
         n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163,
         n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173,
         n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183,
         n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193,
         n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203,
         n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213,
         n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223,
         n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233,
         n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243,
         n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
         n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
         n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273,
         n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
         n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
         n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
         n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
         n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
         n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
         n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
         n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
         n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
         n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
         n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
         n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
         n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083,
         n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
         n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
         n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
         n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
         n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
         n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
         n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
         n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
         n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
         n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
         n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
         n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
         n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
         n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
         n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233,
         n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
         n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
         n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
         n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
         n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
         n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
         n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
         n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
         n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
         n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
         n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
         n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
         n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
         n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
         n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
         n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
         n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
         n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
         n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
         n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
         n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
         n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
         n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
         n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
         n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
         n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
         n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
         n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803,
         n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
         n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823,
         n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833,
         n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843,
         n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853,
         n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
         n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873,
         n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883,
         n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893,
         n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903,
         n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
         n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
         n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
         n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
         n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
         n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
         n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
         n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
         n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
         n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
         n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
         n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
         n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
         n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
         n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
         n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
         n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
         n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
         n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
         n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
         n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
         n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
         n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
         n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
         n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
         n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
         n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
         n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
         n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
         n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
         n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
         n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
         n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
         n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
         n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
         n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
         n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
         n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
         n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
         n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603,
         n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
         n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
         n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
         n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
         n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
         n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
         n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
         n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
         n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
         n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
         n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
         n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
         n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
         n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
         n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
         n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
         n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
         n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803,
         n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813,
         n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
         n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
         n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
         n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853,
         n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
         n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873,
         n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883,
         n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893,
         n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903,
         n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913,
         n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923,
         n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933,
         n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943,
         n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
         n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973,
         n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983,
         n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993,
         n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
         n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
         n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023,
         n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033,
         n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043,
         n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053,
         n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063,
         n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073,
         n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083,
         n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093,
         n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103,
         n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113,
         n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123,
         n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133,
         n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143,
         n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153,
         n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163,
         n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173,
         n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183,
         n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193,
         n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203,
         n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213,
         n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
         n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233,
         n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243,
         n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253,
         n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263,
         n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273,
         n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283,
         n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293,
         n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303,
         n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313,
         n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323,
         n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333,
         n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343,
         n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353,
         n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363,
         n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373,
         n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383,
         n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393,
         n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403,
         n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413,
         n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423,
         n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433,
         n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443,
         n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453,
         n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463,
         n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473,
         n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483,
         n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493,
         n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503,
         n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513,
         n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523,
         n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533,
         n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543,
         n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553,
         n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563,
         n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573,
         n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583,
         n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593,
         n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603,
         n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613,
         n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623,
         n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633,
         n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643,
         n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653,
         n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663,
         n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673,
         n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683,
         n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693,
         n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703,
         n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713,
         n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723,
         n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733,
         n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743,
         n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753,
         n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763,
         n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773,
         n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783,
         n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793,
         n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803,
         n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813,
         n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823,
         n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833,
         n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843,
         n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853,
         n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863,
         n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873,
         n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883,
         n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893,
         n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903,
         n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913,
         n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923,
         n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933,
         n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943,
         n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953,
         n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963,
         n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973,
         n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983,
         n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993,
         n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003,
         n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013,
         n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023,
         n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033,
         n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043,
         n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053,
         n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063,
         n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073,
         n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083,
         n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093,
         n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103,
         n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113,
         n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123,
         n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133,
         n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143,
         n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153,
         n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163,
         n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173,
         n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183,
         n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193,
         n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203,
         n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213,
         n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223,
         n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233,
         n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243,
         n8244, n8245;
  tri   [31:0] do;
  assign test_so8 = N61;
  assign test_so7 = \mem3[242][27] ;
  assign test_so6 = \mem3[77][29] ;
  assign test_so5 = \mem2[168][23] ;
  assign test_so4 = \mem2[4][17] ;
  assign test_so3 = \mem1[95][11] ;
  assign test_so2 = \mem0[186][5] ;
  assign test_so1 = \mem0[21][7] ;

  SDFFX1 \raddr_reg[7]  ( .D(n10411), .SI(N60), .SE(test_se), .CLK(n1737), .Q(
        N61), .QN(n31745) );
  SDFFX1 \raddr_reg[6]  ( .D(n10409), .SI(N59), .SE(test_se), .CLK(n1737), .Q(
        N60), .QN(n31746) );
  SDFFX1 \raddr_reg[5]  ( .D(n10407), .SI(N58), .SE(test_se), .CLK(n1737), .Q(
        N59), .QN(n31747) );
  SDFFX1 \raddr_reg[4]  ( .D(n10405), .SI(N57), .SE(test_se), .CLK(n1737), .Q(
        N58), .QN(n31748) );
  SDFFX1 \raddr_reg[3]  ( .D(n10403), .SI(N56), .SE(test_se), .CLK(n1737), .Q(
        N57), .QN(n31749) );
  SDFFX1 \raddr_reg[2]  ( .D(n10401), .SI(N55), .SE(test_se), .CLK(n1737), .Q(
        N56), .QN(n21496) );
  SDFFX1 \raddr_reg[1]  ( .D(n10399), .SI(N54), .SE(test_se), .CLK(n1737), .Q(
        N55), .QN(n21497) );
  SDFFX1 \raddr_reg[0]  ( .D(n10397), .SI(\mem3[255][31] ), .SE(test_se), 
        .CLK(n1737), .Q(N54), .QN(n31750) );
  SDFFX1 \mem0_reg[255][7]  ( .D(n18603), .SI(\mem0[255][6] ), .SE(test_se), 
        .CLK(n1581), .Q(\mem0[255][7] ), .QN(n23553) );
  SDFFX1 \mem0_reg[255][6]  ( .D(n18602), .SI(\mem0[255][5] ), .SE(test_se), 
        .CLK(n1581), .Q(\mem0[255][6] ), .QN(n23554) );
  SDFFX1 \mem0_reg[255][5]  ( .D(n18601), .SI(\mem0[255][4] ), .SE(test_se), 
        .CLK(n1581), .Q(\mem0[255][5] ), .QN(n23555) );
  SDFFX1 \mem0_reg[255][4]  ( .D(n18600), .SI(\mem0[255][3] ), .SE(test_se), 
        .CLK(n1581), .Q(\mem0[255][4] ), .QN(n23556) );
  SDFFX1 \mem0_reg[255][3]  ( .D(n18599), .SI(\mem0[255][2] ), .SE(test_se), 
        .CLK(n1581), .Q(\mem0[255][3] ), .QN(n23557) );
  SDFFX1 \mem0_reg[255][2]  ( .D(n18598), .SI(\mem0[255][1] ), .SE(test_se), 
        .CLK(n1581), .Q(\mem0[255][2] ), .QN(n23558) );
  SDFFX1 \mem0_reg[255][1]  ( .D(n18597), .SI(\mem0[255][0] ), .SE(test_se), 
        .CLK(n1581), .Q(\mem0[255][1] ), .QN(n23559) );
  SDFFX1 \mem0_reg[255][0]  ( .D(n18596), .SI(\mem0[254][7] ), .SE(test_se), 
        .CLK(n1581), .Q(\mem0[255][0] ), .QN(n23560) );
  SDFFX1 \mem0_reg[254][7]  ( .D(n18595), .SI(\mem0[254][6] ), .SE(test_se), 
        .CLK(n1581), .Q(\mem0[254][7] ), .QN(n23561) );
  SDFFX1 \mem0_reg[254][6]  ( .D(n18594), .SI(\mem0[254][5] ), .SE(test_se), 
        .CLK(n1581), .Q(\mem0[254][6] ), .QN(n23562) );
  SDFFX1 \mem0_reg[254][5]  ( .D(n18593), .SI(\mem0[254][4] ), .SE(test_se), 
        .CLK(n1582), .Q(\mem0[254][5] ), .QN(n23563) );
  SDFFX1 \mem0_reg[254][4]  ( .D(n18592), .SI(\mem0[254][3] ), .SE(test_se), 
        .CLK(n1582), .Q(\mem0[254][4] ), .QN(n23564) );
  SDFFX1 \mem0_reg[254][3]  ( .D(n18591), .SI(\mem0[254][2] ), .SE(test_se), 
        .CLK(n1582), .Q(\mem0[254][3] ), .QN(n23565) );
  SDFFX1 \mem0_reg[254][2]  ( .D(n18590), .SI(\mem0[254][1] ), .SE(test_se), 
        .CLK(n1582), .Q(\mem0[254][2] ), .QN(n23566) );
  SDFFX1 \mem0_reg[254][1]  ( .D(n18589), .SI(\mem0[254][0] ), .SE(test_se), 
        .CLK(n1582), .Q(\mem0[254][1] ), .QN(n23567) );
  SDFFX1 \mem0_reg[254][0]  ( .D(n18588), .SI(\mem0[253][7] ), .SE(test_se), 
        .CLK(n1582), .Q(\mem0[254][0] ), .QN(n23568) );
  SDFFX1 \mem0_reg[253][7]  ( .D(n18587), .SI(\mem0[253][6] ), .SE(test_se), 
        .CLK(n1582), .Q(\mem0[253][7] ), .QN(n23569) );
  SDFFX1 \mem0_reg[253][6]  ( .D(n18586), .SI(\mem0[253][5] ), .SE(test_se), 
        .CLK(n1582), .Q(\mem0[253][6] ), .QN(n23570) );
  SDFFX1 \mem0_reg[253][5]  ( .D(n18585), .SI(\mem0[253][4] ), .SE(test_se), 
        .CLK(n1582), .Q(\mem0[253][5] ), .QN(n23571) );
  SDFFX1 \mem0_reg[253][4]  ( .D(n18584), .SI(\mem0[253][3] ), .SE(test_se), 
        .CLK(n1582), .Q(\mem0[253][4] ), .QN(n23572) );
  SDFFX1 \mem0_reg[253][3]  ( .D(n18583), .SI(\mem0[253][2] ), .SE(test_se), 
        .CLK(n1582), .Q(\mem0[253][3] ), .QN(n23573) );
  SDFFX1 \mem0_reg[253][2]  ( .D(n18582), .SI(\mem0[253][1] ), .SE(test_se), 
        .CLK(n1582), .Q(\mem0[253][2] ), .QN(n23574) );
  SDFFX1 \mem0_reg[253][1]  ( .D(n18581), .SI(\mem0[253][0] ), .SE(test_se), 
        .CLK(n1583), .Q(\mem0[253][1] ), .QN(n23575) );
  SDFFX1 \mem0_reg[253][0]  ( .D(n18580), .SI(\mem0[252][7] ), .SE(test_se), 
        .CLK(n1583), .Q(\mem0[253][0] ), .QN(n23576) );
  SDFFX1 \mem0_reg[252][7]  ( .D(n18579), .SI(\mem0[252][6] ), .SE(test_se), 
        .CLK(n1583), .Q(\mem0[252][7] ), .QN(n23577) );
  SDFFX1 \mem0_reg[252][6]  ( .D(n18578), .SI(\mem0[252][5] ), .SE(test_se), 
        .CLK(n1583), .Q(\mem0[252][6] ), .QN(n23578) );
  SDFFX1 \mem0_reg[252][5]  ( .D(n18577), .SI(\mem0[252][4] ), .SE(test_se), 
        .CLK(n1583), .Q(\mem0[252][5] ), .QN(n23579) );
  SDFFX1 \mem0_reg[252][4]  ( .D(n18576), .SI(\mem0[252][3] ), .SE(test_se), 
        .CLK(n1583), .Q(\mem0[252][4] ), .QN(n23580) );
  SDFFX1 \mem0_reg[252][3]  ( .D(n18575), .SI(\mem0[252][2] ), .SE(test_se), 
        .CLK(n1583), .Q(\mem0[252][3] ), .QN(n23581) );
  SDFFX1 \mem0_reg[252][2]  ( .D(n18574), .SI(\mem0[252][1] ), .SE(test_se), 
        .CLK(n1583), .Q(\mem0[252][2] ), .QN(n23582) );
  SDFFX1 \mem0_reg[252][1]  ( .D(n18573), .SI(\mem0[252][0] ), .SE(test_se), 
        .CLK(n1583), .Q(\mem0[252][1] ), .QN(n23583) );
  SDFFX1 \mem0_reg[252][0]  ( .D(n18572), .SI(\mem0[251][7] ), .SE(test_se), 
        .CLK(n1583), .Q(\mem0[252][0] ), .QN(n23584) );
  SDFFX1 \mem0_reg[251][7]  ( .D(n18571), .SI(\mem0[251][6] ), .SE(test_se), 
        .CLK(n1583), .Q(\mem0[251][7] ), .QN(n23585) );
  SDFFX1 \mem0_reg[251][6]  ( .D(n18570), .SI(\mem0[251][5] ), .SE(test_se), 
        .CLK(n1583), .Q(\mem0[251][6] ), .QN(n23586) );
  SDFFX1 \mem0_reg[251][5]  ( .D(n18569), .SI(\mem0[251][4] ), .SE(test_se), 
        .CLK(n1584), .Q(\mem0[251][5] ), .QN(n23587) );
  SDFFX1 \mem0_reg[251][4]  ( .D(n18568), .SI(\mem0[251][3] ), .SE(test_se), 
        .CLK(n1584), .Q(\mem0[251][4] ), .QN(n23588) );
  SDFFX1 \mem0_reg[251][3]  ( .D(n18567), .SI(\mem0[251][2] ), .SE(test_se), 
        .CLK(n1584), .Q(\mem0[251][3] ), .QN(n23589) );
  SDFFX1 \mem0_reg[251][2]  ( .D(n18566), .SI(\mem0[251][1] ), .SE(test_se), 
        .CLK(n1584), .Q(\mem0[251][2] ), .QN(n23590) );
  SDFFX1 \mem0_reg[251][1]  ( .D(n18565), .SI(\mem0[251][0] ), .SE(test_se), 
        .CLK(n1584), .Q(\mem0[251][1] ), .QN(n23591) );
  SDFFX1 \mem0_reg[251][0]  ( .D(n18564), .SI(\mem0[250][7] ), .SE(test_se), 
        .CLK(n1584), .Q(\mem0[251][0] ), .QN(n23592) );
  SDFFX1 \mem0_reg[250][7]  ( .D(n18563), .SI(\mem0[250][6] ), .SE(test_se), 
        .CLK(n1584), .Q(\mem0[250][7] ), .QN(n23593) );
  SDFFX1 \mem0_reg[250][6]  ( .D(n18562), .SI(\mem0[250][5] ), .SE(test_se), 
        .CLK(n1584), .Q(\mem0[250][6] ), .QN(n23594) );
  SDFFX1 \mem0_reg[250][5]  ( .D(n18561), .SI(\mem0[250][4] ), .SE(test_se), 
        .CLK(n1584), .Q(\mem0[250][5] ), .QN(n23595) );
  SDFFX1 \mem0_reg[250][4]  ( .D(n18560), .SI(\mem0[250][3] ), .SE(test_se), 
        .CLK(n1584), .Q(\mem0[250][4] ), .QN(n23596) );
  SDFFX1 \mem0_reg[250][3]  ( .D(n18559), .SI(\mem0[250][2] ), .SE(test_se), 
        .CLK(n1584), .Q(\mem0[250][3] ), .QN(n23597) );
  SDFFX1 \mem0_reg[250][2]  ( .D(n18558), .SI(\mem0[250][1] ), .SE(test_se), 
        .CLK(n1584), .Q(\mem0[250][2] ), .QN(n23598) );
  SDFFX1 \mem0_reg[250][1]  ( .D(n18557), .SI(\mem0[250][0] ), .SE(test_se), 
        .CLK(n1585), .Q(\mem0[250][1] ), .QN(n23599) );
  SDFFX1 \mem0_reg[250][0]  ( .D(n18556), .SI(\mem0[249][7] ), .SE(test_se), 
        .CLK(n1585), .Q(\mem0[250][0] ), .QN(n23600) );
  SDFFX1 \mem0_reg[249][7]  ( .D(n18555), .SI(\mem0[249][6] ), .SE(test_se), 
        .CLK(n1585), .Q(\mem0[249][7] ), .QN(n23601) );
  SDFFX1 \mem0_reg[249][6]  ( .D(n18554), .SI(\mem0[249][5] ), .SE(test_se), 
        .CLK(n1585), .Q(\mem0[249][6] ), .QN(n23602) );
  SDFFX1 \mem0_reg[249][5]  ( .D(n18553), .SI(\mem0[249][4] ), .SE(test_se), 
        .CLK(n1585), .Q(\mem0[249][5] ), .QN(n23603) );
  SDFFX1 \mem0_reg[249][4]  ( .D(n18552), .SI(\mem0[249][3] ), .SE(test_se), 
        .CLK(n1585), .Q(\mem0[249][4] ), .QN(n23604) );
  SDFFX1 \mem0_reg[249][3]  ( .D(n18551), .SI(\mem0[249][2] ), .SE(test_se), 
        .CLK(n1585), .Q(\mem0[249][3] ), .QN(n23605) );
  SDFFX1 \mem0_reg[249][2]  ( .D(n18550), .SI(\mem0[249][1] ), .SE(test_se), 
        .CLK(n1585), .Q(\mem0[249][2] ), .QN(n23606) );
  SDFFX1 \mem0_reg[249][1]  ( .D(n18549), .SI(\mem0[249][0] ), .SE(test_se), 
        .CLK(n1585), .Q(\mem0[249][1] ), .QN(n23607) );
  SDFFX1 \mem0_reg[249][0]  ( .D(n18548), .SI(\mem0[248][7] ), .SE(test_se), 
        .CLK(n1585), .Q(\mem0[249][0] ), .QN(n23608) );
  SDFFX1 \mem0_reg[248][7]  ( .D(n18547), .SI(\mem0[248][6] ), .SE(test_se), 
        .CLK(n1585), .Q(\mem0[248][7] ), .QN(n23609) );
  SDFFX1 \mem0_reg[248][6]  ( .D(n18546), .SI(\mem0[248][5] ), .SE(test_se), 
        .CLK(n1585), .Q(\mem0[248][6] ), .QN(n23610) );
  SDFFX1 \mem0_reg[248][5]  ( .D(n18545), .SI(\mem0[248][4] ), .SE(test_se), 
        .CLK(n1586), .Q(\mem0[248][5] ), .QN(n23611) );
  SDFFX1 \mem0_reg[248][4]  ( .D(n18544), .SI(\mem0[248][3] ), .SE(test_se), 
        .CLK(n1586), .Q(\mem0[248][4] ), .QN(n23612) );
  SDFFX1 \mem0_reg[248][3]  ( .D(n18543), .SI(\mem0[248][2] ), .SE(test_se), 
        .CLK(n1586), .Q(\mem0[248][3] ), .QN(n23613) );
  SDFFX1 \mem0_reg[248][2]  ( .D(n18542), .SI(\mem0[248][1] ), .SE(test_se), 
        .CLK(n1586), .Q(\mem0[248][2] ), .QN(n23614) );
  SDFFX1 \mem0_reg[248][1]  ( .D(n18541), .SI(\mem0[248][0] ), .SE(test_se), 
        .CLK(n1586), .Q(\mem0[248][1] ), .QN(n23615) );
  SDFFX1 \mem0_reg[248][0]  ( .D(n18540), .SI(\mem0[247][7] ), .SE(test_se), 
        .CLK(n1586), .Q(\mem0[248][0] ), .QN(n23616) );
  SDFFX1 \mem0_reg[247][7]  ( .D(n18539), .SI(\mem0[247][6] ), .SE(test_se), 
        .CLK(n1586), .Q(\mem0[247][7] ), .QN(n23617) );
  SDFFX1 \mem0_reg[247][6]  ( .D(n18538), .SI(\mem0[247][5] ), .SE(test_se), 
        .CLK(n1586), .Q(\mem0[247][6] ), .QN(n23618) );
  SDFFX1 \mem0_reg[247][5]  ( .D(n18537), .SI(\mem0[247][4] ), .SE(test_se), 
        .CLK(n1586), .Q(\mem0[247][5] ), .QN(n23619) );
  SDFFX1 \mem0_reg[247][4]  ( .D(n18536), .SI(\mem0[247][3] ), .SE(test_se), 
        .CLK(n1586), .Q(\mem0[247][4] ), .QN(n23620) );
  SDFFX1 \mem0_reg[247][3]  ( .D(n18535), .SI(\mem0[247][2] ), .SE(test_se), 
        .CLK(n1586), .Q(\mem0[247][3] ), .QN(n23621) );
  SDFFX1 \mem0_reg[247][2]  ( .D(n18534), .SI(\mem0[247][1] ), .SE(test_se), 
        .CLK(n1586), .Q(\mem0[247][2] ), .QN(n23622) );
  SDFFX1 \mem0_reg[247][1]  ( .D(n18533), .SI(\mem0[247][0] ), .SE(test_se), 
        .CLK(n1587), .Q(\mem0[247][1] ), .QN(n23623) );
  SDFFX1 \mem0_reg[247][0]  ( .D(n18532), .SI(\mem0[246][7] ), .SE(test_se), 
        .CLK(n1587), .Q(\mem0[247][0] ), .QN(n23624) );
  SDFFX1 \mem0_reg[246][7]  ( .D(n18531), .SI(\mem0[246][6] ), .SE(test_se), 
        .CLK(n1587), .Q(\mem0[246][7] ), .QN(n23625) );
  SDFFX1 \mem0_reg[246][6]  ( .D(n18530), .SI(\mem0[246][5] ), .SE(test_se), 
        .CLK(n1587), .Q(\mem0[246][6] ), .QN(n23626) );
  SDFFX1 \mem0_reg[246][5]  ( .D(n18529), .SI(\mem0[246][4] ), .SE(test_se), 
        .CLK(n1587), .Q(\mem0[246][5] ), .QN(n23627) );
  SDFFX1 \mem0_reg[246][4]  ( .D(n18528), .SI(\mem0[246][3] ), .SE(test_se), 
        .CLK(n1587), .Q(\mem0[246][4] ), .QN(n23628) );
  SDFFX1 \mem0_reg[246][3]  ( .D(n18527), .SI(\mem0[246][2] ), .SE(test_se), 
        .CLK(n1587), .Q(\mem0[246][3] ), .QN(n23629) );
  SDFFX1 \mem0_reg[246][2]  ( .D(n18526), .SI(\mem0[246][1] ), .SE(test_se), 
        .CLK(n1587), .Q(\mem0[246][2] ), .QN(n23630) );
  SDFFX1 \mem0_reg[246][1]  ( .D(n18525), .SI(\mem0[246][0] ), .SE(test_se), 
        .CLK(n1587), .Q(\mem0[246][1] ), .QN(n23631) );
  SDFFX1 \mem0_reg[246][0]  ( .D(n18524), .SI(\mem0[245][7] ), .SE(test_se), 
        .CLK(n1587), .Q(\mem0[246][0] ), .QN(n23632) );
  SDFFX1 \mem0_reg[245][7]  ( .D(n18523), .SI(\mem0[245][6] ), .SE(test_se), 
        .CLK(n1587), .Q(\mem0[245][7] ), .QN(n23633) );
  SDFFX1 \mem0_reg[245][6]  ( .D(n18522), .SI(\mem0[245][5] ), .SE(test_se), 
        .CLK(n1587), .Q(\mem0[245][6] ), .QN(n23634) );
  SDFFX1 \mem0_reg[245][5]  ( .D(n18521), .SI(\mem0[245][4] ), .SE(test_se), 
        .CLK(n1588), .Q(\mem0[245][5] ), .QN(n23635) );
  SDFFX1 \mem0_reg[245][4]  ( .D(n18520), .SI(\mem0[245][3] ), .SE(test_se), 
        .CLK(n1588), .Q(\mem0[245][4] ), .QN(n23636) );
  SDFFX1 \mem0_reg[245][3]  ( .D(n18519), .SI(\mem0[245][2] ), .SE(test_se), 
        .CLK(n1588), .Q(\mem0[245][3] ), .QN(n23637) );
  SDFFX1 \mem0_reg[245][2]  ( .D(n18518), .SI(\mem0[245][1] ), .SE(test_se), 
        .CLK(n1588), .Q(\mem0[245][2] ), .QN(n23638) );
  SDFFX1 \mem0_reg[245][1]  ( .D(n18517), .SI(\mem0[245][0] ), .SE(test_se), 
        .CLK(n1588), .Q(\mem0[245][1] ), .QN(n23639) );
  SDFFX1 \mem0_reg[245][0]  ( .D(n18516), .SI(\mem0[244][7] ), .SE(test_se), 
        .CLK(n1588), .Q(\mem0[245][0] ), .QN(n23640) );
  SDFFX1 \mem0_reg[244][7]  ( .D(n18515), .SI(\mem0[244][6] ), .SE(test_se), 
        .CLK(n1588), .Q(\mem0[244][7] ), .QN(n23641) );
  SDFFX1 \mem0_reg[244][6]  ( .D(n18514), .SI(\mem0[244][5] ), .SE(test_se), 
        .CLK(n1588), .Q(\mem0[244][6] ), .QN(n23642) );
  SDFFX1 \mem0_reg[244][5]  ( .D(n18513), .SI(\mem0[244][4] ), .SE(test_se), 
        .CLK(n1588), .Q(\mem0[244][5] ), .QN(n23643) );
  SDFFX1 \mem0_reg[244][4]  ( .D(n18512), .SI(\mem0[244][3] ), .SE(test_se), 
        .CLK(n1588), .Q(\mem0[244][4] ), .QN(n23644) );
  SDFFX1 \mem0_reg[244][3]  ( .D(n18511), .SI(\mem0[244][2] ), .SE(test_se), 
        .CLK(n1588), .Q(\mem0[244][3] ), .QN(n23645) );
  SDFFX1 \mem0_reg[244][2]  ( .D(n18510), .SI(\mem0[244][1] ), .SE(test_se), 
        .CLK(n1588), .Q(\mem0[244][2] ), .QN(n23646) );
  SDFFX1 \mem0_reg[244][1]  ( .D(n18509), .SI(\mem0[244][0] ), .SE(test_se), 
        .CLK(n1589), .Q(\mem0[244][1] ), .QN(n23647) );
  SDFFX1 \mem0_reg[244][0]  ( .D(n18508), .SI(\mem0[243][7] ), .SE(test_se), 
        .CLK(n1589), .Q(\mem0[244][0] ), .QN(n23648) );
  SDFFX1 \mem0_reg[243][7]  ( .D(n18507), .SI(\mem0[243][6] ), .SE(test_se), 
        .CLK(n1589), .Q(\mem0[243][7] ), .QN(n23649) );
  SDFFX1 \mem0_reg[243][6]  ( .D(n18506), .SI(\mem0[243][5] ), .SE(test_se), 
        .CLK(n1589), .Q(\mem0[243][6] ), .QN(n23650) );
  SDFFX1 \mem0_reg[243][5]  ( .D(n18505), .SI(\mem0[243][4] ), .SE(test_se), 
        .CLK(n1589), .Q(\mem0[243][5] ), .QN(n23651) );
  SDFFX1 \mem0_reg[243][4]  ( .D(n18504), .SI(\mem0[243][3] ), .SE(test_se), 
        .CLK(n1589), .Q(\mem0[243][4] ), .QN(n23652) );
  SDFFX1 \mem0_reg[243][3]  ( .D(n18503), .SI(\mem0[243][2] ), .SE(test_se), 
        .CLK(n1589), .Q(\mem0[243][3] ), .QN(n23653) );
  SDFFX1 \mem0_reg[243][2]  ( .D(n18502), .SI(\mem0[243][1] ), .SE(test_se), 
        .CLK(n1589), .Q(\mem0[243][2] ), .QN(n23654) );
  SDFFX1 \mem0_reg[243][1]  ( .D(n18501), .SI(\mem0[243][0] ), .SE(test_se), 
        .CLK(n1589), .Q(\mem0[243][1] ), .QN(n23655) );
  SDFFX1 \mem0_reg[243][0]  ( .D(n18500), .SI(\mem0[242][7] ), .SE(test_se), 
        .CLK(n1589), .Q(\mem0[243][0] ), .QN(n23656) );
  SDFFX1 \mem0_reg[242][7]  ( .D(n18499), .SI(\mem0[242][6] ), .SE(test_se), 
        .CLK(n1589), .Q(\mem0[242][7] ), .QN(n23657) );
  SDFFX1 \mem0_reg[242][6]  ( .D(n18498), .SI(\mem0[242][5] ), .SE(test_se), 
        .CLK(n1589), .Q(\mem0[242][6] ), .QN(n23658) );
  SDFFX1 \mem0_reg[242][5]  ( .D(n18497), .SI(\mem0[242][4] ), .SE(test_se), 
        .CLK(n1590), .Q(\mem0[242][5] ), .QN(n23659) );
  SDFFX1 \mem0_reg[242][4]  ( .D(n18496), .SI(\mem0[242][3] ), .SE(test_se), 
        .CLK(n1590), .Q(\mem0[242][4] ), .QN(n23660) );
  SDFFX1 \mem0_reg[242][3]  ( .D(n18495), .SI(\mem0[242][2] ), .SE(test_se), 
        .CLK(n1590), .Q(\mem0[242][3] ), .QN(n23661) );
  SDFFX1 \mem0_reg[242][2]  ( .D(n18494), .SI(\mem0[242][1] ), .SE(test_se), 
        .CLK(n1590), .Q(\mem0[242][2] ), .QN(n23662) );
  SDFFX1 \mem0_reg[242][1]  ( .D(n18493), .SI(\mem0[242][0] ), .SE(test_se), 
        .CLK(n1590), .Q(\mem0[242][1] ), .QN(n23663) );
  SDFFX1 \mem0_reg[242][0]  ( .D(n18492), .SI(\mem0[241][7] ), .SE(test_se), 
        .CLK(n1590), .Q(\mem0[242][0] ), .QN(n23664) );
  SDFFX1 \mem0_reg[241][7]  ( .D(n18491), .SI(\mem0[241][6] ), .SE(test_se), 
        .CLK(n1590), .Q(\mem0[241][7] ), .QN(n23665) );
  SDFFX1 \mem0_reg[241][6]  ( .D(n18490), .SI(\mem0[241][5] ), .SE(test_se), 
        .CLK(n1590), .Q(\mem0[241][6] ), .QN(n23666) );
  SDFFX1 \mem0_reg[241][5]  ( .D(n18489), .SI(\mem0[241][4] ), .SE(test_se), 
        .CLK(n1590), .Q(\mem0[241][5] ), .QN(n23667) );
  SDFFX1 \mem0_reg[241][4]  ( .D(n18488), .SI(\mem0[241][3] ), .SE(test_se), 
        .CLK(n1590), .Q(\mem0[241][4] ), .QN(n23668) );
  SDFFX1 \mem0_reg[241][3]  ( .D(n18487), .SI(\mem0[241][2] ), .SE(test_se), 
        .CLK(n1590), .Q(\mem0[241][3] ), .QN(n23669) );
  SDFFX1 \mem0_reg[241][2]  ( .D(n18486), .SI(\mem0[241][1] ), .SE(test_se), 
        .CLK(n1590), .Q(\mem0[241][2] ), .QN(n23670) );
  SDFFX1 \mem0_reg[241][1]  ( .D(n18485), .SI(\mem0[241][0] ), .SE(test_se), 
        .CLK(n1591), .Q(\mem0[241][1] ), .QN(n23671) );
  SDFFX1 \mem0_reg[241][0]  ( .D(n18484), .SI(\mem0[240][7] ), .SE(test_se), 
        .CLK(n1591), .Q(\mem0[241][0] ), .QN(n23672) );
  SDFFX1 \mem0_reg[240][7]  ( .D(n18483), .SI(\mem0[240][6] ), .SE(test_se), 
        .CLK(n1591), .Q(\mem0[240][7] ), .QN(n23673) );
  SDFFX1 \mem0_reg[240][6]  ( .D(n18482), .SI(\mem0[240][5] ), .SE(test_se), 
        .CLK(n1591), .Q(\mem0[240][6] ), .QN(n23674) );
  SDFFX1 \mem0_reg[240][5]  ( .D(n18481), .SI(\mem0[240][4] ), .SE(test_se), 
        .CLK(n1591), .Q(\mem0[240][5] ), .QN(n23675) );
  SDFFX1 \mem0_reg[240][4]  ( .D(n18480), .SI(\mem0[240][3] ), .SE(test_se), 
        .CLK(n1591), .Q(\mem0[240][4] ), .QN(n23676) );
  SDFFX1 \mem0_reg[240][3]  ( .D(n18479), .SI(\mem0[240][2] ), .SE(test_se), 
        .CLK(n1591), .Q(\mem0[240][3] ), .QN(n23677) );
  SDFFX1 \mem0_reg[240][2]  ( .D(n18478), .SI(\mem0[240][1] ), .SE(test_se), 
        .CLK(n1591), .Q(\mem0[240][2] ), .QN(n23678) );
  SDFFX1 \mem0_reg[240][1]  ( .D(n18477), .SI(\mem0[240][0] ), .SE(test_se), 
        .CLK(n1591), .Q(\mem0[240][1] ), .QN(n23679) );
  SDFFX1 \mem0_reg[240][0]  ( .D(n18476), .SI(\mem0[239][7] ), .SE(test_se), 
        .CLK(n1591), .Q(\mem0[240][0] ), .QN(n23680) );
  SDFFX1 \mem0_reg[239][7]  ( .D(n18475), .SI(\mem0[239][6] ), .SE(test_se), 
        .CLK(n1591), .Q(\mem0[239][7] ), .QN(n23681) );
  SDFFX1 \mem0_reg[239][6]  ( .D(n18474), .SI(\mem0[239][5] ), .SE(test_se), 
        .CLK(n1591), .Q(\mem0[239][6] ), .QN(n23682) );
  SDFFX1 \mem0_reg[239][5]  ( .D(n18473), .SI(\mem0[239][4] ), .SE(test_se), 
        .CLK(n1592), .Q(\mem0[239][5] ), .QN(n23683) );
  SDFFX1 \mem0_reg[239][4]  ( .D(n18472), .SI(\mem0[239][3] ), .SE(test_se), 
        .CLK(n1592), .Q(\mem0[239][4] ), .QN(n23684) );
  SDFFX1 \mem0_reg[239][3]  ( .D(n18471), .SI(\mem0[239][2] ), .SE(test_se), 
        .CLK(n1592), .Q(\mem0[239][3] ), .QN(n23685) );
  SDFFX1 \mem0_reg[239][2]  ( .D(n18470), .SI(\mem0[239][1] ), .SE(test_se), 
        .CLK(n1592), .Q(\mem0[239][2] ), .QN(n23686) );
  SDFFX1 \mem0_reg[239][1]  ( .D(n18469), .SI(\mem0[239][0] ), .SE(test_se), 
        .CLK(n1592), .Q(\mem0[239][1] ), .QN(n23687) );
  SDFFX1 \mem0_reg[239][0]  ( .D(n18468), .SI(\mem0[238][7] ), .SE(test_se), 
        .CLK(n1592), .Q(\mem0[239][0] ), .QN(n23688) );
  SDFFX1 \mem0_reg[238][7]  ( .D(n18467), .SI(\mem0[238][6] ), .SE(test_se), 
        .CLK(n1592), .Q(\mem0[238][7] ), .QN(n23689) );
  SDFFX1 \mem0_reg[238][6]  ( .D(n18466), .SI(\mem0[238][5] ), .SE(test_se), 
        .CLK(n1592), .Q(\mem0[238][6] ), .QN(n23690) );
  SDFFX1 \mem0_reg[238][5]  ( .D(n18465), .SI(\mem0[238][4] ), .SE(test_se), 
        .CLK(n1592), .Q(\mem0[238][5] ), .QN(n23691) );
  SDFFX1 \mem0_reg[238][4]  ( .D(n18464), .SI(\mem0[238][3] ), .SE(test_se), 
        .CLK(n1592), .Q(\mem0[238][4] ), .QN(n23692) );
  SDFFX1 \mem0_reg[238][3]  ( .D(n18463), .SI(\mem0[238][2] ), .SE(test_se), 
        .CLK(n1592), .Q(\mem0[238][3] ), .QN(n23693) );
  SDFFX1 \mem0_reg[238][2]  ( .D(n18462), .SI(\mem0[238][1] ), .SE(test_se), 
        .CLK(n1592), .Q(\mem0[238][2] ), .QN(n23694) );
  SDFFX1 \mem0_reg[238][1]  ( .D(n18461), .SI(\mem0[238][0] ), .SE(test_se), 
        .CLK(n1593), .Q(\mem0[238][1] ), .QN(n23695) );
  SDFFX1 \mem0_reg[238][0]  ( .D(n18460), .SI(\mem0[237][7] ), .SE(test_se), 
        .CLK(n1593), .Q(\mem0[238][0] ), .QN(n23696) );
  SDFFX1 \mem0_reg[237][7]  ( .D(n18459), .SI(\mem0[237][6] ), .SE(test_se), 
        .CLK(n1593), .Q(\mem0[237][7] ), .QN(n23697) );
  SDFFX1 \mem0_reg[237][6]  ( .D(n18458), .SI(\mem0[237][5] ), .SE(test_se), 
        .CLK(n1593), .Q(\mem0[237][6] ), .QN(n23698) );
  SDFFX1 \mem0_reg[237][5]  ( .D(n18457), .SI(\mem0[237][4] ), .SE(test_se), 
        .CLK(n1593), .Q(\mem0[237][5] ), .QN(n23699) );
  SDFFX1 \mem0_reg[237][4]  ( .D(n18456), .SI(\mem0[237][3] ), .SE(test_se), 
        .CLK(n1593), .Q(\mem0[237][4] ), .QN(n23700) );
  SDFFX1 \mem0_reg[237][3]  ( .D(n18455), .SI(\mem0[237][2] ), .SE(test_se), 
        .CLK(n1593), .Q(\mem0[237][3] ), .QN(n23701) );
  SDFFX1 \mem0_reg[237][2]  ( .D(n18454), .SI(\mem0[237][1] ), .SE(test_se), 
        .CLK(n1593), .Q(\mem0[237][2] ), .QN(n23702) );
  SDFFX1 \mem0_reg[237][1]  ( .D(n18453), .SI(\mem0[237][0] ), .SE(test_se), 
        .CLK(n1593), .Q(\mem0[237][1] ), .QN(n23703) );
  SDFFX1 \mem0_reg[237][0]  ( .D(n18452), .SI(\mem0[236][7] ), .SE(test_se), 
        .CLK(n1593), .Q(\mem0[237][0] ), .QN(n23704) );
  SDFFX1 \mem0_reg[236][7]  ( .D(n18451), .SI(\mem0[236][6] ), .SE(test_se), 
        .CLK(n1593), .Q(\mem0[236][7] ), .QN(n23705) );
  SDFFX1 \mem0_reg[236][6]  ( .D(n18450), .SI(\mem0[236][5] ), .SE(test_se), 
        .CLK(n1593), .Q(\mem0[236][6] ), .QN(n23706) );
  SDFFX1 \mem0_reg[236][5]  ( .D(n18449), .SI(\mem0[236][4] ), .SE(test_se), 
        .CLK(n1594), .Q(\mem0[236][5] ), .QN(n23707) );
  SDFFX1 \mem0_reg[236][4]  ( .D(n18448), .SI(\mem0[236][3] ), .SE(test_se), 
        .CLK(n1594), .Q(\mem0[236][4] ), .QN(n23708) );
  SDFFX1 \mem0_reg[236][3]  ( .D(n18447), .SI(\mem0[236][2] ), .SE(test_se), 
        .CLK(n1594), .Q(\mem0[236][3] ), .QN(n23709) );
  SDFFX1 \mem0_reg[236][2]  ( .D(n18446), .SI(\mem0[236][1] ), .SE(test_se), 
        .CLK(n1594), .Q(\mem0[236][2] ), .QN(n23710) );
  SDFFX1 \mem0_reg[236][1]  ( .D(n18445), .SI(\mem0[236][0] ), .SE(test_se), 
        .CLK(n1594), .Q(\mem0[236][1] ), .QN(n23711) );
  SDFFX1 \mem0_reg[236][0]  ( .D(n18444), .SI(\mem0[235][7] ), .SE(test_se), 
        .CLK(n1594), .Q(\mem0[236][0] ), .QN(n23712) );
  SDFFX1 \mem0_reg[235][7]  ( .D(n18443), .SI(\mem0[235][6] ), .SE(test_se), 
        .CLK(n1594), .Q(\mem0[235][7] ), .QN(n23713) );
  SDFFX1 \mem0_reg[235][6]  ( .D(n18442), .SI(\mem0[235][5] ), .SE(test_se), 
        .CLK(n1594), .Q(\mem0[235][6] ), .QN(n23714) );
  SDFFX1 \mem0_reg[235][5]  ( .D(n18441), .SI(\mem0[235][4] ), .SE(test_se), 
        .CLK(n1594), .Q(\mem0[235][5] ), .QN(n23715) );
  SDFFX1 \mem0_reg[235][4]  ( .D(n18440), .SI(\mem0[235][3] ), .SE(test_se), 
        .CLK(n1594), .Q(\mem0[235][4] ), .QN(n23716) );
  SDFFX1 \mem0_reg[235][3]  ( .D(n18439), .SI(\mem0[235][2] ), .SE(test_se), 
        .CLK(n1594), .Q(\mem0[235][3] ), .QN(n23717) );
  SDFFX1 \mem0_reg[235][2]  ( .D(n18438), .SI(\mem0[235][1] ), .SE(test_se), 
        .CLK(n1594), .Q(\mem0[235][2] ), .QN(n23718) );
  SDFFX1 \mem0_reg[235][1]  ( .D(n18437), .SI(\mem0[235][0] ), .SE(test_se), 
        .CLK(n1595), .Q(\mem0[235][1] ), .QN(n23719) );
  SDFFX1 \mem0_reg[235][0]  ( .D(n18436), .SI(\mem0[234][7] ), .SE(test_se), 
        .CLK(n1595), .Q(\mem0[235][0] ), .QN(n23720) );
  SDFFX1 \mem0_reg[234][7]  ( .D(n18435), .SI(\mem0[234][6] ), .SE(test_se), 
        .CLK(n1595), .Q(\mem0[234][7] ), .QN(n23721) );
  SDFFX1 \mem0_reg[234][6]  ( .D(n18434), .SI(\mem0[234][5] ), .SE(test_se), 
        .CLK(n1595), .Q(\mem0[234][6] ), .QN(n23722) );
  SDFFX1 \mem0_reg[234][5]  ( .D(n18433), .SI(\mem0[234][4] ), .SE(test_se), 
        .CLK(n1595), .Q(\mem0[234][5] ), .QN(n23723) );
  SDFFX1 \mem0_reg[234][4]  ( .D(n18432), .SI(\mem0[234][3] ), .SE(test_se), 
        .CLK(n1595), .Q(\mem0[234][4] ), .QN(n23724) );
  SDFFX1 \mem0_reg[234][3]  ( .D(n18431), .SI(\mem0[234][2] ), .SE(test_se), 
        .CLK(n1595), .Q(\mem0[234][3] ), .QN(n23725) );
  SDFFX1 \mem0_reg[234][2]  ( .D(n18430), .SI(\mem0[234][1] ), .SE(test_se), 
        .CLK(n1595), .Q(\mem0[234][2] ), .QN(n23726) );
  SDFFX1 \mem0_reg[234][1]  ( .D(n18429), .SI(\mem0[234][0] ), .SE(test_se), 
        .CLK(n1595), .Q(\mem0[234][1] ), .QN(n23727) );
  SDFFX1 \mem0_reg[234][0]  ( .D(n18428), .SI(\mem0[233][7] ), .SE(test_se), 
        .CLK(n1595), .Q(\mem0[234][0] ), .QN(n23728) );
  SDFFX1 \mem0_reg[233][7]  ( .D(n18427), .SI(\mem0[233][6] ), .SE(test_se), 
        .CLK(n1595), .Q(\mem0[233][7] ), .QN(n23729) );
  SDFFX1 \mem0_reg[233][6]  ( .D(n18426), .SI(\mem0[233][5] ), .SE(test_se), 
        .CLK(n1595), .Q(\mem0[233][6] ), .QN(n23730) );
  SDFFX1 \mem0_reg[233][5]  ( .D(n18425), .SI(\mem0[233][4] ), .SE(test_se), 
        .CLK(n1596), .Q(\mem0[233][5] ), .QN(n23731) );
  SDFFX1 \mem0_reg[233][4]  ( .D(n18424), .SI(\mem0[233][3] ), .SE(test_se), 
        .CLK(n1596), .Q(\mem0[233][4] ), .QN(n23732) );
  SDFFX1 \mem0_reg[233][3]  ( .D(n18423), .SI(\mem0[233][2] ), .SE(test_se), 
        .CLK(n1596), .Q(\mem0[233][3] ), .QN(n23733) );
  SDFFX1 \mem0_reg[233][2]  ( .D(n18422), .SI(\mem0[233][1] ), .SE(test_se), 
        .CLK(n1596), .Q(\mem0[233][2] ), .QN(n23734) );
  SDFFX1 \mem0_reg[233][1]  ( .D(n18421), .SI(\mem0[233][0] ), .SE(test_se), 
        .CLK(n1596), .Q(\mem0[233][1] ), .QN(n23735) );
  SDFFX1 \mem0_reg[233][0]  ( .D(n18420), .SI(\mem0[232][7] ), .SE(test_se), 
        .CLK(n1596), .Q(\mem0[233][0] ), .QN(n23736) );
  SDFFX1 \mem0_reg[232][7]  ( .D(n18419), .SI(\mem0[232][6] ), .SE(test_se), 
        .CLK(n1596), .Q(\mem0[232][7] ), .QN(n23737) );
  SDFFX1 \mem0_reg[232][6]  ( .D(n18418), .SI(\mem0[232][5] ), .SE(test_se), 
        .CLK(n1596), .Q(\mem0[232][6] ), .QN(n23738) );
  SDFFX1 \mem0_reg[232][5]  ( .D(n18417), .SI(\mem0[232][4] ), .SE(test_se), 
        .CLK(n1596), .Q(\mem0[232][5] ), .QN(n23739) );
  SDFFX1 \mem0_reg[232][4]  ( .D(n18416), .SI(\mem0[232][3] ), .SE(test_se), 
        .CLK(n1596), .Q(\mem0[232][4] ), .QN(n23740) );
  SDFFX1 \mem0_reg[232][3]  ( .D(n18415), .SI(\mem0[232][2] ), .SE(test_se), 
        .CLK(n1596), .Q(\mem0[232][3] ), .QN(n23741) );
  SDFFX1 \mem0_reg[232][2]  ( .D(n18414), .SI(\mem0[232][1] ), .SE(test_se), 
        .CLK(n1596), .Q(\mem0[232][2] ), .QN(n23742) );
  SDFFX1 \mem0_reg[232][1]  ( .D(n18413), .SI(\mem0[232][0] ), .SE(test_se), 
        .CLK(n1597), .Q(\mem0[232][1] ), .QN(n23743) );
  SDFFX1 \mem0_reg[232][0]  ( .D(n18412), .SI(\mem0[231][7] ), .SE(test_se), 
        .CLK(n1597), .Q(\mem0[232][0] ), .QN(n23744) );
  SDFFX1 \mem0_reg[231][7]  ( .D(n18411), .SI(\mem0[231][6] ), .SE(test_se), 
        .CLK(n1597), .Q(\mem0[231][7] ), .QN(n23745) );
  SDFFX1 \mem0_reg[231][6]  ( .D(n18410), .SI(\mem0[231][5] ), .SE(test_se), 
        .CLK(n1597), .Q(\mem0[231][6] ), .QN(n23746) );
  SDFFX1 \mem0_reg[231][5]  ( .D(n18409), .SI(\mem0[231][4] ), .SE(test_se), 
        .CLK(n1597), .Q(\mem0[231][5] ), .QN(n23747) );
  SDFFX1 \mem0_reg[231][4]  ( .D(n18408), .SI(\mem0[231][3] ), .SE(test_se), 
        .CLK(n1597), .Q(\mem0[231][4] ), .QN(n23748) );
  SDFFX1 \mem0_reg[231][3]  ( .D(n18407), .SI(\mem0[231][2] ), .SE(test_se), 
        .CLK(n1597), .Q(\mem0[231][3] ), .QN(n23749) );
  SDFFX1 \mem0_reg[231][2]  ( .D(n18406), .SI(\mem0[231][1] ), .SE(test_se), 
        .CLK(n1597), .Q(\mem0[231][2] ), .QN(n23750) );
  SDFFX1 \mem0_reg[231][1]  ( .D(n18405), .SI(\mem0[231][0] ), .SE(test_se), 
        .CLK(n1597), .Q(\mem0[231][1] ), .QN(n23751) );
  SDFFX1 \mem0_reg[231][0]  ( .D(n18404), .SI(\mem0[230][7] ), .SE(test_se), 
        .CLK(n1597), .Q(\mem0[231][0] ), .QN(n23752) );
  SDFFX1 \mem0_reg[230][7]  ( .D(n18403), .SI(\mem0[230][6] ), .SE(test_se), 
        .CLK(n1597), .Q(\mem0[230][7] ), .QN(n23753) );
  SDFFX1 \mem0_reg[230][6]  ( .D(n18402), .SI(\mem0[230][5] ), .SE(test_se), 
        .CLK(n1597), .Q(\mem0[230][6] ), .QN(n23754) );
  SDFFX1 \mem0_reg[230][5]  ( .D(n18401), .SI(\mem0[230][4] ), .SE(test_se), 
        .CLK(n1598), .Q(\mem0[230][5] ), .QN(n23755) );
  SDFFX1 \mem0_reg[230][4]  ( .D(n18400), .SI(\mem0[230][3] ), .SE(test_se), 
        .CLK(n1598), .Q(\mem0[230][4] ), .QN(n23756) );
  SDFFX1 \mem0_reg[230][3]  ( .D(n18399), .SI(\mem0[230][2] ), .SE(test_se), 
        .CLK(n1598), .Q(\mem0[230][3] ), .QN(n23757) );
  SDFFX1 \mem0_reg[230][2]  ( .D(n18398), .SI(\mem0[230][1] ), .SE(test_se), 
        .CLK(n1598), .Q(\mem0[230][2] ), .QN(n23758) );
  SDFFX1 \mem0_reg[230][1]  ( .D(n18397), .SI(\mem0[230][0] ), .SE(test_se), 
        .CLK(n1598), .Q(\mem0[230][1] ), .QN(n23759) );
  SDFFX1 \mem0_reg[230][0]  ( .D(n18396), .SI(\mem0[229][7] ), .SE(test_se), 
        .CLK(n1598), .Q(\mem0[230][0] ), .QN(n23760) );
  SDFFX1 \mem0_reg[229][7]  ( .D(n18395), .SI(\mem0[229][6] ), .SE(test_se), 
        .CLK(n1598), .Q(\mem0[229][7] ), .QN(n23761) );
  SDFFX1 \mem0_reg[229][6]  ( .D(n18394), .SI(\mem0[229][5] ), .SE(test_se), 
        .CLK(n1598), .Q(\mem0[229][6] ), .QN(n23762) );
  SDFFX1 \mem0_reg[229][5]  ( .D(n18393), .SI(\mem0[229][4] ), .SE(test_se), 
        .CLK(n1598), .Q(\mem0[229][5] ), .QN(n23763) );
  SDFFX1 \mem0_reg[229][4]  ( .D(n18392), .SI(\mem0[229][3] ), .SE(test_se), 
        .CLK(n1598), .Q(\mem0[229][4] ), .QN(n23764) );
  SDFFX1 \mem0_reg[229][3]  ( .D(n18391), .SI(\mem0[229][2] ), .SE(test_se), 
        .CLK(n1598), .Q(\mem0[229][3] ), .QN(n23765) );
  SDFFX1 \mem0_reg[229][2]  ( .D(n18390), .SI(\mem0[229][1] ), .SE(test_se), 
        .CLK(n1598), .Q(\mem0[229][2] ), .QN(n23766) );
  SDFFX1 \mem0_reg[229][1]  ( .D(n18389), .SI(\mem0[229][0] ), .SE(test_se), 
        .CLK(n1599), .Q(\mem0[229][1] ), .QN(n23767) );
  SDFFX1 \mem0_reg[229][0]  ( .D(n18388), .SI(\mem0[228][7] ), .SE(test_se), 
        .CLK(n1599), .Q(\mem0[229][0] ), .QN(n23768) );
  SDFFX1 \mem0_reg[228][7]  ( .D(n18387), .SI(\mem0[228][6] ), .SE(test_se), 
        .CLK(n1599), .Q(\mem0[228][7] ), .QN(n23769) );
  SDFFX1 \mem0_reg[228][6]  ( .D(n18386), .SI(\mem0[228][5] ), .SE(test_se), 
        .CLK(n1599), .Q(\mem0[228][6] ), .QN(n23770) );
  SDFFX1 \mem0_reg[228][5]  ( .D(n18385), .SI(\mem0[228][4] ), .SE(test_se), 
        .CLK(n1599), .Q(\mem0[228][5] ), .QN(n23771) );
  SDFFX1 \mem0_reg[228][4]  ( .D(n18384), .SI(\mem0[228][3] ), .SE(test_se), 
        .CLK(n1599), .Q(\mem0[228][4] ), .QN(n23772) );
  SDFFX1 \mem0_reg[228][3]  ( .D(n18383), .SI(\mem0[228][2] ), .SE(test_se), 
        .CLK(n1599), .Q(\mem0[228][3] ), .QN(n23773) );
  SDFFX1 \mem0_reg[228][2]  ( .D(n18382), .SI(\mem0[228][1] ), .SE(test_se), 
        .CLK(n1599), .Q(\mem0[228][2] ), .QN(n23774) );
  SDFFX1 \mem0_reg[228][1]  ( .D(n18381), .SI(\mem0[228][0] ), .SE(test_se), 
        .CLK(n1599), .Q(\mem0[228][1] ), .QN(n23775) );
  SDFFX1 \mem0_reg[228][0]  ( .D(n18380), .SI(\mem0[227][7] ), .SE(test_se), 
        .CLK(n1599), .Q(\mem0[228][0] ), .QN(n23776) );
  SDFFX1 \mem0_reg[227][7]  ( .D(n18379), .SI(\mem0[227][6] ), .SE(test_se), 
        .CLK(n1599), .Q(\mem0[227][7] ), .QN(n23777) );
  SDFFX1 \mem0_reg[227][6]  ( .D(n18378), .SI(\mem0[227][5] ), .SE(test_se), 
        .CLK(n1599), .Q(\mem0[227][6] ), .QN(n23778) );
  SDFFX1 \mem0_reg[227][5]  ( .D(n18377), .SI(\mem0[227][4] ), .SE(test_se), 
        .CLK(n1600), .Q(\mem0[227][5] ), .QN(n23779) );
  SDFFX1 \mem0_reg[227][4]  ( .D(n18376), .SI(\mem0[227][3] ), .SE(test_se), 
        .CLK(n1600), .Q(\mem0[227][4] ), .QN(n23780) );
  SDFFX1 \mem0_reg[227][3]  ( .D(n18375), .SI(\mem0[227][2] ), .SE(test_se), 
        .CLK(n1600), .Q(\mem0[227][3] ), .QN(n23781) );
  SDFFX1 \mem0_reg[227][2]  ( .D(n18374), .SI(\mem0[227][1] ), .SE(test_se), 
        .CLK(n1600), .Q(\mem0[227][2] ), .QN(n23782) );
  SDFFX1 \mem0_reg[227][1]  ( .D(n18373), .SI(\mem0[227][0] ), .SE(test_se), 
        .CLK(n1600), .Q(\mem0[227][1] ), .QN(n23783) );
  SDFFX1 \mem0_reg[227][0]  ( .D(n18372), .SI(\mem0[226][7] ), .SE(test_se), 
        .CLK(n1600), .Q(\mem0[227][0] ), .QN(n23784) );
  SDFFX1 \mem0_reg[226][7]  ( .D(n18371), .SI(\mem0[226][6] ), .SE(test_se), 
        .CLK(n1600), .Q(\mem0[226][7] ), .QN(n23785) );
  SDFFX1 \mem0_reg[226][6]  ( .D(n18370), .SI(\mem0[226][5] ), .SE(test_se), 
        .CLK(n1600), .Q(\mem0[226][6] ), .QN(n23786) );
  SDFFX1 \mem0_reg[226][5]  ( .D(n18369), .SI(\mem0[226][4] ), .SE(test_se), 
        .CLK(n1600), .Q(\mem0[226][5] ), .QN(n23787) );
  SDFFX1 \mem0_reg[226][4]  ( .D(n18368), .SI(\mem0[226][3] ), .SE(test_se), 
        .CLK(n1600), .Q(\mem0[226][4] ), .QN(n23788) );
  SDFFX1 \mem0_reg[226][3]  ( .D(n18367), .SI(\mem0[226][2] ), .SE(test_se), 
        .CLK(n1600), .Q(\mem0[226][3] ), .QN(n23789) );
  SDFFX1 \mem0_reg[226][2]  ( .D(n18366), .SI(\mem0[226][1] ), .SE(test_se), 
        .CLK(n1600), .Q(\mem0[226][2] ), .QN(n23790) );
  SDFFX1 \mem0_reg[226][1]  ( .D(n18365), .SI(\mem0[226][0] ), .SE(test_se), 
        .CLK(n1601), .Q(\mem0[226][1] ), .QN(n23791) );
  SDFFX1 \mem0_reg[226][0]  ( .D(n18364), .SI(\mem0[225][7] ), .SE(test_se), 
        .CLK(n1601), .Q(\mem0[226][0] ), .QN(n23792) );
  SDFFX1 \mem0_reg[225][7]  ( .D(n18363), .SI(\mem0[225][6] ), .SE(test_se), 
        .CLK(n1601), .Q(\mem0[225][7] ), .QN(n23793) );
  SDFFX1 \mem0_reg[225][6]  ( .D(n18362), .SI(\mem0[225][5] ), .SE(test_se), 
        .CLK(n1601), .Q(\mem0[225][6] ), .QN(n23794) );
  SDFFX1 \mem0_reg[225][5]  ( .D(n18361), .SI(\mem0[225][4] ), .SE(test_se), 
        .CLK(n1601), .Q(\mem0[225][5] ), .QN(n23795) );
  SDFFX1 \mem0_reg[225][4]  ( .D(n18360), .SI(\mem0[225][3] ), .SE(test_se), 
        .CLK(n1601), .Q(\mem0[225][4] ), .QN(n23796) );
  SDFFX1 \mem0_reg[225][3]  ( .D(n18359), .SI(\mem0[225][2] ), .SE(test_se), 
        .CLK(n1601), .Q(\mem0[225][3] ), .QN(n23797) );
  SDFFX1 \mem0_reg[225][2]  ( .D(n18358), .SI(\mem0[225][1] ), .SE(test_se), 
        .CLK(n1601), .Q(\mem0[225][2] ), .QN(n23798) );
  SDFFX1 \mem0_reg[225][1]  ( .D(n18357), .SI(\mem0[225][0] ), .SE(test_se), 
        .CLK(n1601), .Q(\mem0[225][1] ), .QN(n23799) );
  SDFFX1 \mem0_reg[225][0]  ( .D(n18356), .SI(\mem0[224][7] ), .SE(test_se), 
        .CLK(n1601), .Q(\mem0[225][0] ), .QN(n23800) );
  SDFFX1 \mem0_reg[224][7]  ( .D(n18355), .SI(\mem0[224][6] ), .SE(test_se), 
        .CLK(n1601), .Q(\mem0[224][7] ), .QN(n23801) );
  SDFFX1 \mem0_reg[224][6]  ( .D(n18354), .SI(\mem0[224][5] ), .SE(test_se), 
        .CLK(n1601), .Q(\mem0[224][6] ), .QN(n23802) );
  SDFFX1 \mem0_reg[224][5]  ( .D(n18353), .SI(\mem0[224][4] ), .SE(test_se), 
        .CLK(n1602), .Q(\mem0[224][5] ), .QN(n23803) );
  SDFFX1 \mem0_reg[224][4]  ( .D(n18352), .SI(\mem0[224][3] ), .SE(test_se), 
        .CLK(n1602), .Q(\mem0[224][4] ), .QN(n23804) );
  SDFFX1 \mem0_reg[224][3]  ( .D(n18351), .SI(\mem0[224][2] ), .SE(test_se), 
        .CLK(n1602), .Q(\mem0[224][3] ), .QN(n23805) );
  SDFFX1 \mem0_reg[224][2]  ( .D(n18350), .SI(\mem0[224][1] ), .SE(test_se), 
        .CLK(n1602), .Q(\mem0[224][2] ), .QN(n23806) );
  SDFFX1 \mem0_reg[224][1]  ( .D(n18349), .SI(\mem0[224][0] ), .SE(test_se), 
        .CLK(n1602), .Q(\mem0[224][1] ), .QN(n23807) );
  SDFFX1 \mem0_reg[224][0]  ( .D(n18348), .SI(\mem0[223][7] ), .SE(test_se), 
        .CLK(n1602), .Q(\mem0[224][0] ), .QN(n23808) );
  SDFFX1 \mem0_reg[223][7]  ( .D(n18347), .SI(\mem0[223][6] ), .SE(test_se), 
        .CLK(n1602), .Q(\mem0[223][7] ), .QN(n23809) );
  SDFFX1 \mem0_reg[223][6]  ( .D(n18346), .SI(\mem0[223][5] ), .SE(test_se), 
        .CLK(n1602), .Q(\mem0[223][6] ), .QN(n23810) );
  SDFFX1 \mem0_reg[223][5]  ( .D(n18345), .SI(\mem0[223][4] ), .SE(test_se), 
        .CLK(n1602), .Q(\mem0[223][5] ), .QN(n23811) );
  SDFFX1 \mem0_reg[223][4]  ( .D(n18344), .SI(\mem0[223][3] ), .SE(test_se), 
        .CLK(n1602), .Q(\mem0[223][4] ), .QN(n23812) );
  SDFFX1 \mem0_reg[223][3]  ( .D(n18343), .SI(\mem0[223][2] ), .SE(test_se), 
        .CLK(n1602), .Q(\mem0[223][3] ), .QN(n23813) );
  SDFFX1 \mem0_reg[223][2]  ( .D(n18342), .SI(\mem0[223][1] ), .SE(test_se), 
        .CLK(n1602), .Q(\mem0[223][2] ), .QN(n23814) );
  SDFFX1 \mem0_reg[223][1]  ( .D(n18341), .SI(\mem0[223][0] ), .SE(test_se), 
        .CLK(n1603), .Q(\mem0[223][1] ), .QN(n23815) );
  SDFFX1 \mem0_reg[223][0]  ( .D(n18340), .SI(\mem0[222][7] ), .SE(test_se), 
        .CLK(n1603), .Q(\mem0[223][0] ), .QN(n23816) );
  SDFFX1 \mem0_reg[222][7]  ( .D(n18339), .SI(\mem0[222][6] ), .SE(test_se), 
        .CLK(n1603), .Q(\mem0[222][7] ), .QN(n23817) );
  SDFFX1 \mem0_reg[222][6]  ( .D(n18338), .SI(\mem0[222][5] ), .SE(test_se), 
        .CLK(n1603), .Q(\mem0[222][6] ), .QN(n23818) );
  SDFFX1 \mem0_reg[222][5]  ( .D(n18337), .SI(\mem0[222][4] ), .SE(test_se), 
        .CLK(n1603), .Q(\mem0[222][5] ), .QN(n23819) );
  SDFFX1 \mem0_reg[222][4]  ( .D(n18336), .SI(\mem0[222][3] ), .SE(test_se), 
        .CLK(n1603), .Q(\mem0[222][4] ), .QN(n23820) );
  SDFFX1 \mem0_reg[222][3]  ( .D(n18335), .SI(\mem0[222][2] ), .SE(test_se), 
        .CLK(n1603), .Q(\mem0[222][3] ), .QN(n23821) );
  SDFFX1 \mem0_reg[222][2]  ( .D(n18334), .SI(\mem0[222][1] ), .SE(test_se), 
        .CLK(n1603), .Q(\mem0[222][2] ), .QN(n23822) );
  SDFFX1 \mem0_reg[222][1]  ( .D(n18333), .SI(\mem0[222][0] ), .SE(test_se), 
        .CLK(n1603), .Q(\mem0[222][1] ), .QN(n23823) );
  SDFFX1 \mem0_reg[222][0]  ( .D(n18332), .SI(\mem0[221][7] ), .SE(test_se), 
        .CLK(n1603), .Q(\mem0[222][0] ), .QN(n23824) );
  SDFFX1 \mem0_reg[221][7]  ( .D(n18331), .SI(\mem0[221][6] ), .SE(test_se), 
        .CLK(n1603), .Q(\mem0[221][7] ), .QN(n23825) );
  SDFFX1 \mem0_reg[221][6]  ( .D(n18330), .SI(\mem0[221][5] ), .SE(test_se), 
        .CLK(n1603), .Q(\mem0[221][6] ), .QN(n23826) );
  SDFFX1 \mem0_reg[221][5]  ( .D(n18329), .SI(\mem0[221][4] ), .SE(test_se), 
        .CLK(n1604), .Q(\mem0[221][5] ), .QN(n23827) );
  SDFFX1 \mem0_reg[221][4]  ( .D(n18328), .SI(\mem0[221][3] ), .SE(test_se), 
        .CLK(n1604), .Q(\mem0[221][4] ), .QN(n23828) );
  SDFFX1 \mem0_reg[221][3]  ( .D(n18327), .SI(\mem0[221][2] ), .SE(test_se), 
        .CLK(n1604), .Q(\mem0[221][3] ), .QN(n23829) );
  SDFFX1 \mem0_reg[221][2]  ( .D(n18326), .SI(\mem0[221][1] ), .SE(test_se), 
        .CLK(n1604), .Q(\mem0[221][2] ), .QN(n23830) );
  SDFFX1 \mem0_reg[221][1]  ( .D(n18325), .SI(\mem0[221][0] ), .SE(test_se), 
        .CLK(n1604), .Q(\mem0[221][1] ), .QN(n23831) );
  SDFFX1 \mem0_reg[221][0]  ( .D(n18324), .SI(\mem0[220][7] ), .SE(test_se), 
        .CLK(n1604), .Q(\mem0[221][0] ), .QN(n23832) );
  SDFFX1 \mem0_reg[220][7]  ( .D(n18323), .SI(\mem0[220][6] ), .SE(test_se), 
        .CLK(n1604), .Q(\mem0[220][7] ), .QN(n23833) );
  SDFFX1 \mem0_reg[220][6]  ( .D(n18322), .SI(\mem0[220][5] ), .SE(test_se), 
        .CLK(n1604), .Q(\mem0[220][6] ), .QN(n23834) );
  SDFFX1 \mem0_reg[220][5]  ( .D(n18321), .SI(\mem0[220][4] ), .SE(test_se), 
        .CLK(n1604), .Q(\mem0[220][5] ), .QN(n23835) );
  SDFFX1 \mem0_reg[220][4]  ( .D(n18320), .SI(\mem0[220][3] ), .SE(test_se), 
        .CLK(n1604), .Q(\mem0[220][4] ), .QN(n23836) );
  SDFFX1 \mem0_reg[220][3]  ( .D(n18319), .SI(\mem0[220][2] ), .SE(test_se), 
        .CLK(n1604), .Q(\mem0[220][3] ), .QN(n23837) );
  SDFFX1 \mem0_reg[220][2]  ( .D(n18318), .SI(\mem0[220][1] ), .SE(test_se), 
        .CLK(n1604), .Q(\mem0[220][2] ), .QN(n23838) );
  SDFFX1 \mem0_reg[220][1]  ( .D(n18317), .SI(\mem0[220][0] ), .SE(test_se), 
        .CLK(n1605), .Q(\mem0[220][1] ), .QN(n23839) );
  SDFFX1 \mem0_reg[220][0]  ( .D(n18316), .SI(\mem0[219][7] ), .SE(test_se), 
        .CLK(n1605), .Q(\mem0[220][0] ), .QN(n23840) );
  SDFFX1 \mem0_reg[219][7]  ( .D(n18315), .SI(\mem0[219][6] ), .SE(test_se), 
        .CLK(n1605), .Q(\mem0[219][7] ), .QN(n23841) );
  SDFFX1 \mem0_reg[219][6]  ( .D(n18314), .SI(\mem0[219][5] ), .SE(test_se), 
        .CLK(n1605), .Q(\mem0[219][6] ), .QN(n23842) );
  SDFFX1 \mem0_reg[219][5]  ( .D(n18313), .SI(\mem0[219][4] ), .SE(test_se), 
        .CLK(n1605), .Q(\mem0[219][5] ), .QN(n23843) );
  SDFFX1 \mem0_reg[219][4]  ( .D(n18312), .SI(\mem0[219][3] ), .SE(test_se), 
        .CLK(n1605), .Q(\mem0[219][4] ), .QN(n23844) );
  SDFFX1 \mem0_reg[219][3]  ( .D(n18311), .SI(\mem0[219][2] ), .SE(test_se), 
        .CLK(n1605), .Q(\mem0[219][3] ), .QN(n23845) );
  SDFFX1 \mem0_reg[219][2]  ( .D(n18310), .SI(\mem0[219][1] ), .SE(test_se), 
        .CLK(n1605), .Q(\mem0[219][2] ), .QN(n23846) );
  SDFFX1 \mem0_reg[219][1]  ( .D(n18309), .SI(\mem0[219][0] ), .SE(test_se), 
        .CLK(n1605), .Q(\mem0[219][1] ), .QN(n23847) );
  SDFFX1 \mem0_reg[219][0]  ( .D(n18308), .SI(\mem0[218][7] ), .SE(test_se), 
        .CLK(n1605), .Q(\mem0[219][0] ), .QN(n23848) );
  SDFFX1 \mem0_reg[218][7]  ( .D(n18307), .SI(\mem0[218][6] ), .SE(test_se), 
        .CLK(n1605), .Q(\mem0[218][7] ), .QN(n23849) );
  SDFFX1 \mem0_reg[218][6]  ( .D(n18306), .SI(\mem0[218][5] ), .SE(test_se), 
        .CLK(n1605), .Q(\mem0[218][6] ), .QN(n23850) );
  SDFFX1 \mem0_reg[218][5]  ( .D(n18305), .SI(\mem0[218][4] ), .SE(test_se), 
        .CLK(n1606), .Q(\mem0[218][5] ), .QN(n23851) );
  SDFFX1 \mem0_reg[218][4]  ( .D(n18304), .SI(\mem0[218][3] ), .SE(test_se), 
        .CLK(n1606), .Q(\mem0[218][4] ), .QN(n23852) );
  SDFFX1 \mem0_reg[218][3]  ( .D(n18303), .SI(\mem0[218][2] ), .SE(test_se), 
        .CLK(n1606), .Q(\mem0[218][3] ), .QN(n23853) );
  SDFFX1 \mem0_reg[218][2]  ( .D(n18302), .SI(\mem0[218][1] ), .SE(test_se), 
        .CLK(n1606), .Q(\mem0[218][2] ), .QN(n23854) );
  SDFFX1 \mem0_reg[218][1]  ( .D(n18301), .SI(\mem0[218][0] ), .SE(test_se), 
        .CLK(n1606), .Q(\mem0[218][1] ), .QN(n23855) );
  SDFFX1 \mem0_reg[218][0]  ( .D(n18300), .SI(\mem0[217][7] ), .SE(test_se), 
        .CLK(n1606), .Q(\mem0[218][0] ), .QN(n23856) );
  SDFFX1 \mem0_reg[217][7]  ( .D(n18299), .SI(\mem0[217][6] ), .SE(test_se), 
        .CLK(n1606), .Q(\mem0[217][7] ), .QN(n23857) );
  SDFFX1 \mem0_reg[217][6]  ( .D(n18298), .SI(\mem0[217][5] ), .SE(test_se), 
        .CLK(n1606), .Q(\mem0[217][6] ), .QN(n23858) );
  SDFFX1 \mem0_reg[217][5]  ( .D(n18297), .SI(\mem0[217][4] ), .SE(test_se), 
        .CLK(n1606), .Q(\mem0[217][5] ), .QN(n23859) );
  SDFFX1 \mem0_reg[217][4]  ( .D(n18296), .SI(\mem0[217][3] ), .SE(test_se), 
        .CLK(n1606), .Q(\mem0[217][4] ), .QN(n23860) );
  SDFFX1 \mem0_reg[217][3]  ( .D(n18295), .SI(\mem0[217][2] ), .SE(test_se), 
        .CLK(n1606), .Q(\mem0[217][3] ), .QN(n23861) );
  SDFFX1 \mem0_reg[217][2]  ( .D(n18294), .SI(\mem0[217][1] ), .SE(test_se), 
        .CLK(n1606), .Q(\mem0[217][2] ), .QN(n23862) );
  SDFFX1 \mem0_reg[217][1]  ( .D(n18293), .SI(\mem0[217][0] ), .SE(test_se), 
        .CLK(n1607), .Q(\mem0[217][1] ), .QN(n23863) );
  SDFFX1 \mem0_reg[217][0]  ( .D(n18292), .SI(\mem0[216][7] ), .SE(test_se), 
        .CLK(n1607), .Q(\mem0[217][0] ), .QN(n23864) );
  SDFFX1 \mem0_reg[216][7]  ( .D(n18291), .SI(\mem0[216][6] ), .SE(test_se), 
        .CLK(n1607), .Q(\mem0[216][7] ), .QN(n23865) );
  SDFFX1 \mem0_reg[216][6]  ( .D(n18290), .SI(\mem0[216][5] ), .SE(test_se), 
        .CLK(n1607), .Q(\mem0[216][6] ), .QN(n23866) );
  SDFFX1 \mem0_reg[216][5]  ( .D(n18289), .SI(\mem0[216][4] ), .SE(test_se), 
        .CLK(n1607), .Q(\mem0[216][5] ), .QN(n23867) );
  SDFFX1 \mem0_reg[216][4]  ( .D(n18288), .SI(\mem0[216][3] ), .SE(test_se), 
        .CLK(n1607), .Q(\mem0[216][4] ), .QN(n23868) );
  SDFFX1 \mem0_reg[216][3]  ( .D(n18287), .SI(\mem0[216][2] ), .SE(test_se), 
        .CLK(n1607), .Q(\mem0[216][3] ), .QN(n23869) );
  SDFFX1 \mem0_reg[216][2]  ( .D(n18286), .SI(\mem0[216][1] ), .SE(test_se), 
        .CLK(n1607), .Q(\mem0[216][2] ), .QN(n23870) );
  SDFFX1 \mem0_reg[216][1]  ( .D(n18285), .SI(\mem0[216][0] ), .SE(test_se), 
        .CLK(n1607), .Q(\mem0[216][1] ), .QN(n23871) );
  SDFFX1 \mem0_reg[216][0]  ( .D(n18284), .SI(\mem0[215][7] ), .SE(test_se), 
        .CLK(n1607), .Q(\mem0[216][0] ), .QN(n23872) );
  SDFFX1 \mem0_reg[215][7]  ( .D(n18283), .SI(\mem0[215][6] ), .SE(test_se), 
        .CLK(n1607), .Q(\mem0[215][7] ), .QN(n23873) );
  SDFFX1 \mem0_reg[215][6]  ( .D(n18282), .SI(\mem0[215][5] ), .SE(test_se), 
        .CLK(n1607), .Q(\mem0[215][6] ), .QN(n23874) );
  SDFFX1 \mem0_reg[215][5]  ( .D(n18281), .SI(\mem0[215][4] ), .SE(test_se), 
        .CLK(n1608), .Q(\mem0[215][5] ), .QN(n23875) );
  SDFFX1 \mem0_reg[215][4]  ( .D(n18280), .SI(\mem0[215][3] ), .SE(test_se), 
        .CLK(n1608), .Q(\mem0[215][4] ), .QN(n23876) );
  SDFFX1 \mem0_reg[215][3]  ( .D(n18279), .SI(\mem0[215][2] ), .SE(test_se), 
        .CLK(n1608), .Q(\mem0[215][3] ), .QN(n23877) );
  SDFFX1 \mem0_reg[215][2]  ( .D(n18278), .SI(\mem0[215][1] ), .SE(test_se), 
        .CLK(n1608), .Q(\mem0[215][2] ), .QN(n23878) );
  SDFFX1 \mem0_reg[215][1]  ( .D(n18277), .SI(\mem0[215][0] ), .SE(test_se), 
        .CLK(n1608), .Q(\mem0[215][1] ), .QN(n23879) );
  SDFFX1 \mem0_reg[215][0]  ( .D(n18276), .SI(\mem0[214][7] ), .SE(test_se), 
        .CLK(n1608), .Q(\mem0[215][0] ), .QN(n23880) );
  SDFFX1 \mem0_reg[214][7]  ( .D(n18275), .SI(\mem0[214][6] ), .SE(test_se), 
        .CLK(n1608), .Q(\mem0[214][7] ), .QN(n23881) );
  SDFFX1 \mem0_reg[214][6]  ( .D(n18274), .SI(\mem0[214][5] ), .SE(test_se), 
        .CLK(n1608), .Q(\mem0[214][6] ), .QN(n23882) );
  SDFFX1 \mem0_reg[214][5]  ( .D(n18273), .SI(\mem0[214][4] ), .SE(test_se), 
        .CLK(n1608), .Q(\mem0[214][5] ), .QN(n23883) );
  SDFFX1 \mem0_reg[214][4]  ( .D(n18272), .SI(\mem0[214][3] ), .SE(test_se), 
        .CLK(n1608), .Q(\mem0[214][4] ), .QN(n23884) );
  SDFFX1 \mem0_reg[214][3]  ( .D(n18271), .SI(\mem0[214][2] ), .SE(test_se), 
        .CLK(n1608), .Q(\mem0[214][3] ), .QN(n23885) );
  SDFFX1 \mem0_reg[214][2]  ( .D(n18270), .SI(\mem0[214][1] ), .SE(test_se), 
        .CLK(n1608), .Q(\mem0[214][2] ), .QN(n23886) );
  SDFFX1 \mem0_reg[214][1]  ( .D(n18269), .SI(\mem0[214][0] ), .SE(test_se), 
        .CLK(n1609), .Q(\mem0[214][1] ), .QN(n23887) );
  SDFFX1 \mem0_reg[214][0]  ( .D(n18268), .SI(\mem0[213][7] ), .SE(test_se), 
        .CLK(n1609), .Q(\mem0[214][0] ), .QN(n23888) );
  SDFFX1 \mem0_reg[213][7]  ( .D(n18267), .SI(\mem0[213][6] ), .SE(test_se), 
        .CLK(n1609), .Q(\mem0[213][7] ), .QN(n23889) );
  SDFFX1 \mem0_reg[213][6]  ( .D(n18266), .SI(\mem0[213][5] ), .SE(test_se), 
        .CLK(n1609), .Q(\mem0[213][6] ), .QN(n23890) );
  SDFFX1 \mem0_reg[213][5]  ( .D(n18265), .SI(\mem0[213][4] ), .SE(test_se), 
        .CLK(n1609), .Q(\mem0[213][5] ), .QN(n23891) );
  SDFFX1 \mem0_reg[213][4]  ( .D(n18264), .SI(\mem0[213][3] ), .SE(test_se), 
        .CLK(n1609), .Q(\mem0[213][4] ), .QN(n23892) );
  SDFFX1 \mem0_reg[213][3]  ( .D(n18263), .SI(\mem0[213][2] ), .SE(test_se), 
        .CLK(n1609), .Q(\mem0[213][3] ), .QN(n23893) );
  SDFFX1 \mem0_reg[213][2]  ( .D(n18262), .SI(\mem0[213][1] ), .SE(test_se), 
        .CLK(n1609), .Q(\mem0[213][2] ), .QN(n23894) );
  SDFFX1 \mem0_reg[213][1]  ( .D(n18261), .SI(\mem0[213][0] ), .SE(test_se), 
        .CLK(n1609), .Q(\mem0[213][1] ), .QN(n23895) );
  SDFFX1 \mem0_reg[213][0]  ( .D(n18260), .SI(\mem0[212][7] ), .SE(test_se), 
        .CLK(n1609), .Q(\mem0[213][0] ), .QN(n23896) );
  SDFFX1 \mem0_reg[212][7]  ( .D(n18259), .SI(\mem0[212][6] ), .SE(test_se), 
        .CLK(n1609), .Q(\mem0[212][7] ), .QN(n23897) );
  SDFFX1 \mem0_reg[212][6]  ( .D(n18258), .SI(\mem0[212][5] ), .SE(test_se), 
        .CLK(n1609), .Q(\mem0[212][6] ), .QN(n23898) );
  SDFFX1 \mem0_reg[212][5]  ( .D(n18257), .SI(\mem0[212][4] ), .SE(test_se), 
        .CLK(n1610), .Q(\mem0[212][5] ), .QN(n23899) );
  SDFFX1 \mem0_reg[212][4]  ( .D(n18256), .SI(\mem0[212][3] ), .SE(test_se), 
        .CLK(n1610), .Q(\mem0[212][4] ), .QN(n23900) );
  SDFFX1 \mem0_reg[212][3]  ( .D(n18255), .SI(\mem0[212][2] ), .SE(test_se), 
        .CLK(n1610), .Q(\mem0[212][3] ), .QN(n23901) );
  SDFFX1 \mem0_reg[212][2]  ( .D(n18254), .SI(\mem0[212][1] ), .SE(test_se), 
        .CLK(n1610), .Q(\mem0[212][2] ), .QN(n23902) );
  SDFFX1 \mem0_reg[212][1]  ( .D(n18253), .SI(\mem0[212][0] ), .SE(test_se), 
        .CLK(n1610), .Q(\mem0[212][1] ), .QN(n23903) );
  SDFFX1 \mem0_reg[212][0]  ( .D(n18252), .SI(\mem0[211][7] ), .SE(test_se), 
        .CLK(n1610), .Q(\mem0[212][0] ), .QN(n23904) );
  SDFFX1 \mem0_reg[211][7]  ( .D(n18251), .SI(\mem0[211][6] ), .SE(test_se), 
        .CLK(n1610), .Q(\mem0[211][7] ), .QN(n23905) );
  SDFFX1 \mem0_reg[211][6]  ( .D(n18250), .SI(\mem0[211][5] ), .SE(test_se), 
        .CLK(n1610), .Q(\mem0[211][6] ), .QN(n23906) );
  SDFFX1 \mem0_reg[211][5]  ( .D(n18249), .SI(\mem0[211][4] ), .SE(test_se), 
        .CLK(n1610), .Q(\mem0[211][5] ), .QN(n23907) );
  SDFFX1 \mem0_reg[211][4]  ( .D(n18248), .SI(\mem0[211][3] ), .SE(test_se), 
        .CLK(n1610), .Q(\mem0[211][4] ), .QN(n23908) );
  SDFFX1 \mem0_reg[211][3]  ( .D(n18247), .SI(\mem0[211][2] ), .SE(test_se), 
        .CLK(n1610), .Q(\mem0[211][3] ), .QN(n23909) );
  SDFFX1 \mem0_reg[211][2]  ( .D(n18246), .SI(\mem0[211][1] ), .SE(test_se), 
        .CLK(n1610), .Q(\mem0[211][2] ), .QN(n23910) );
  SDFFX1 \mem0_reg[211][1]  ( .D(n18245), .SI(\mem0[211][0] ), .SE(test_se), 
        .CLK(n1611), .Q(\mem0[211][1] ), .QN(n23911) );
  SDFFX1 \mem0_reg[211][0]  ( .D(n18244), .SI(\mem0[210][7] ), .SE(test_se), 
        .CLK(n1611), .Q(\mem0[211][0] ), .QN(n23912) );
  SDFFX1 \mem0_reg[210][7]  ( .D(n18243), .SI(\mem0[210][6] ), .SE(test_se), 
        .CLK(n1611), .Q(\mem0[210][7] ), .QN(n23913) );
  SDFFX1 \mem0_reg[210][6]  ( .D(n18242), .SI(\mem0[210][5] ), .SE(test_se), 
        .CLK(n1611), .Q(\mem0[210][6] ), .QN(n23914) );
  SDFFX1 \mem0_reg[210][5]  ( .D(n18241), .SI(\mem0[210][4] ), .SE(test_se), 
        .CLK(n1611), .Q(\mem0[210][5] ), .QN(n23915) );
  SDFFX1 \mem0_reg[210][4]  ( .D(n18240), .SI(\mem0[210][3] ), .SE(test_se), 
        .CLK(n1611), .Q(\mem0[210][4] ), .QN(n23916) );
  SDFFX1 \mem0_reg[210][3]  ( .D(n18239), .SI(\mem0[210][2] ), .SE(test_se), 
        .CLK(n1611), .Q(\mem0[210][3] ), .QN(n23917) );
  SDFFX1 \mem0_reg[210][2]  ( .D(n18238), .SI(\mem0[210][1] ), .SE(test_se), 
        .CLK(n1611), .Q(\mem0[210][2] ), .QN(n23918) );
  SDFFX1 \mem0_reg[210][1]  ( .D(n18237), .SI(\mem0[210][0] ), .SE(test_se), 
        .CLK(n1611), .Q(\mem0[210][1] ), .QN(n23919) );
  SDFFX1 \mem0_reg[210][0]  ( .D(n18236), .SI(\mem0[209][7] ), .SE(test_se), 
        .CLK(n1611), .Q(\mem0[210][0] ), .QN(n23920) );
  SDFFX1 \mem0_reg[209][7]  ( .D(n18235), .SI(\mem0[209][6] ), .SE(test_se), 
        .CLK(n1611), .Q(\mem0[209][7] ), .QN(n23921) );
  SDFFX1 \mem0_reg[209][6]  ( .D(n18234), .SI(\mem0[209][5] ), .SE(test_se), 
        .CLK(n1611), .Q(\mem0[209][6] ), .QN(n23922) );
  SDFFX1 \mem0_reg[209][5]  ( .D(n18233), .SI(\mem0[209][4] ), .SE(test_se), 
        .CLK(n1612), .Q(\mem0[209][5] ), .QN(n23923) );
  SDFFX1 \mem0_reg[209][4]  ( .D(n18232), .SI(\mem0[209][3] ), .SE(test_se), 
        .CLK(n1612), .Q(\mem0[209][4] ), .QN(n23924) );
  SDFFX1 \mem0_reg[209][3]  ( .D(n18231), .SI(\mem0[209][2] ), .SE(test_se), 
        .CLK(n1612), .Q(\mem0[209][3] ), .QN(n23925) );
  SDFFX1 \mem0_reg[209][2]  ( .D(n18230), .SI(\mem0[209][1] ), .SE(test_se), 
        .CLK(n1612), .Q(\mem0[209][2] ), .QN(n23926) );
  SDFFX1 \mem0_reg[209][1]  ( .D(n18229), .SI(\mem0[209][0] ), .SE(test_se), 
        .CLK(n1612), .Q(\mem0[209][1] ), .QN(n23927) );
  SDFFX1 \mem0_reg[209][0]  ( .D(n18228), .SI(\mem0[208][7] ), .SE(test_se), 
        .CLK(n1612), .Q(\mem0[209][0] ), .QN(n23928) );
  SDFFX1 \mem0_reg[208][7]  ( .D(n18227), .SI(\mem0[208][6] ), .SE(test_se), 
        .CLK(n1612), .Q(\mem0[208][7] ), .QN(n23929) );
  SDFFX1 \mem0_reg[208][6]  ( .D(n18226), .SI(\mem0[208][5] ), .SE(test_se), 
        .CLK(n1612), .Q(\mem0[208][6] ), .QN(n23930) );
  SDFFX1 \mem0_reg[208][5]  ( .D(n18225), .SI(\mem0[208][4] ), .SE(test_se), 
        .CLK(n1612), .Q(\mem0[208][5] ), .QN(n23931) );
  SDFFX1 \mem0_reg[208][4]  ( .D(n18224), .SI(\mem0[208][3] ), .SE(test_se), 
        .CLK(n1612), .Q(\mem0[208][4] ), .QN(n23932) );
  SDFFX1 \mem0_reg[208][3]  ( .D(n18223), .SI(\mem0[208][2] ), .SE(test_se), 
        .CLK(n1612), .Q(\mem0[208][3] ), .QN(n23933) );
  SDFFX1 \mem0_reg[208][2]  ( .D(n18222), .SI(\mem0[208][1] ), .SE(test_se), 
        .CLK(n1612), .Q(\mem0[208][2] ), .QN(n23934) );
  SDFFX1 \mem0_reg[208][1]  ( .D(n18221), .SI(\mem0[208][0] ), .SE(test_se), 
        .CLK(n1613), .Q(\mem0[208][1] ), .QN(n23935) );
  SDFFX1 \mem0_reg[208][0]  ( .D(n18220), .SI(\mem0[207][7] ), .SE(test_se), 
        .CLK(n1613), .Q(\mem0[208][0] ), .QN(n23936) );
  SDFFX1 \mem0_reg[207][7]  ( .D(n18219), .SI(\mem0[207][6] ), .SE(test_se), 
        .CLK(n1613), .Q(\mem0[207][7] ), .QN(n23937) );
  SDFFX1 \mem0_reg[207][6]  ( .D(n18218), .SI(\mem0[207][5] ), .SE(test_se), 
        .CLK(n1613), .Q(\mem0[207][6] ), .QN(n23938) );
  SDFFX1 \mem0_reg[207][5]  ( .D(n18217), .SI(\mem0[207][4] ), .SE(test_se), 
        .CLK(n1613), .Q(\mem0[207][5] ), .QN(n23939) );
  SDFFX1 \mem0_reg[207][4]  ( .D(n18216), .SI(\mem0[207][3] ), .SE(test_se), 
        .CLK(n1613), .Q(\mem0[207][4] ), .QN(n23940) );
  SDFFX1 \mem0_reg[207][3]  ( .D(n18215), .SI(\mem0[207][2] ), .SE(test_se), 
        .CLK(n1613), .Q(\mem0[207][3] ), .QN(n23941) );
  SDFFX1 \mem0_reg[207][2]  ( .D(n18214), .SI(\mem0[207][1] ), .SE(test_se), 
        .CLK(n1613), .Q(\mem0[207][2] ), .QN(n23942) );
  SDFFX1 \mem0_reg[207][1]  ( .D(n18213), .SI(\mem0[207][0] ), .SE(test_se), 
        .CLK(n1613), .Q(\mem0[207][1] ), .QN(n23943) );
  SDFFX1 \mem0_reg[207][0]  ( .D(n18212), .SI(\mem0[206][7] ), .SE(test_se), 
        .CLK(n1613), .Q(\mem0[207][0] ), .QN(n23944) );
  SDFFX1 \mem0_reg[206][7]  ( .D(n18211), .SI(\mem0[206][6] ), .SE(test_se), 
        .CLK(n1613), .Q(\mem0[206][7] ), .QN(n23945) );
  SDFFX1 \mem0_reg[206][6]  ( .D(n18210), .SI(\mem0[206][5] ), .SE(test_se), 
        .CLK(n1613), .Q(\mem0[206][6] ), .QN(n23946) );
  SDFFX1 \mem0_reg[206][5]  ( .D(n18209), .SI(\mem0[206][4] ), .SE(test_se), 
        .CLK(n1614), .Q(\mem0[206][5] ), .QN(n23947) );
  SDFFX1 \mem0_reg[206][4]  ( .D(n18208), .SI(\mem0[206][3] ), .SE(test_se), 
        .CLK(n1614), .Q(\mem0[206][4] ), .QN(n23948) );
  SDFFX1 \mem0_reg[206][3]  ( .D(n18207), .SI(\mem0[206][2] ), .SE(test_se), 
        .CLK(n1614), .Q(\mem0[206][3] ), .QN(n23949) );
  SDFFX1 \mem0_reg[206][2]  ( .D(n18206), .SI(\mem0[206][1] ), .SE(test_se), 
        .CLK(n1614), .Q(\mem0[206][2] ), .QN(n23950) );
  SDFFX1 \mem0_reg[206][1]  ( .D(n18205), .SI(\mem0[206][0] ), .SE(test_se), 
        .CLK(n1614), .Q(\mem0[206][1] ), .QN(n23951) );
  SDFFX1 \mem0_reg[206][0]  ( .D(n18204), .SI(\mem0[205][7] ), .SE(test_se), 
        .CLK(n1614), .Q(\mem0[206][0] ), .QN(n23952) );
  SDFFX1 \mem0_reg[205][7]  ( .D(n18203), .SI(\mem0[205][6] ), .SE(test_se), 
        .CLK(n1614), .Q(\mem0[205][7] ), .QN(n23953) );
  SDFFX1 \mem0_reg[205][6]  ( .D(n18202), .SI(\mem0[205][5] ), .SE(test_se), 
        .CLK(n1614), .Q(\mem0[205][6] ), .QN(n23954) );
  SDFFX1 \mem0_reg[205][5]  ( .D(n18201), .SI(\mem0[205][4] ), .SE(test_se), 
        .CLK(n1614), .Q(\mem0[205][5] ), .QN(n23955) );
  SDFFX1 \mem0_reg[205][4]  ( .D(n18200), .SI(\mem0[205][3] ), .SE(test_se), 
        .CLK(n1614), .Q(\mem0[205][4] ), .QN(n23956) );
  SDFFX1 \mem0_reg[205][3]  ( .D(n18199), .SI(\mem0[205][2] ), .SE(test_se), 
        .CLK(n1614), .Q(\mem0[205][3] ), .QN(n23957) );
  SDFFX1 \mem0_reg[205][2]  ( .D(n18198), .SI(\mem0[205][1] ), .SE(test_se), 
        .CLK(n1614), .Q(\mem0[205][2] ), .QN(n23958) );
  SDFFX1 \mem0_reg[205][1]  ( .D(n18197), .SI(\mem0[205][0] ), .SE(test_se), 
        .CLK(n1615), .Q(\mem0[205][1] ), .QN(n23959) );
  SDFFX1 \mem0_reg[205][0]  ( .D(n18196), .SI(\mem0[204][7] ), .SE(test_se), 
        .CLK(n1615), .Q(\mem0[205][0] ), .QN(n23960) );
  SDFFX1 \mem0_reg[204][7]  ( .D(n18195), .SI(\mem0[204][6] ), .SE(test_se), 
        .CLK(n1615), .Q(\mem0[204][7] ), .QN(n23961) );
  SDFFX1 \mem0_reg[204][6]  ( .D(n18194), .SI(\mem0[204][5] ), .SE(test_se), 
        .CLK(n1615), .Q(\mem0[204][6] ), .QN(n23962) );
  SDFFX1 \mem0_reg[204][5]  ( .D(n18193), .SI(\mem0[204][4] ), .SE(test_se), 
        .CLK(n1615), .Q(\mem0[204][5] ), .QN(n23963) );
  SDFFX1 \mem0_reg[204][4]  ( .D(n18192), .SI(\mem0[204][3] ), .SE(test_se), 
        .CLK(n1615), .Q(\mem0[204][4] ), .QN(n23964) );
  SDFFX1 \mem0_reg[204][3]  ( .D(n18191), .SI(\mem0[204][2] ), .SE(test_se), 
        .CLK(n1615), .Q(\mem0[204][3] ), .QN(n23965) );
  SDFFX1 \mem0_reg[204][2]  ( .D(n18190), .SI(\mem0[204][1] ), .SE(test_se), 
        .CLK(n1615), .Q(\mem0[204][2] ), .QN(n23966) );
  SDFFX1 \mem0_reg[204][1]  ( .D(n18189), .SI(\mem0[204][0] ), .SE(test_se), 
        .CLK(n1615), .Q(\mem0[204][1] ), .QN(n23967) );
  SDFFX1 \mem0_reg[204][0]  ( .D(n18188), .SI(\mem0[203][7] ), .SE(test_se), 
        .CLK(n1615), .Q(\mem0[204][0] ), .QN(n23968) );
  SDFFX1 \mem0_reg[203][7]  ( .D(n18187), .SI(\mem0[203][6] ), .SE(test_se), 
        .CLK(n1615), .Q(\mem0[203][7] ), .QN(n23969) );
  SDFFX1 \mem0_reg[203][6]  ( .D(n18186), .SI(\mem0[203][5] ), .SE(test_se), 
        .CLK(n1615), .Q(\mem0[203][6] ), .QN(n23970) );
  SDFFX1 \mem0_reg[203][5]  ( .D(n18185), .SI(\mem0[203][4] ), .SE(test_se), 
        .CLK(n1616), .Q(\mem0[203][5] ), .QN(n23971) );
  SDFFX1 \mem0_reg[203][4]  ( .D(n18184), .SI(\mem0[203][3] ), .SE(test_se), 
        .CLK(n1616), .Q(\mem0[203][4] ), .QN(n23972) );
  SDFFX1 \mem0_reg[203][3]  ( .D(n18183), .SI(\mem0[203][2] ), .SE(test_se), 
        .CLK(n1616), .Q(\mem0[203][3] ), .QN(n23973) );
  SDFFX1 \mem0_reg[203][2]  ( .D(n18182), .SI(\mem0[203][1] ), .SE(test_se), 
        .CLK(n1616), .Q(\mem0[203][2] ), .QN(n23974) );
  SDFFX1 \mem0_reg[203][1]  ( .D(n18181), .SI(\mem0[203][0] ), .SE(test_se), 
        .CLK(n1616), .Q(\mem0[203][1] ), .QN(n23975) );
  SDFFX1 \mem0_reg[203][0]  ( .D(n18180), .SI(\mem0[202][7] ), .SE(test_se), 
        .CLK(n1616), .Q(\mem0[203][0] ), .QN(n23976) );
  SDFFX1 \mem0_reg[202][7]  ( .D(n18179), .SI(\mem0[202][6] ), .SE(test_se), 
        .CLK(n1616), .Q(\mem0[202][7] ), .QN(n23977) );
  SDFFX1 \mem0_reg[202][6]  ( .D(n18178), .SI(\mem0[202][5] ), .SE(test_se), 
        .CLK(n1616), .Q(\mem0[202][6] ), .QN(n23978) );
  SDFFX1 \mem0_reg[202][5]  ( .D(n18177), .SI(\mem0[202][4] ), .SE(test_se), 
        .CLK(n1616), .Q(\mem0[202][5] ), .QN(n23979) );
  SDFFX1 \mem0_reg[202][4]  ( .D(n18176), .SI(\mem0[202][3] ), .SE(test_se), 
        .CLK(n1616), .Q(\mem0[202][4] ), .QN(n23980) );
  SDFFX1 \mem0_reg[202][3]  ( .D(n18175), .SI(\mem0[202][2] ), .SE(test_se), 
        .CLK(n1616), .Q(\mem0[202][3] ), .QN(n23981) );
  SDFFX1 \mem0_reg[202][2]  ( .D(n18174), .SI(\mem0[202][1] ), .SE(test_se), 
        .CLK(n1616), .Q(\mem0[202][2] ), .QN(n23982) );
  SDFFX1 \mem0_reg[202][1]  ( .D(n18173), .SI(\mem0[202][0] ), .SE(test_se), 
        .CLK(n1617), .Q(\mem0[202][1] ), .QN(n23983) );
  SDFFX1 \mem0_reg[202][0]  ( .D(n18172), .SI(\mem0[201][7] ), .SE(test_se), 
        .CLK(n1617), .Q(\mem0[202][0] ), .QN(n23984) );
  SDFFX1 \mem0_reg[201][7]  ( .D(n18171), .SI(\mem0[201][6] ), .SE(test_se), 
        .CLK(n1617), .Q(\mem0[201][7] ), .QN(n23985) );
  SDFFX1 \mem0_reg[201][6]  ( .D(n18170), .SI(\mem0[201][5] ), .SE(test_se), 
        .CLK(n1617), .Q(\mem0[201][6] ), .QN(n23986) );
  SDFFX1 \mem0_reg[201][5]  ( .D(n18169), .SI(\mem0[201][4] ), .SE(test_se), 
        .CLK(n1617), .Q(\mem0[201][5] ), .QN(n23987) );
  SDFFX1 \mem0_reg[201][4]  ( .D(n18168), .SI(\mem0[201][3] ), .SE(test_se), 
        .CLK(n1617), .Q(\mem0[201][4] ), .QN(n23988) );
  SDFFX1 \mem0_reg[201][3]  ( .D(n18167), .SI(\mem0[201][2] ), .SE(test_se), 
        .CLK(n1617), .Q(\mem0[201][3] ), .QN(n23989) );
  SDFFX1 \mem0_reg[201][2]  ( .D(n18166), .SI(\mem0[201][1] ), .SE(test_se), 
        .CLK(n1617), .Q(\mem0[201][2] ), .QN(n23990) );
  SDFFX1 \mem0_reg[201][1]  ( .D(n18165), .SI(\mem0[201][0] ), .SE(test_se), 
        .CLK(n1617), .Q(\mem0[201][1] ), .QN(n23991) );
  SDFFX1 \mem0_reg[201][0]  ( .D(n18164), .SI(\mem0[200][7] ), .SE(test_se), 
        .CLK(n1617), .Q(\mem0[201][0] ), .QN(n23992) );
  SDFFX1 \mem0_reg[200][7]  ( .D(n18163), .SI(\mem0[200][6] ), .SE(test_se), 
        .CLK(n1617), .Q(\mem0[200][7] ), .QN(n23993) );
  SDFFX1 \mem0_reg[200][6]  ( .D(n18162), .SI(\mem0[200][5] ), .SE(test_se), 
        .CLK(n1617), .Q(\mem0[200][6] ), .QN(n23994) );
  SDFFX1 \mem0_reg[200][5]  ( .D(n18161), .SI(\mem0[200][4] ), .SE(test_se), 
        .CLK(n1618), .Q(\mem0[200][5] ), .QN(n23995) );
  SDFFX1 \mem0_reg[200][4]  ( .D(n18160), .SI(\mem0[200][3] ), .SE(test_se), 
        .CLK(n1618), .Q(\mem0[200][4] ), .QN(n23996) );
  SDFFX1 \mem0_reg[200][3]  ( .D(n18159), .SI(\mem0[200][2] ), .SE(test_se), 
        .CLK(n1618), .Q(\mem0[200][3] ), .QN(n23997) );
  SDFFX1 \mem0_reg[200][2]  ( .D(n18158), .SI(\mem0[200][1] ), .SE(test_se), 
        .CLK(n1618), .Q(\mem0[200][2] ), .QN(n23998) );
  SDFFX1 \mem0_reg[200][1]  ( .D(n18157), .SI(\mem0[200][0] ), .SE(test_se), 
        .CLK(n1618), .Q(\mem0[200][1] ), .QN(n23999) );
  SDFFX1 \mem0_reg[200][0]  ( .D(n18156), .SI(\mem0[199][7] ), .SE(test_se), 
        .CLK(n1618), .Q(\mem0[200][0] ), .QN(n24000) );
  SDFFX1 \mem0_reg[199][7]  ( .D(n18155), .SI(\mem0[199][6] ), .SE(test_se), 
        .CLK(n1618), .Q(\mem0[199][7] ), .QN(n24001) );
  SDFFX1 \mem0_reg[199][6]  ( .D(n18154), .SI(\mem0[199][5] ), .SE(test_se), 
        .CLK(n1618), .Q(\mem0[199][6] ), .QN(n24002) );
  SDFFX1 \mem0_reg[199][5]  ( .D(n18153), .SI(\mem0[199][4] ), .SE(test_se), 
        .CLK(n1618), .Q(\mem0[199][5] ), .QN(n24003) );
  SDFFX1 \mem0_reg[199][4]  ( .D(n18152), .SI(\mem0[199][3] ), .SE(test_se), 
        .CLK(n1618), .Q(\mem0[199][4] ), .QN(n24004) );
  SDFFX1 \mem0_reg[199][3]  ( .D(n18151), .SI(\mem0[199][2] ), .SE(test_se), 
        .CLK(n1618), .Q(\mem0[199][3] ), .QN(n24005) );
  SDFFX1 \mem0_reg[199][2]  ( .D(n18150), .SI(\mem0[199][1] ), .SE(test_se), 
        .CLK(n1618), .Q(\mem0[199][2] ), .QN(n24006) );
  SDFFX1 \mem0_reg[199][1]  ( .D(n18149), .SI(\mem0[199][0] ), .SE(test_se), 
        .CLK(n1619), .Q(\mem0[199][1] ), .QN(n24007) );
  SDFFX1 \mem0_reg[199][0]  ( .D(n18148), .SI(\mem0[198][7] ), .SE(test_se), 
        .CLK(n1619), .Q(\mem0[199][0] ), .QN(n24008) );
  SDFFX1 \mem0_reg[198][7]  ( .D(n18147), .SI(\mem0[198][6] ), .SE(test_se), 
        .CLK(n1619), .Q(\mem0[198][7] ), .QN(n24009) );
  SDFFX1 \mem0_reg[198][6]  ( .D(n18146), .SI(\mem0[198][5] ), .SE(test_se), 
        .CLK(n1619), .Q(\mem0[198][6] ), .QN(n24010) );
  SDFFX1 \mem0_reg[198][5]  ( .D(n18145), .SI(\mem0[198][4] ), .SE(test_se), 
        .CLK(n1619), .Q(\mem0[198][5] ), .QN(n24011) );
  SDFFX1 \mem0_reg[198][4]  ( .D(n18144), .SI(\mem0[198][3] ), .SE(test_se), 
        .CLK(n1619), .Q(\mem0[198][4] ), .QN(n24012) );
  SDFFX1 \mem0_reg[198][3]  ( .D(n18143), .SI(\mem0[198][2] ), .SE(test_se), 
        .CLK(n1619), .Q(\mem0[198][3] ), .QN(n24013) );
  SDFFX1 \mem0_reg[198][2]  ( .D(n18142), .SI(\mem0[198][1] ), .SE(test_se), 
        .CLK(n1619), .Q(\mem0[198][2] ), .QN(n24014) );
  SDFFX1 \mem0_reg[198][1]  ( .D(n18141), .SI(\mem0[198][0] ), .SE(test_se), 
        .CLK(n1619), .Q(\mem0[198][1] ), .QN(n24015) );
  SDFFX1 \mem0_reg[198][0]  ( .D(n18140), .SI(\mem0[197][7] ), .SE(test_se), 
        .CLK(n1619), .Q(\mem0[198][0] ), .QN(n24016) );
  SDFFX1 \mem0_reg[197][7]  ( .D(n18139), .SI(\mem0[197][6] ), .SE(test_se), 
        .CLK(n1619), .Q(\mem0[197][7] ), .QN(n24017) );
  SDFFX1 \mem0_reg[197][6]  ( .D(n18138), .SI(\mem0[197][5] ), .SE(test_se), 
        .CLK(n1619), .Q(\mem0[197][6] ), .QN(n24018) );
  SDFFX1 \mem0_reg[197][5]  ( .D(n18137), .SI(\mem0[197][4] ), .SE(test_se), 
        .CLK(n1620), .Q(\mem0[197][5] ), .QN(n24019) );
  SDFFX1 \mem0_reg[197][4]  ( .D(n18136), .SI(\mem0[197][3] ), .SE(test_se), 
        .CLK(n1620), .Q(\mem0[197][4] ), .QN(n24020) );
  SDFFX1 \mem0_reg[197][3]  ( .D(n18135), .SI(\mem0[197][2] ), .SE(test_se), 
        .CLK(n1620), .Q(\mem0[197][3] ), .QN(n24021) );
  SDFFX1 \mem0_reg[197][2]  ( .D(n18134), .SI(\mem0[197][1] ), .SE(test_se), 
        .CLK(n1620), .Q(\mem0[197][2] ), .QN(n24022) );
  SDFFX1 \mem0_reg[197][1]  ( .D(n18133), .SI(\mem0[197][0] ), .SE(test_se), 
        .CLK(n1620), .Q(\mem0[197][1] ), .QN(n24023) );
  SDFFX1 \mem0_reg[197][0]  ( .D(n18132), .SI(\mem0[196][7] ), .SE(test_se), 
        .CLK(n1620), .Q(\mem0[197][0] ), .QN(n24024) );
  SDFFX1 \mem0_reg[196][7]  ( .D(n18131), .SI(\mem0[196][6] ), .SE(test_se), 
        .CLK(n1620), .Q(\mem0[196][7] ), .QN(n24025) );
  SDFFX1 \mem0_reg[196][6]  ( .D(n18130), .SI(\mem0[196][5] ), .SE(test_se), 
        .CLK(n1620), .Q(\mem0[196][6] ), .QN(n24026) );
  SDFFX1 \mem0_reg[196][5]  ( .D(n18129), .SI(\mem0[196][4] ), .SE(test_se), 
        .CLK(n1620), .Q(\mem0[196][5] ), .QN(n24027) );
  SDFFX1 \mem0_reg[196][4]  ( .D(n18128), .SI(\mem0[196][3] ), .SE(test_se), 
        .CLK(n1620), .Q(\mem0[196][4] ), .QN(n24028) );
  SDFFX1 \mem0_reg[196][3]  ( .D(n18127), .SI(\mem0[196][2] ), .SE(test_se), 
        .CLK(n1620), .Q(\mem0[196][3] ), .QN(n24029) );
  SDFFX1 \mem0_reg[196][2]  ( .D(n18126), .SI(\mem0[196][1] ), .SE(test_se), 
        .CLK(n1620), .Q(\mem0[196][2] ), .QN(n24030) );
  SDFFX1 \mem0_reg[196][1]  ( .D(n18125), .SI(\mem0[196][0] ), .SE(test_se), 
        .CLK(n1621), .Q(\mem0[196][1] ), .QN(n24031) );
  SDFFX1 \mem0_reg[196][0]  ( .D(n18124), .SI(\mem0[195][7] ), .SE(test_se), 
        .CLK(n1621), .Q(\mem0[196][0] ), .QN(n24032) );
  SDFFX1 \mem0_reg[195][7]  ( .D(n18123), .SI(\mem0[195][6] ), .SE(test_se), 
        .CLK(n1621), .Q(\mem0[195][7] ), .QN(n24033) );
  SDFFX1 \mem0_reg[195][6]  ( .D(n18122), .SI(\mem0[195][5] ), .SE(test_se), 
        .CLK(n1621), .Q(\mem0[195][6] ), .QN(n24034) );
  SDFFX1 \mem0_reg[195][5]  ( .D(n18121), .SI(\mem0[195][4] ), .SE(test_se), 
        .CLK(n1621), .Q(\mem0[195][5] ), .QN(n24035) );
  SDFFX1 \mem0_reg[195][4]  ( .D(n18120), .SI(\mem0[195][3] ), .SE(test_se), 
        .CLK(n1621), .Q(\mem0[195][4] ), .QN(n24036) );
  SDFFX1 \mem0_reg[195][3]  ( .D(n18119), .SI(\mem0[195][2] ), .SE(test_se), 
        .CLK(n1621), .Q(\mem0[195][3] ), .QN(n24037) );
  SDFFX1 \mem0_reg[195][2]  ( .D(n18118), .SI(\mem0[195][1] ), .SE(test_se), 
        .CLK(n1621), .Q(\mem0[195][2] ), .QN(n24038) );
  SDFFX1 \mem0_reg[195][1]  ( .D(n18117), .SI(\mem0[195][0] ), .SE(test_se), 
        .CLK(n1621), .Q(\mem0[195][1] ), .QN(n24039) );
  SDFFX1 \mem0_reg[195][0]  ( .D(n18116), .SI(\mem0[194][7] ), .SE(test_se), 
        .CLK(n1621), .Q(\mem0[195][0] ), .QN(n24040) );
  SDFFX1 \mem0_reg[194][7]  ( .D(n18115), .SI(\mem0[194][6] ), .SE(test_se), 
        .CLK(n1621), .Q(\mem0[194][7] ), .QN(n24041) );
  SDFFX1 \mem0_reg[194][6]  ( .D(n18114), .SI(\mem0[194][5] ), .SE(test_se), 
        .CLK(n1621), .Q(\mem0[194][6] ), .QN(n24042) );
  SDFFX1 \mem0_reg[194][5]  ( .D(n18113), .SI(\mem0[194][4] ), .SE(test_se), 
        .CLK(n1622), .Q(\mem0[194][5] ), .QN(n24043) );
  SDFFX1 \mem0_reg[194][4]  ( .D(n18112), .SI(\mem0[194][3] ), .SE(test_se), 
        .CLK(n1622), .Q(\mem0[194][4] ), .QN(n24044) );
  SDFFX1 \mem0_reg[194][3]  ( .D(n18111), .SI(\mem0[194][2] ), .SE(test_se), 
        .CLK(n1622), .Q(\mem0[194][3] ), .QN(n24045) );
  SDFFX1 \mem0_reg[194][2]  ( .D(n18110), .SI(\mem0[194][1] ), .SE(test_se), 
        .CLK(n1622), .Q(\mem0[194][2] ), .QN(n24046) );
  SDFFX1 \mem0_reg[194][1]  ( .D(n18109), .SI(\mem0[194][0] ), .SE(test_se), 
        .CLK(n1622), .Q(\mem0[194][1] ), .QN(n24047) );
  SDFFX1 \mem0_reg[194][0]  ( .D(n18108), .SI(\mem0[193][7] ), .SE(test_se), 
        .CLK(n1622), .Q(\mem0[194][0] ), .QN(n24048) );
  SDFFX1 \mem0_reg[193][7]  ( .D(n18107), .SI(\mem0[193][6] ), .SE(test_se), 
        .CLK(n1622), .Q(\mem0[193][7] ), .QN(n24049) );
  SDFFX1 \mem0_reg[193][6]  ( .D(n18106), .SI(\mem0[193][5] ), .SE(test_se), 
        .CLK(n1622), .Q(\mem0[193][6] ), .QN(n24050) );
  SDFFX1 \mem0_reg[193][5]  ( .D(n18105), .SI(\mem0[193][4] ), .SE(test_se), 
        .CLK(n1622), .Q(\mem0[193][5] ), .QN(n24051) );
  SDFFX1 \mem0_reg[193][4]  ( .D(n18104), .SI(\mem0[193][3] ), .SE(test_se), 
        .CLK(n1622), .Q(\mem0[193][4] ), .QN(n24052) );
  SDFFX1 \mem0_reg[193][3]  ( .D(n18103), .SI(\mem0[193][2] ), .SE(test_se), 
        .CLK(n1622), .Q(\mem0[193][3] ), .QN(n24053) );
  SDFFX1 \mem0_reg[193][2]  ( .D(n18102), .SI(\mem0[193][1] ), .SE(test_se), 
        .CLK(n1622), .Q(\mem0[193][2] ), .QN(n24054) );
  SDFFX1 \mem0_reg[193][1]  ( .D(n18101), .SI(\mem0[193][0] ), .SE(test_se), 
        .CLK(n1623), .Q(\mem0[193][1] ), .QN(n24055) );
  SDFFX1 \mem0_reg[193][0]  ( .D(n18100), .SI(\mem0[192][7] ), .SE(test_se), 
        .CLK(n1623), .Q(\mem0[193][0] ), .QN(n24056) );
  SDFFX1 \mem0_reg[192][7]  ( .D(n18099), .SI(\mem0[192][6] ), .SE(test_se), 
        .CLK(n1623), .Q(\mem0[192][7] ), .QN(n24057) );
  SDFFX1 \mem0_reg[192][6]  ( .D(n18098), .SI(\mem0[192][5] ), .SE(test_se), 
        .CLK(n1623), .Q(\mem0[192][6] ), .QN(n24058) );
  SDFFX1 \mem0_reg[192][5]  ( .D(n18097), .SI(\mem0[192][4] ), .SE(test_se), 
        .CLK(n1623), .Q(\mem0[192][5] ), .QN(n24059) );
  SDFFX1 \mem0_reg[192][4]  ( .D(n18096), .SI(\mem0[192][3] ), .SE(test_se), 
        .CLK(n1623), .Q(\mem0[192][4] ), .QN(n24060) );
  SDFFX1 \mem0_reg[192][3]  ( .D(n18095), .SI(\mem0[192][2] ), .SE(test_se), 
        .CLK(n1623), .Q(\mem0[192][3] ), .QN(n24061) );
  SDFFX1 \mem0_reg[192][2]  ( .D(n18094), .SI(\mem0[192][1] ), .SE(test_se), 
        .CLK(n1623), .Q(\mem0[192][2] ), .QN(n24062) );
  SDFFX1 \mem0_reg[192][1]  ( .D(n18093), .SI(\mem0[192][0] ), .SE(test_se), 
        .CLK(n1623), .Q(\mem0[192][1] ), .QN(n24063) );
  SDFFX1 \mem0_reg[192][0]  ( .D(n18092), .SI(\mem0[191][7] ), .SE(test_se), 
        .CLK(n1623), .Q(\mem0[192][0] ), .QN(n24064) );
  SDFFX1 \mem0_reg[191][7]  ( .D(n18091), .SI(\mem0[191][6] ), .SE(test_se), 
        .CLK(n1623), .Q(\mem0[191][7] ), .QN(n24065) );
  SDFFX1 \mem0_reg[191][6]  ( .D(n18090), .SI(\mem0[191][5] ), .SE(test_se), 
        .CLK(n1623), .Q(\mem0[191][6] ), .QN(n24066) );
  SDFFX1 \mem0_reg[191][5]  ( .D(n18089), .SI(\mem0[191][4] ), .SE(test_se), 
        .CLK(n1624), .Q(\mem0[191][5] ), .QN(n24067) );
  SDFFX1 \mem0_reg[191][4]  ( .D(n18088), .SI(\mem0[191][3] ), .SE(test_se), 
        .CLK(n1624), .Q(\mem0[191][4] ), .QN(n24068) );
  SDFFX1 \mem0_reg[191][3]  ( .D(n18087), .SI(\mem0[191][2] ), .SE(test_se), 
        .CLK(n1624), .Q(\mem0[191][3] ), .QN(n24069) );
  SDFFX1 \mem0_reg[191][2]  ( .D(n18086), .SI(\mem0[191][1] ), .SE(test_se), 
        .CLK(n1624), .Q(\mem0[191][2] ), .QN(n24070) );
  SDFFX1 \mem0_reg[191][1]  ( .D(n18085), .SI(\mem0[191][0] ), .SE(test_se), 
        .CLK(n1624), .Q(\mem0[191][1] ), .QN(n24071) );
  SDFFX1 \mem0_reg[191][0]  ( .D(n18084), .SI(\mem0[190][7] ), .SE(test_se), 
        .CLK(n1624), .Q(\mem0[191][0] ), .QN(n24072) );
  SDFFX1 \mem0_reg[190][7]  ( .D(n18083), .SI(\mem0[190][6] ), .SE(test_se), 
        .CLK(n1624), .Q(\mem0[190][7] ), .QN(n24073) );
  SDFFX1 \mem0_reg[190][6]  ( .D(n18082), .SI(\mem0[190][5] ), .SE(test_se), 
        .CLK(n1624), .Q(\mem0[190][6] ), .QN(n24074) );
  SDFFX1 \mem0_reg[190][5]  ( .D(n18081), .SI(\mem0[190][4] ), .SE(test_se), 
        .CLK(n1624), .Q(\mem0[190][5] ), .QN(n24075) );
  SDFFX1 \mem0_reg[190][4]  ( .D(n18080), .SI(\mem0[190][3] ), .SE(test_se), 
        .CLK(n1624), .Q(\mem0[190][4] ), .QN(n24076) );
  SDFFX1 \mem0_reg[190][3]  ( .D(n18079), .SI(\mem0[190][2] ), .SE(test_se), 
        .CLK(n1624), .Q(\mem0[190][3] ), .QN(n24077) );
  SDFFX1 \mem0_reg[190][2]  ( .D(n18078), .SI(\mem0[190][1] ), .SE(test_se), 
        .CLK(n1624), .Q(\mem0[190][2] ), .QN(n24078) );
  SDFFX1 \mem0_reg[190][1]  ( .D(n18077), .SI(\mem0[190][0] ), .SE(test_se), 
        .CLK(n1625), .Q(\mem0[190][1] ), .QN(n24079) );
  SDFFX1 \mem0_reg[190][0]  ( .D(n18076), .SI(\mem0[189][7] ), .SE(test_se), 
        .CLK(n1625), .Q(\mem0[190][0] ), .QN(n24080) );
  SDFFX1 \mem0_reg[189][7]  ( .D(n18075), .SI(\mem0[189][6] ), .SE(test_se), 
        .CLK(n1625), .Q(\mem0[189][7] ), .QN(n24081) );
  SDFFX1 \mem0_reg[189][6]  ( .D(n18074), .SI(\mem0[189][5] ), .SE(test_se), 
        .CLK(n1625), .Q(\mem0[189][6] ), .QN(n24082) );
  SDFFX1 \mem0_reg[189][5]  ( .D(n18073), .SI(\mem0[189][4] ), .SE(test_se), 
        .CLK(n1625), .Q(\mem0[189][5] ), .QN(n24083) );
  SDFFX1 \mem0_reg[189][4]  ( .D(n18072), .SI(\mem0[189][3] ), .SE(test_se), 
        .CLK(n1625), .Q(\mem0[189][4] ), .QN(n24084) );
  SDFFX1 \mem0_reg[189][3]  ( .D(n18071), .SI(\mem0[189][2] ), .SE(test_se), 
        .CLK(n1625), .Q(\mem0[189][3] ), .QN(n24085) );
  SDFFX1 \mem0_reg[189][2]  ( .D(n18070), .SI(\mem0[189][1] ), .SE(test_se), 
        .CLK(n1625), .Q(\mem0[189][2] ), .QN(n24086) );
  SDFFX1 \mem0_reg[189][1]  ( .D(n18069), .SI(\mem0[189][0] ), .SE(test_se), 
        .CLK(n1625), .Q(\mem0[189][1] ), .QN(n24087) );
  SDFFX1 \mem0_reg[189][0]  ( .D(n18068), .SI(\mem0[188][7] ), .SE(test_se), 
        .CLK(n1625), .Q(\mem0[189][0] ), .QN(n24088) );
  SDFFX1 \mem0_reg[188][7]  ( .D(n18067), .SI(\mem0[188][6] ), .SE(test_se), 
        .CLK(n1625), .Q(\mem0[188][7] ), .QN(n24089) );
  SDFFX1 \mem0_reg[188][6]  ( .D(n18066), .SI(\mem0[188][5] ), .SE(test_se), 
        .CLK(n1625), .Q(\mem0[188][6] ), .QN(n24090) );
  SDFFX1 \mem0_reg[188][5]  ( .D(n18065), .SI(\mem0[188][4] ), .SE(test_se), 
        .CLK(n1626), .Q(\mem0[188][5] ), .QN(n24091) );
  SDFFX1 \mem0_reg[188][4]  ( .D(n18064), .SI(\mem0[188][3] ), .SE(test_se), 
        .CLK(n1626), .Q(\mem0[188][4] ), .QN(n24092) );
  SDFFX1 \mem0_reg[188][3]  ( .D(n18063), .SI(\mem0[188][2] ), .SE(test_se), 
        .CLK(n1626), .Q(\mem0[188][3] ), .QN(n24093) );
  SDFFX1 \mem0_reg[188][2]  ( .D(n18062), .SI(\mem0[188][1] ), .SE(test_se), 
        .CLK(n1626), .Q(\mem0[188][2] ), .QN(n24094) );
  SDFFX1 \mem0_reg[188][1]  ( .D(n18061), .SI(\mem0[188][0] ), .SE(test_se), 
        .CLK(n1626), .Q(\mem0[188][1] ), .QN(n24095) );
  SDFFX1 \mem0_reg[188][0]  ( .D(n18060), .SI(\mem0[187][7] ), .SE(test_se), 
        .CLK(n1626), .Q(\mem0[188][0] ), .QN(n24096) );
  SDFFX1 \mem0_reg[187][7]  ( .D(n18059), .SI(\mem0[187][6] ), .SE(test_se), 
        .CLK(n1626), .Q(\mem0[187][7] ), .QN(n24097) );
  SDFFX1 \mem0_reg[187][6]  ( .D(n18058), .SI(\mem0[187][5] ), .SE(test_se), 
        .CLK(n1626), .Q(\mem0[187][6] ), .QN(n24098) );
  SDFFX1 \mem0_reg[187][5]  ( .D(n18057), .SI(\mem0[187][4] ), .SE(test_se), 
        .CLK(n1626), .Q(\mem0[187][5] ), .QN(n24099) );
  SDFFX1 \mem0_reg[187][4]  ( .D(n18056), .SI(\mem0[187][3] ), .SE(test_se), 
        .CLK(n1626), .Q(\mem0[187][4] ), .QN(n24100) );
  SDFFX1 \mem0_reg[187][3]  ( .D(n18055), .SI(\mem0[187][2] ), .SE(test_se), 
        .CLK(n1626), .Q(\mem0[187][3] ), .QN(n24101) );
  SDFFX1 \mem0_reg[187][2]  ( .D(n18054), .SI(\mem0[187][1] ), .SE(test_se), 
        .CLK(n1626), .Q(\mem0[187][2] ), .QN(n24102) );
  SDFFX1 \mem0_reg[187][1]  ( .D(n18053), .SI(\mem0[187][0] ), .SE(test_se), 
        .CLK(n1627), .Q(\mem0[187][1] ), .QN(n24103) );
  SDFFX1 \mem0_reg[187][0]  ( .D(n18052), .SI(\mem0[186][7] ), .SE(test_se), 
        .CLK(n1627), .Q(\mem0[187][0] ), .QN(n24104) );
  SDFFX1 \mem0_reg[186][7]  ( .D(n18051), .SI(\mem0[186][6] ), .SE(test_se), 
        .CLK(n1627), .Q(\mem0[186][7] ), .QN(n24105) );
  SDFFX1 \mem0_reg[186][6]  ( .D(n18050), .SI(test_si3), .SE(test_se), .CLK(
        n1627), .Q(\mem0[186][6] ), .QN(n24106) );
  SDFFX1 \mem0_reg[186][5]  ( .D(n18049), .SI(\mem0[186][4] ), .SE(test_se), 
        .CLK(n1627), .Q(\mem0[186][5] ), .QN(n24107) );
  SDFFX1 \mem0_reg[186][4]  ( .D(n18048), .SI(\mem0[186][3] ), .SE(test_se), 
        .CLK(n1627), .Q(\mem0[186][4] ), .QN(n24108) );
  SDFFX1 \mem0_reg[186][3]  ( .D(n18047), .SI(\mem0[186][2] ), .SE(test_se), 
        .CLK(n1627), .Q(\mem0[186][3] ), .QN(n24109) );
  SDFFX1 \mem0_reg[186][2]  ( .D(n18046), .SI(\mem0[186][1] ), .SE(test_se), 
        .CLK(n1627), .Q(\mem0[186][2] ), .QN(n24110) );
  SDFFX1 \mem0_reg[186][1]  ( .D(n18045), .SI(\mem0[186][0] ), .SE(test_se), 
        .CLK(n1627), .Q(\mem0[186][1] ), .QN(n24111) );
  SDFFX1 \mem0_reg[186][0]  ( .D(n18044), .SI(\mem0[185][7] ), .SE(test_se), 
        .CLK(n1627), .Q(\mem0[186][0] ), .QN(n24112) );
  SDFFX1 \mem0_reg[185][7]  ( .D(n18043), .SI(\mem0[185][6] ), .SE(test_se), 
        .CLK(n1627), .Q(\mem0[185][7] ), .QN(n24113) );
  SDFFX1 \mem0_reg[185][6]  ( .D(n18042), .SI(\mem0[185][5] ), .SE(test_se), 
        .CLK(n1627), .Q(\mem0[185][6] ), .QN(n24114) );
  SDFFX1 \mem0_reg[185][5]  ( .D(n18041), .SI(\mem0[185][4] ), .SE(test_se), 
        .CLK(n1628), .Q(\mem0[185][5] ), .QN(n24115) );
  SDFFX1 \mem0_reg[185][4]  ( .D(n18040), .SI(\mem0[185][3] ), .SE(test_se), 
        .CLK(n1628), .Q(\mem0[185][4] ), .QN(n24116) );
  SDFFX1 \mem0_reg[185][3]  ( .D(n18039), .SI(\mem0[185][2] ), .SE(test_se), 
        .CLK(n1628), .Q(\mem0[185][3] ), .QN(n24117) );
  SDFFX1 \mem0_reg[185][2]  ( .D(n18038), .SI(\mem0[185][1] ), .SE(test_se), 
        .CLK(n1628), .Q(\mem0[185][2] ), .QN(n24118) );
  SDFFX1 \mem0_reg[185][1]  ( .D(n18037), .SI(\mem0[185][0] ), .SE(test_se), 
        .CLK(n1628), .Q(\mem0[185][1] ), .QN(n24119) );
  SDFFX1 \mem0_reg[185][0]  ( .D(n18036), .SI(\mem0[184][7] ), .SE(test_se), 
        .CLK(n1628), .Q(\mem0[185][0] ), .QN(n24120) );
  SDFFX1 \mem0_reg[184][7]  ( .D(n18035), .SI(\mem0[184][6] ), .SE(test_se), 
        .CLK(n1628), .Q(\mem0[184][7] ), .QN(n24121) );
  SDFFX1 \mem0_reg[184][6]  ( .D(n18034), .SI(\mem0[184][5] ), .SE(test_se), 
        .CLK(n1628), .Q(\mem0[184][6] ), .QN(n24122) );
  SDFFX1 \mem0_reg[184][5]  ( .D(n18033), .SI(\mem0[184][4] ), .SE(test_se), 
        .CLK(n1628), .Q(\mem0[184][5] ), .QN(n24123) );
  SDFFX1 \mem0_reg[184][4]  ( .D(n18032), .SI(\mem0[184][3] ), .SE(test_se), 
        .CLK(n1628), .Q(\mem0[184][4] ), .QN(n24124) );
  SDFFX1 \mem0_reg[184][3]  ( .D(n18031), .SI(\mem0[184][2] ), .SE(test_se), 
        .CLK(n1628), .Q(\mem0[184][3] ), .QN(n24125) );
  SDFFX1 \mem0_reg[184][2]  ( .D(n18030), .SI(\mem0[184][1] ), .SE(test_se), 
        .CLK(n1628), .Q(\mem0[184][2] ), .QN(n24126) );
  SDFFX1 \mem0_reg[184][1]  ( .D(n18029), .SI(\mem0[184][0] ), .SE(test_se), 
        .CLK(n1629), .Q(\mem0[184][1] ), .QN(n24127) );
  SDFFX1 \mem0_reg[184][0]  ( .D(n18028), .SI(\mem0[183][7] ), .SE(test_se), 
        .CLK(n1629), .Q(\mem0[184][0] ), .QN(n24128) );
  SDFFX1 \mem0_reg[183][7]  ( .D(n18027), .SI(\mem0[183][6] ), .SE(test_se), 
        .CLK(n1629), .Q(\mem0[183][7] ), .QN(n24129) );
  SDFFX1 \mem0_reg[183][6]  ( .D(n18026), .SI(\mem0[183][5] ), .SE(test_se), 
        .CLK(n1629), .Q(\mem0[183][6] ), .QN(n24130) );
  SDFFX1 \mem0_reg[183][5]  ( .D(n18025), .SI(\mem0[183][4] ), .SE(test_se), 
        .CLK(n1629), .Q(\mem0[183][5] ), .QN(n24131) );
  SDFFX1 \mem0_reg[183][4]  ( .D(n18024), .SI(\mem0[183][3] ), .SE(test_se), 
        .CLK(n1629), .Q(\mem0[183][4] ), .QN(n24132) );
  SDFFX1 \mem0_reg[183][3]  ( .D(n18023), .SI(\mem0[183][2] ), .SE(test_se), 
        .CLK(n1629), .Q(\mem0[183][3] ), .QN(n24133) );
  SDFFX1 \mem0_reg[183][2]  ( .D(n18022), .SI(\mem0[183][1] ), .SE(test_se), 
        .CLK(n1629), .Q(\mem0[183][2] ), .QN(n24134) );
  SDFFX1 \mem0_reg[183][1]  ( .D(n18021), .SI(\mem0[183][0] ), .SE(test_se), 
        .CLK(n1629), .Q(\mem0[183][1] ), .QN(n24135) );
  SDFFX1 \mem0_reg[183][0]  ( .D(n18020), .SI(\mem0[182][7] ), .SE(test_se), 
        .CLK(n1629), .Q(\mem0[183][0] ), .QN(n24136) );
  SDFFX1 \mem0_reg[182][7]  ( .D(n18019), .SI(\mem0[182][6] ), .SE(test_se), 
        .CLK(n1629), .Q(\mem0[182][7] ), .QN(n24137) );
  SDFFX1 \mem0_reg[182][6]  ( .D(n18018), .SI(\mem0[182][5] ), .SE(test_se), 
        .CLK(n1629), .Q(\mem0[182][6] ), .QN(n24138) );
  SDFFX1 \mem0_reg[182][5]  ( .D(n18017), .SI(\mem0[182][4] ), .SE(test_se), 
        .CLK(n1630), .Q(\mem0[182][5] ), .QN(n24139) );
  SDFFX1 \mem0_reg[182][4]  ( .D(n18016), .SI(\mem0[182][3] ), .SE(test_se), 
        .CLK(n1630), .Q(\mem0[182][4] ), .QN(n24140) );
  SDFFX1 \mem0_reg[182][3]  ( .D(n18015), .SI(\mem0[182][2] ), .SE(test_se), 
        .CLK(n1630), .Q(\mem0[182][3] ), .QN(n24141) );
  SDFFX1 \mem0_reg[182][2]  ( .D(n18014), .SI(\mem0[182][1] ), .SE(test_se), 
        .CLK(n1630), .Q(\mem0[182][2] ), .QN(n24142) );
  SDFFX1 \mem0_reg[182][1]  ( .D(n18013), .SI(\mem0[182][0] ), .SE(test_se), 
        .CLK(n1630), .Q(\mem0[182][1] ), .QN(n24143) );
  SDFFX1 \mem0_reg[182][0]  ( .D(n18012), .SI(\mem0[181][7] ), .SE(test_se), 
        .CLK(n1630), .Q(\mem0[182][0] ), .QN(n24144) );
  SDFFX1 \mem0_reg[181][7]  ( .D(n18011), .SI(\mem0[181][6] ), .SE(test_se), 
        .CLK(n1630), .Q(\mem0[181][7] ), .QN(n24145) );
  SDFFX1 \mem0_reg[181][6]  ( .D(n18010), .SI(\mem0[181][5] ), .SE(test_se), 
        .CLK(n1630), .Q(\mem0[181][6] ), .QN(n24146) );
  SDFFX1 \mem0_reg[181][5]  ( .D(n18009), .SI(\mem0[181][4] ), .SE(test_se), 
        .CLK(n1630), .Q(\mem0[181][5] ), .QN(n24147) );
  SDFFX1 \mem0_reg[181][4]  ( .D(n18008), .SI(\mem0[181][3] ), .SE(test_se), 
        .CLK(n1630), .Q(\mem0[181][4] ), .QN(n24148) );
  SDFFX1 \mem0_reg[181][3]  ( .D(n18007), .SI(\mem0[181][2] ), .SE(test_se), 
        .CLK(n1630), .Q(\mem0[181][3] ), .QN(n24149) );
  SDFFX1 \mem0_reg[181][2]  ( .D(n18006), .SI(\mem0[181][1] ), .SE(test_se), 
        .CLK(n1630), .Q(\mem0[181][2] ), .QN(n24150) );
  SDFFX1 \mem0_reg[181][1]  ( .D(n18005), .SI(\mem0[181][0] ), .SE(test_se), 
        .CLK(n1631), .Q(\mem0[181][1] ), .QN(n24151) );
  SDFFX1 \mem0_reg[181][0]  ( .D(n18004), .SI(\mem0[180][7] ), .SE(test_se), 
        .CLK(n1631), .Q(\mem0[181][0] ), .QN(n24152) );
  SDFFX1 \mem0_reg[180][7]  ( .D(n18003), .SI(\mem0[180][6] ), .SE(test_se), 
        .CLK(n1631), .Q(\mem0[180][7] ), .QN(n24153) );
  SDFFX1 \mem0_reg[180][6]  ( .D(n18002), .SI(\mem0[180][5] ), .SE(test_se), 
        .CLK(n1631), .Q(\mem0[180][6] ), .QN(n24154) );
  SDFFX1 \mem0_reg[180][5]  ( .D(n18001), .SI(\mem0[180][4] ), .SE(test_se), 
        .CLK(n1631), .Q(\mem0[180][5] ), .QN(n24155) );
  SDFFX1 \mem0_reg[180][4]  ( .D(n18000), .SI(\mem0[180][3] ), .SE(test_se), 
        .CLK(n1631), .Q(\mem0[180][4] ), .QN(n24156) );
  SDFFX1 \mem0_reg[180][3]  ( .D(n17999), .SI(\mem0[180][2] ), .SE(test_se), 
        .CLK(n1631), .Q(\mem0[180][3] ), .QN(n24157) );
  SDFFX1 \mem0_reg[180][2]  ( .D(n17998), .SI(\mem0[180][1] ), .SE(test_se), 
        .CLK(n1631), .Q(\mem0[180][2] ), .QN(n24158) );
  SDFFX1 \mem0_reg[180][1]  ( .D(n17997), .SI(\mem0[180][0] ), .SE(test_se), 
        .CLK(n1631), .Q(\mem0[180][1] ), .QN(n24159) );
  SDFFX1 \mem0_reg[180][0]  ( .D(n17996), .SI(\mem0[179][7] ), .SE(test_se), 
        .CLK(n1631), .Q(\mem0[180][0] ), .QN(n24160) );
  SDFFX1 \mem0_reg[179][7]  ( .D(n17995), .SI(\mem0[179][6] ), .SE(test_se), 
        .CLK(n1631), .Q(\mem0[179][7] ), .QN(n24161) );
  SDFFX1 \mem0_reg[179][6]  ( .D(n17994), .SI(\mem0[179][5] ), .SE(test_se), 
        .CLK(n1631), .Q(\mem0[179][6] ), .QN(n24162) );
  SDFFX1 \mem0_reg[179][5]  ( .D(n17993), .SI(\mem0[179][4] ), .SE(test_se), 
        .CLK(n1632), .Q(\mem0[179][5] ), .QN(n24163) );
  SDFFX1 \mem0_reg[179][4]  ( .D(n17992), .SI(\mem0[179][3] ), .SE(test_se), 
        .CLK(n1632), .Q(\mem0[179][4] ), .QN(n24164) );
  SDFFX1 \mem0_reg[179][3]  ( .D(n17991), .SI(\mem0[179][2] ), .SE(test_se), 
        .CLK(n1632), .Q(\mem0[179][3] ), .QN(n24165) );
  SDFFX1 \mem0_reg[179][2]  ( .D(n17990), .SI(\mem0[179][1] ), .SE(test_se), 
        .CLK(n1632), .Q(\mem0[179][2] ), .QN(n24166) );
  SDFFX1 \mem0_reg[179][1]  ( .D(n17989), .SI(\mem0[179][0] ), .SE(test_se), 
        .CLK(n1632), .Q(\mem0[179][1] ), .QN(n24167) );
  SDFFX1 \mem0_reg[179][0]  ( .D(n17988), .SI(\mem0[178][7] ), .SE(test_se), 
        .CLK(n1632), .Q(\mem0[179][0] ), .QN(n24168) );
  SDFFX1 \mem0_reg[178][7]  ( .D(n17987), .SI(\mem0[178][6] ), .SE(test_se), 
        .CLK(n1632), .Q(\mem0[178][7] ), .QN(n24169) );
  SDFFX1 \mem0_reg[178][6]  ( .D(n17986), .SI(\mem0[178][5] ), .SE(test_se), 
        .CLK(n1632), .Q(\mem0[178][6] ), .QN(n24170) );
  SDFFX1 \mem0_reg[178][5]  ( .D(n17985), .SI(\mem0[178][4] ), .SE(test_se), 
        .CLK(n1632), .Q(\mem0[178][5] ), .QN(n24171) );
  SDFFX1 \mem0_reg[178][4]  ( .D(n17984), .SI(\mem0[178][3] ), .SE(test_se), 
        .CLK(n1632), .Q(\mem0[178][4] ), .QN(n24172) );
  SDFFX1 \mem0_reg[178][3]  ( .D(n17983), .SI(\mem0[178][2] ), .SE(test_se), 
        .CLK(n1632), .Q(\mem0[178][3] ), .QN(n24173) );
  SDFFX1 \mem0_reg[178][2]  ( .D(n17982), .SI(\mem0[178][1] ), .SE(test_se), 
        .CLK(n1632), .Q(\mem0[178][2] ), .QN(n24174) );
  SDFFX1 \mem0_reg[178][1]  ( .D(n17981), .SI(\mem0[178][0] ), .SE(test_se), 
        .CLK(n1633), .Q(\mem0[178][1] ), .QN(n24175) );
  SDFFX1 \mem0_reg[178][0]  ( .D(n17980), .SI(\mem0[177][7] ), .SE(test_se), 
        .CLK(n1633), .Q(\mem0[178][0] ), .QN(n24176) );
  SDFFX1 \mem0_reg[177][7]  ( .D(n17979), .SI(\mem0[177][6] ), .SE(test_se), 
        .CLK(n1633), .Q(\mem0[177][7] ), .QN(n24177) );
  SDFFX1 \mem0_reg[177][6]  ( .D(n17978), .SI(\mem0[177][5] ), .SE(test_se), 
        .CLK(n1633), .Q(\mem0[177][6] ), .QN(n24178) );
  SDFFX1 \mem0_reg[177][5]  ( .D(n17977), .SI(\mem0[177][4] ), .SE(test_se), 
        .CLK(n1633), .Q(\mem0[177][5] ), .QN(n24179) );
  SDFFX1 \mem0_reg[177][4]  ( .D(n17976), .SI(\mem0[177][3] ), .SE(test_se), 
        .CLK(n1633), .Q(\mem0[177][4] ), .QN(n24180) );
  SDFFX1 \mem0_reg[177][3]  ( .D(n17975), .SI(\mem0[177][2] ), .SE(test_se), 
        .CLK(n1633), .Q(\mem0[177][3] ), .QN(n24181) );
  SDFFX1 \mem0_reg[177][2]  ( .D(n17974), .SI(\mem0[177][1] ), .SE(test_se), 
        .CLK(n1633), .Q(\mem0[177][2] ), .QN(n24182) );
  SDFFX1 \mem0_reg[177][1]  ( .D(n17973), .SI(\mem0[177][0] ), .SE(test_se), 
        .CLK(n1633), .Q(\mem0[177][1] ), .QN(n24183) );
  SDFFX1 \mem0_reg[177][0]  ( .D(n17972), .SI(\mem0[176][7] ), .SE(test_se), 
        .CLK(n1633), .Q(\mem0[177][0] ), .QN(n24184) );
  SDFFX1 \mem0_reg[176][7]  ( .D(n17971), .SI(\mem0[176][6] ), .SE(test_se), 
        .CLK(n1633), .Q(\mem0[176][7] ), .QN(n24185) );
  SDFFX1 \mem0_reg[176][6]  ( .D(n17970), .SI(\mem0[176][5] ), .SE(test_se), 
        .CLK(n1633), .Q(\mem0[176][6] ), .QN(n24186) );
  SDFFX1 \mem0_reg[176][5]  ( .D(n17969), .SI(\mem0[176][4] ), .SE(test_se), 
        .CLK(n1634), .Q(\mem0[176][5] ), .QN(n24187) );
  SDFFX1 \mem0_reg[176][4]  ( .D(n17968), .SI(\mem0[176][3] ), .SE(test_se), 
        .CLK(n1634), .Q(\mem0[176][4] ), .QN(n24188) );
  SDFFX1 \mem0_reg[176][3]  ( .D(n17967), .SI(\mem0[176][2] ), .SE(test_se), 
        .CLK(n1634), .Q(\mem0[176][3] ), .QN(n24189) );
  SDFFX1 \mem0_reg[176][2]  ( .D(n17966), .SI(\mem0[176][1] ), .SE(test_se), 
        .CLK(n1634), .Q(\mem0[176][2] ), .QN(n24190) );
  SDFFX1 \mem0_reg[176][1]  ( .D(n17965), .SI(\mem0[176][0] ), .SE(test_se), 
        .CLK(n1634), .Q(\mem0[176][1] ), .QN(n24191) );
  SDFFX1 \mem0_reg[176][0]  ( .D(n17964), .SI(\mem0[175][7] ), .SE(test_se), 
        .CLK(n1634), .Q(\mem0[176][0] ), .QN(n24192) );
  SDFFX1 \mem0_reg[175][7]  ( .D(n17963), .SI(\mem0[175][6] ), .SE(test_se), 
        .CLK(n1634), .Q(\mem0[175][7] ), .QN(n24193) );
  SDFFX1 \mem0_reg[175][6]  ( .D(n17962), .SI(\mem0[175][5] ), .SE(test_se), 
        .CLK(n1634), .Q(\mem0[175][6] ), .QN(n24194) );
  SDFFX1 \mem0_reg[175][5]  ( .D(n17961), .SI(\mem0[175][4] ), .SE(test_se), 
        .CLK(n1634), .Q(\mem0[175][5] ), .QN(n24195) );
  SDFFX1 \mem0_reg[175][4]  ( .D(n17960), .SI(\mem0[175][3] ), .SE(test_se), 
        .CLK(n1634), .Q(\mem0[175][4] ), .QN(n24196) );
  SDFFX1 \mem0_reg[175][3]  ( .D(n17959), .SI(\mem0[175][2] ), .SE(test_se), 
        .CLK(n1634), .Q(\mem0[175][3] ), .QN(n24197) );
  SDFFX1 \mem0_reg[175][2]  ( .D(n17958), .SI(\mem0[175][1] ), .SE(test_se), 
        .CLK(n1634), .Q(\mem0[175][2] ), .QN(n24198) );
  SDFFX1 \mem0_reg[175][1]  ( .D(n17957), .SI(\mem0[175][0] ), .SE(test_se), 
        .CLK(n1635), .Q(\mem0[175][1] ), .QN(n24199) );
  SDFFX1 \mem0_reg[175][0]  ( .D(n17956), .SI(\mem0[174][7] ), .SE(test_se), 
        .CLK(n1635), .Q(\mem0[175][0] ), .QN(n24200) );
  SDFFX1 \mem0_reg[174][7]  ( .D(n17955), .SI(\mem0[174][6] ), .SE(test_se), 
        .CLK(n1635), .Q(\mem0[174][7] ), .QN(n24201) );
  SDFFX1 \mem0_reg[174][6]  ( .D(n17954), .SI(\mem0[174][5] ), .SE(test_se), 
        .CLK(n1635), .Q(\mem0[174][6] ), .QN(n24202) );
  SDFFX1 \mem0_reg[174][5]  ( .D(n17953), .SI(\mem0[174][4] ), .SE(test_se), 
        .CLK(n1635), .Q(\mem0[174][5] ), .QN(n24203) );
  SDFFX1 \mem0_reg[174][4]  ( .D(n17952), .SI(\mem0[174][3] ), .SE(test_se), 
        .CLK(n1635), .Q(\mem0[174][4] ), .QN(n24204) );
  SDFFX1 \mem0_reg[174][3]  ( .D(n17951), .SI(\mem0[174][2] ), .SE(test_se), 
        .CLK(n1635), .Q(\mem0[174][3] ), .QN(n24205) );
  SDFFX1 \mem0_reg[174][2]  ( .D(n17950), .SI(\mem0[174][1] ), .SE(test_se), 
        .CLK(n1635), .Q(\mem0[174][2] ), .QN(n24206) );
  SDFFX1 \mem0_reg[174][1]  ( .D(n17949), .SI(\mem0[174][0] ), .SE(test_se), 
        .CLK(n1635), .Q(\mem0[174][1] ), .QN(n24207) );
  SDFFX1 \mem0_reg[174][0]  ( .D(n17948), .SI(\mem0[173][7] ), .SE(test_se), 
        .CLK(n1635), .Q(\mem0[174][0] ), .QN(n24208) );
  SDFFX1 \mem0_reg[173][7]  ( .D(n17947), .SI(\mem0[173][6] ), .SE(test_se), 
        .CLK(n1635), .Q(\mem0[173][7] ), .QN(n24209) );
  SDFFX1 \mem0_reg[173][6]  ( .D(n17946), .SI(\mem0[173][5] ), .SE(test_se), 
        .CLK(n1635), .Q(\mem0[173][6] ), .QN(n24210) );
  SDFFX1 \mem0_reg[173][5]  ( .D(n17945), .SI(\mem0[173][4] ), .SE(test_se), 
        .CLK(n1636), .Q(\mem0[173][5] ), .QN(n24211) );
  SDFFX1 \mem0_reg[173][4]  ( .D(n17944), .SI(\mem0[173][3] ), .SE(test_se), 
        .CLK(n1636), .Q(\mem0[173][4] ), .QN(n24212) );
  SDFFX1 \mem0_reg[173][3]  ( .D(n17943), .SI(\mem0[173][2] ), .SE(test_se), 
        .CLK(n1636), .Q(\mem0[173][3] ), .QN(n24213) );
  SDFFX1 \mem0_reg[173][2]  ( .D(n17942), .SI(\mem0[173][1] ), .SE(test_se), 
        .CLK(n1636), .Q(\mem0[173][2] ), .QN(n24214) );
  SDFFX1 \mem0_reg[173][1]  ( .D(n17941), .SI(\mem0[173][0] ), .SE(test_se), 
        .CLK(n1636), .Q(\mem0[173][1] ), .QN(n24215) );
  SDFFX1 \mem0_reg[173][0]  ( .D(n17940), .SI(\mem0[172][7] ), .SE(test_se), 
        .CLK(n1636), .Q(\mem0[173][0] ), .QN(n24216) );
  SDFFX1 \mem0_reg[172][7]  ( .D(n17939), .SI(\mem0[172][6] ), .SE(test_se), 
        .CLK(n1636), .Q(\mem0[172][7] ), .QN(n24217) );
  SDFFX1 \mem0_reg[172][6]  ( .D(n17938), .SI(\mem0[172][5] ), .SE(test_se), 
        .CLK(n1636), .Q(\mem0[172][6] ), .QN(n24218) );
  SDFFX1 \mem0_reg[172][5]  ( .D(n17937), .SI(\mem0[172][4] ), .SE(test_se), 
        .CLK(n1636), .Q(\mem0[172][5] ), .QN(n24219) );
  SDFFX1 \mem0_reg[172][4]  ( .D(n17936), .SI(\mem0[172][3] ), .SE(test_se), 
        .CLK(n1636), .Q(\mem0[172][4] ), .QN(n24220) );
  SDFFX1 \mem0_reg[172][3]  ( .D(n17935), .SI(\mem0[172][2] ), .SE(test_se), 
        .CLK(n1636), .Q(\mem0[172][3] ), .QN(n24221) );
  SDFFX1 \mem0_reg[172][2]  ( .D(n17934), .SI(\mem0[172][1] ), .SE(test_se), 
        .CLK(n1636), .Q(\mem0[172][2] ), .QN(n24222) );
  SDFFX1 \mem0_reg[172][1]  ( .D(n17933), .SI(\mem0[172][0] ), .SE(test_se), 
        .CLK(n1637), .Q(\mem0[172][1] ), .QN(n24223) );
  SDFFX1 \mem0_reg[172][0]  ( .D(n17932), .SI(\mem0[171][7] ), .SE(test_se), 
        .CLK(n1637), .Q(\mem0[172][0] ), .QN(n24224) );
  SDFFX1 \mem0_reg[171][7]  ( .D(n17931), .SI(\mem0[171][6] ), .SE(test_se), 
        .CLK(n1637), .Q(\mem0[171][7] ), .QN(n24225) );
  SDFFX1 \mem0_reg[171][6]  ( .D(n17930), .SI(\mem0[171][5] ), .SE(test_se), 
        .CLK(n1637), .Q(\mem0[171][6] ), .QN(n24226) );
  SDFFX1 \mem0_reg[171][5]  ( .D(n17929), .SI(\mem0[171][4] ), .SE(test_se), 
        .CLK(n1637), .Q(\mem0[171][5] ), .QN(n24227) );
  SDFFX1 \mem0_reg[171][4]  ( .D(n17928), .SI(\mem0[171][3] ), .SE(test_se), 
        .CLK(n1637), .Q(\mem0[171][4] ), .QN(n24228) );
  SDFFX1 \mem0_reg[171][3]  ( .D(n17927), .SI(\mem0[171][2] ), .SE(test_se), 
        .CLK(n1637), .Q(\mem0[171][3] ), .QN(n24229) );
  SDFFX1 \mem0_reg[171][2]  ( .D(n17926), .SI(\mem0[171][1] ), .SE(test_se), 
        .CLK(n1637), .Q(\mem0[171][2] ), .QN(n24230) );
  SDFFX1 \mem0_reg[171][1]  ( .D(n17925), .SI(\mem0[171][0] ), .SE(test_se), 
        .CLK(n1637), .Q(\mem0[171][1] ), .QN(n24231) );
  SDFFX1 \mem0_reg[171][0]  ( .D(n17924), .SI(\mem0[170][7] ), .SE(test_se), 
        .CLK(n1637), .Q(\mem0[171][0] ), .QN(n24232) );
  SDFFX1 \mem0_reg[170][7]  ( .D(n17923), .SI(\mem0[170][6] ), .SE(test_se), 
        .CLK(n1637), .Q(\mem0[170][7] ), .QN(n24233) );
  SDFFX1 \mem0_reg[170][6]  ( .D(n17922), .SI(\mem0[170][5] ), .SE(test_se), 
        .CLK(n1637), .Q(\mem0[170][6] ), .QN(n24234) );
  SDFFX1 \mem0_reg[170][5]  ( .D(n17921), .SI(\mem0[170][4] ), .SE(test_se), 
        .CLK(n1638), .Q(\mem0[170][5] ), .QN(n24235) );
  SDFFX1 \mem0_reg[170][4]  ( .D(n17920), .SI(\mem0[170][3] ), .SE(test_se), 
        .CLK(n1638), .Q(\mem0[170][4] ), .QN(n24236) );
  SDFFX1 \mem0_reg[170][3]  ( .D(n17919), .SI(\mem0[170][2] ), .SE(test_se), 
        .CLK(n1638), .Q(\mem0[170][3] ), .QN(n24237) );
  SDFFX1 \mem0_reg[170][2]  ( .D(n17918), .SI(\mem0[170][1] ), .SE(test_se), 
        .CLK(n1638), .Q(\mem0[170][2] ), .QN(n24238) );
  SDFFX1 \mem0_reg[170][1]  ( .D(n17917), .SI(\mem0[170][0] ), .SE(test_se), 
        .CLK(n1638), .Q(\mem0[170][1] ), .QN(n24239) );
  SDFFX1 \mem0_reg[170][0]  ( .D(n17916), .SI(\mem0[169][7] ), .SE(test_se), 
        .CLK(n1638), .Q(\mem0[170][0] ), .QN(n24240) );
  SDFFX1 \mem0_reg[169][7]  ( .D(n17915), .SI(\mem0[169][6] ), .SE(test_se), 
        .CLK(n1638), .Q(\mem0[169][7] ), .QN(n24241) );
  SDFFX1 \mem0_reg[169][6]  ( .D(n17914), .SI(\mem0[169][5] ), .SE(test_se), 
        .CLK(n1638), .Q(\mem0[169][6] ), .QN(n24242) );
  SDFFX1 \mem0_reg[169][5]  ( .D(n17913), .SI(\mem0[169][4] ), .SE(test_se), 
        .CLK(n1638), .Q(\mem0[169][5] ), .QN(n24243) );
  SDFFX1 \mem0_reg[169][4]  ( .D(n17912), .SI(\mem0[169][3] ), .SE(test_se), 
        .CLK(n1638), .Q(\mem0[169][4] ), .QN(n24244) );
  SDFFX1 \mem0_reg[169][3]  ( .D(n17911), .SI(\mem0[169][2] ), .SE(test_se), 
        .CLK(n1638), .Q(\mem0[169][3] ), .QN(n24245) );
  SDFFX1 \mem0_reg[169][2]  ( .D(n17910), .SI(\mem0[169][1] ), .SE(test_se), 
        .CLK(n1638), .Q(\mem0[169][2] ), .QN(n24246) );
  SDFFX1 \mem0_reg[169][1]  ( .D(n17909), .SI(\mem0[169][0] ), .SE(test_se), 
        .CLK(n1639), .Q(\mem0[169][1] ), .QN(n24247) );
  SDFFX1 \mem0_reg[169][0]  ( .D(n17908), .SI(\mem0[168][7] ), .SE(test_se), 
        .CLK(n1639), .Q(\mem0[169][0] ), .QN(n24248) );
  SDFFX1 \mem0_reg[168][7]  ( .D(n17907), .SI(\mem0[168][6] ), .SE(test_se), 
        .CLK(n1639), .Q(\mem0[168][7] ), .QN(n24249) );
  SDFFX1 \mem0_reg[168][6]  ( .D(n17906), .SI(\mem0[168][5] ), .SE(test_se), 
        .CLK(n1639), .Q(\mem0[168][6] ), .QN(n24250) );
  SDFFX1 \mem0_reg[168][5]  ( .D(n17905), .SI(\mem0[168][4] ), .SE(test_se), 
        .CLK(n1639), .Q(\mem0[168][5] ), .QN(n24251) );
  SDFFX1 \mem0_reg[168][4]  ( .D(n17904), .SI(\mem0[168][3] ), .SE(test_se), 
        .CLK(n1639), .Q(\mem0[168][4] ), .QN(n24252) );
  SDFFX1 \mem0_reg[168][3]  ( .D(n17903), .SI(\mem0[168][2] ), .SE(test_se), 
        .CLK(n1639), .Q(\mem0[168][3] ), .QN(n24253) );
  SDFFX1 \mem0_reg[168][2]  ( .D(n17902), .SI(\mem0[168][1] ), .SE(test_se), 
        .CLK(n1639), .Q(\mem0[168][2] ), .QN(n24254) );
  SDFFX1 \mem0_reg[168][1]  ( .D(n17901), .SI(\mem0[168][0] ), .SE(test_se), 
        .CLK(n1639), .Q(\mem0[168][1] ), .QN(n24255) );
  SDFFX1 \mem0_reg[168][0]  ( .D(n17900), .SI(\mem0[167][7] ), .SE(test_se), 
        .CLK(n1639), .Q(\mem0[168][0] ), .QN(n24256) );
  SDFFX1 \mem0_reg[167][7]  ( .D(n17899), .SI(\mem0[167][6] ), .SE(test_se), 
        .CLK(n1639), .Q(\mem0[167][7] ), .QN(n24257) );
  SDFFX1 \mem0_reg[167][6]  ( .D(n17898), .SI(\mem0[167][5] ), .SE(test_se), 
        .CLK(n1639), .Q(\mem0[167][6] ), .QN(n24258) );
  SDFFX1 \mem0_reg[167][5]  ( .D(n17897), .SI(\mem0[167][4] ), .SE(test_se), 
        .CLK(n1640), .Q(\mem0[167][5] ), .QN(n24259) );
  SDFFX1 \mem0_reg[167][4]  ( .D(n17896), .SI(\mem0[167][3] ), .SE(test_se), 
        .CLK(n1640), .Q(\mem0[167][4] ), .QN(n24260) );
  SDFFX1 \mem0_reg[167][3]  ( .D(n17895), .SI(\mem0[167][2] ), .SE(test_se), 
        .CLK(n1640), .Q(\mem0[167][3] ), .QN(n24261) );
  SDFFX1 \mem0_reg[167][2]  ( .D(n17894), .SI(\mem0[167][1] ), .SE(test_se), 
        .CLK(n1640), .Q(\mem0[167][2] ), .QN(n24262) );
  SDFFX1 \mem0_reg[167][1]  ( .D(n17893), .SI(\mem0[167][0] ), .SE(test_se), 
        .CLK(n1640), .Q(\mem0[167][1] ), .QN(n24263) );
  SDFFX1 \mem0_reg[167][0]  ( .D(n17892), .SI(\mem0[166][7] ), .SE(test_se), 
        .CLK(n1640), .Q(\mem0[167][0] ), .QN(n24264) );
  SDFFX1 \mem0_reg[166][7]  ( .D(n17891), .SI(\mem0[166][6] ), .SE(test_se), 
        .CLK(n1640), .Q(\mem0[166][7] ), .QN(n24265) );
  SDFFX1 \mem0_reg[166][6]  ( .D(n17890), .SI(\mem0[166][5] ), .SE(test_se), 
        .CLK(n1640), .Q(\mem0[166][6] ), .QN(n24266) );
  SDFFX1 \mem0_reg[166][5]  ( .D(n17889), .SI(\mem0[166][4] ), .SE(test_se), 
        .CLK(n1640), .Q(\mem0[166][5] ), .QN(n24267) );
  SDFFX1 \mem0_reg[166][4]  ( .D(n17888), .SI(\mem0[166][3] ), .SE(test_se), 
        .CLK(n1640), .Q(\mem0[166][4] ), .QN(n24268) );
  SDFFX1 \mem0_reg[166][3]  ( .D(n17887), .SI(\mem0[166][2] ), .SE(test_se), 
        .CLK(n1640), .Q(\mem0[166][3] ), .QN(n24269) );
  SDFFX1 \mem0_reg[166][2]  ( .D(n17886), .SI(\mem0[166][1] ), .SE(test_se), 
        .CLK(n1640), .Q(\mem0[166][2] ), .QN(n24270) );
  SDFFX1 \mem0_reg[166][1]  ( .D(n17885), .SI(\mem0[166][0] ), .SE(test_se), 
        .CLK(n1641), .Q(\mem0[166][1] ), .QN(n24271) );
  SDFFX1 \mem0_reg[166][0]  ( .D(n17884), .SI(\mem0[165][7] ), .SE(test_se), 
        .CLK(n1641), .Q(\mem0[166][0] ), .QN(n24272) );
  SDFFX1 \mem0_reg[165][7]  ( .D(n17883), .SI(\mem0[165][6] ), .SE(test_se), 
        .CLK(n1641), .Q(\mem0[165][7] ), .QN(n24273) );
  SDFFX1 \mem0_reg[165][6]  ( .D(n17882), .SI(\mem0[165][5] ), .SE(test_se), 
        .CLK(n1641), .Q(\mem0[165][6] ), .QN(n24274) );
  SDFFX1 \mem0_reg[165][5]  ( .D(n17881), .SI(\mem0[165][4] ), .SE(test_se), 
        .CLK(n1641), .Q(\mem0[165][5] ), .QN(n24275) );
  SDFFX1 \mem0_reg[165][4]  ( .D(n17880), .SI(\mem0[165][3] ), .SE(test_se), 
        .CLK(n1641), .Q(\mem0[165][4] ), .QN(n24276) );
  SDFFX1 \mem0_reg[165][3]  ( .D(n17879), .SI(\mem0[165][2] ), .SE(test_se), 
        .CLK(n1641), .Q(\mem0[165][3] ), .QN(n24277) );
  SDFFX1 \mem0_reg[165][2]  ( .D(n17878), .SI(\mem0[165][1] ), .SE(test_se), 
        .CLK(n1641), .Q(\mem0[165][2] ), .QN(n24278) );
  SDFFX1 \mem0_reg[165][1]  ( .D(n17877), .SI(\mem0[165][0] ), .SE(test_se), 
        .CLK(n1641), .Q(\mem0[165][1] ), .QN(n24279) );
  SDFFX1 \mem0_reg[165][0]  ( .D(n17876), .SI(\mem0[164][7] ), .SE(test_se), 
        .CLK(n1641), .Q(\mem0[165][0] ), .QN(n24280) );
  SDFFX1 \mem0_reg[164][7]  ( .D(n17875), .SI(\mem0[164][6] ), .SE(test_se), 
        .CLK(n1641), .Q(\mem0[164][7] ), .QN(n24281) );
  SDFFX1 \mem0_reg[164][6]  ( .D(n17874), .SI(\mem0[164][5] ), .SE(test_se), 
        .CLK(n1641), .Q(\mem0[164][6] ), .QN(n24282) );
  SDFFX1 \mem0_reg[164][5]  ( .D(n17873), .SI(\mem0[164][4] ), .SE(test_se), 
        .CLK(n1642), .Q(\mem0[164][5] ), .QN(n24283) );
  SDFFX1 \mem0_reg[164][4]  ( .D(n17872), .SI(\mem0[164][3] ), .SE(test_se), 
        .CLK(n1642), .Q(\mem0[164][4] ), .QN(n24284) );
  SDFFX1 \mem0_reg[164][3]  ( .D(n17871), .SI(\mem0[164][2] ), .SE(test_se), 
        .CLK(n1642), .Q(\mem0[164][3] ), .QN(n24285) );
  SDFFX1 \mem0_reg[164][2]  ( .D(n17870), .SI(\mem0[164][1] ), .SE(test_se), 
        .CLK(n1642), .Q(\mem0[164][2] ), .QN(n24286) );
  SDFFX1 \mem0_reg[164][1]  ( .D(n17869), .SI(\mem0[164][0] ), .SE(test_se), 
        .CLK(n1642), .Q(\mem0[164][1] ), .QN(n24287) );
  SDFFX1 \mem0_reg[164][0]  ( .D(n17868), .SI(\mem0[163][7] ), .SE(test_se), 
        .CLK(n1642), .Q(\mem0[164][0] ), .QN(n24288) );
  SDFFX1 \mem0_reg[163][7]  ( .D(n17867), .SI(\mem0[163][6] ), .SE(test_se), 
        .CLK(n1642), .Q(\mem0[163][7] ), .QN(n24289) );
  SDFFX1 \mem0_reg[163][6]  ( .D(n17866), .SI(\mem0[163][5] ), .SE(test_se), 
        .CLK(n1642), .Q(\mem0[163][6] ), .QN(n24290) );
  SDFFX1 \mem0_reg[163][5]  ( .D(n17865), .SI(\mem0[163][4] ), .SE(test_se), 
        .CLK(n1642), .Q(\mem0[163][5] ), .QN(n24291) );
  SDFFX1 \mem0_reg[163][4]  ( .D(n17864), .SI(\mem0[163][3] ), .SE(test_se), 
        .CLK(n1642), .Q(\mem0[163][4] ), .QN(n24292) );
  SDFFX1 \mem0_reg[163][3]  ( .D(n17863), .SI(\mem0[163][2] ), .SE(test_se), 
        .CLK(n1642), .Q(\mem0[163][3] ), .QN(n24293) );
  SDFFX1 \mem0_reg[163][2]  ( .D(n17862), .SI(\mem0[163][1] ), .SE(test_se), 
        .CLK(n1642), .Q(\mem0[163][2] ), .QN(n24294) );
  SDFFX1 \mem0_reg[163][1]  ( .D(n17861), .SI(\mem0[163][0] ), .SE(test_se), 
        .CLK(n1643), .Q(\mem0[163][1] ), .QN(n24295) );
  SDFFX1 \mem0_reg[163][0]  ( .D(n17860), .SI(\mem0[162][7] ), .SE(test_se), 
        .CLK(n1643), .Q(\mem0[163][0] ), .QN(n24296) );
  SDFFX1 \mem0_reg[162][7]  ( .D(n17859), .SI(\mem0[162][6] ), .SE(test_se), 
        .CLK(n1643), .Q(\mem0[162][7] ), .QN(n24297) );
  SDFFX1 \mem0_reg[162][6]  ( .D(n17858), .SI(\mem0[162][5] ), .SE(test_se), 
        .CLK(n1643), .Q(\mem0[162][6] ), .QN(n24298) );
  SDFFX1 \mem0_reg[162][5]  ( .D(n17857), .SI(\mem0[162][4] ), .SE(test_se), 
        .CLK(n1643), .Q(\mem0[162][5] ), .QN(n24299) );
  SDFFX1 \mem0_reg[162][4]  ( .D(n17856), .SI(\mem0[162][3] ), .SE(test_se), 
        .CLK(n1643), .Q(\mem0[162][4] ), .QN(n24300) );
  SDFFX1 \mem0_reg[162][3]  ( .D(n17855), .SI(\mem0[162][2] ), .SE(test_se), 
        .CLK(n1643), .Q(\mem0[162][3] ), .QN(n24301) );
  SDFFX1 \mem0_reg[162][2]  ( .D(n17854), .SI(\mem0[162][1] ), .SE(test_se), 
        .CLK(n1643), .Q(\mem0[162][2] ), .QN(n24302) );
  SDFFX1 \mem0_reg[162][1]  ( .D(n17853), .SI(\mem0[162][0] ), .SE(test_se), 
        .CLK(n1643), .Q(\mem0[162][1] ), .QN(n24303) );
  SDFFX1 \mem0_reg[162][0]  ( .D(n17852), .SI(\mem0[161][7] ), .SE(test_se), 
        .CLK(n1643), .Q(\mem0[162][0] ), .QN(n24304) );
  SDFFX1 \mem0_reg[161][7]  ( .D(n17851), .SI(\mem0[161][6] ), .SE(test_se), 
        .CLK(n1643), .Q(\mem0[161][7] ), .QN(n24305) );
  SDFFX1 \mem0_reg[161][6]  ( .D(n17850), .SI(\mem0[161][5] ), .SE(test_se), 
        .CLK(n1643), .Q(\mem0[161][6] ), .QN(n24306) );
  SDFFX1 \mem0_reg[161][5]  ( .D(n17849), .SI(\mem0[161][4] ), .SE(test_se), 
        .CLK(n1644), .Q(\mem0[161][5] ), .QN(n24307) );
  SDFFX1 \mem0_reg[161][4]  ( .D(n17848), .SI(\mem0[161][3] ), .SE(test_se), 
        .CLK(n1644), .Q(\mem0[161][4] ), .QN(n24308) );
  SDFFX1 \mem0_reg[161][3]  ( .D(n17847), .SI(\mem0[161][2] ), .SE(test_se), 
        .CLK(n1644), .Q(\mem0[161][3] ), .QN(n24309) );
  SDFFX1 \mem0_reg[161][2]  ( .D(n17846), .SI(\mem0[161][1] ), .SE(test_se), 
        .CLK(n1644), .Q(\mem0[161][2] ), .QN(n24310) );
  SDFFX1 \mem0_reg[161][1]  ( .D(n17845), .SI(\mem0[161][0] ), .SE(test_se), 
        .CLK(n1644), .Q(\mem0[161][1] ), .QN(n24311) );
  SDFFX1 \mem0_reg[161][0]  ( .D(n17844), .SI(\mem0[160][7] ), .SE(test_se), 
        .CLK(n1644), .Q(\mem0[161][0] ), .QN(n24312) );
  SDFFX1 \mem0_reg[160][7]  ( .D(n17843), .SI(\mem0[160][6] ), .SE(test_se), 
        .CLK(n1644), .Q(\mem0[160][7] ), .QN(n24313) );
  SDFFX1 \mem0_reg[160][6]  ( .D(n17842), .SI(\mem0[160][5] ), .SE(test_se), 
        .CLK(n1644), .Q(\mem0[160][6] ), .QN(n24314) );
  SDFFX1 \mem0_reg[160][5]  ( .D(n17841), .SI(\mem0[160][4] ), .SE(test_se), 
        .CLK(n1644), .Q(\mem0[160][5] ), .QN(n24315) );
  SDFFX1 \mem0_reg[160][4]  ( .D(n17840), .SI(\mem0[160][3] ), .SE(test_se), 
        .CLK(n1644), .Q(\mem0[160][4] ), .QN(n24316) );
  SDFFX1 \mem0_reg[160][3]  ( .D(n17839), .SI(\mem0[160][2] ), .SE(test_se), 
        .CLK(n1644), .Q(\mem0[160][3] ), .QN(n24317) );
  SDFFX1 \mem0_reg[160][2]  ( .D(n17838), .SI(\mem0[160][1] ), .SE(test_se), 
        .CLK(n1644), .Q(\mem0[160][2] ), .QN(n24318) );
  SDFFX1 \mem0_reg[160][1]  ( .D(n17837), .SI(\mem0[160][0] ), .SE(test_se), 
        .CLK(n1645), .Q(\mem0[160][1] ), .QN(n24319) );
  SDFFX1 \mem0_reg[160][0]  ( .D(n17836), .SI(\mem0[159][7] ), .SE(test_se), 
        .CLK(n1645), .Q(\mem0[160][0] ), .QN(n24320) );
  SDFFX1 \mem0_reg[159][7]  ( .D(n17835), .SI(\mem0[159][6] ), .SE(test_se), 
        .CLK(n1645), .Q(\mem0[159][7] ), .QN(n24321) );
  SDFFX1 \mem0_reg[159][6]  ( .D(n17834), .SI(\mem0[159][5] ), .SE(test_se), 
        .CLK(n1645), .Q(\mem0[159][6] ), .QN(n24322) );
  SDFFX1 \mem0_reg[159][5]  ( .D(n17833), .SI(\mem0[159][4] ), .SE(test_se), 
        .CLK(n1645), .Q(\mem0[159][5] ), .QN(n24323) );
  SDFFX1 \mem0_reg[159][4]  ( .D(n17832), .SI(\mem0[159][3] ), .SE(test_se), 
        .CLK(n1645), .Q(\mem0[159][4] ), .QN(n24324) );
  SDFFX1 \mem0_reg[159][3]  ( .D(n17831), .SI(\mem0[159][2] ), .SE(test_se), 
        .CLK(n1645), .Q(\mem0[159][3] ), .QN(n24325) );
  SDFFX1 \mem0_reg[159][2]  ( .D(n17830), .SI(\mem0[159][1] ), .SE(test_se), 
        .CLK(n1645), .Q(\mem0[159][2] ), .QN(n24326) );
  SDFFX1 \mem0_reg[159][1]  ( .D(n17829), .SI(\mem0[159][0] ), .SE(test_se), 
        .CLK(n1645), .Q(\mem0[159][1] ), .QN(n24327) );
  SDFFX1 \mem0_reg[159][0]  ( .D(n17828), .SI(\mem0[158][7] ), .SE(test_se), 
        .CLK(n1645), .Q(\mem0[159][0] ), .QN(n24328) );
  SDFFX1 \mem0_reg[158][7]  ( .D(n17827), .SI(\mem0[158][6] ), .SE(test_se), 
        .CLK(n1645), .Q(\mem0[158][7] ), .QN(n24329) );
  SDFFX1 \mem0_reg[158][6]  ( .D(n17826), .SI(\mem0[158][5] ), .SE(test_se), 
        .CLK(n1645), .Q(\mem0[158][6] ), .QN(n24330) );
  SDFFX1 \mem0_reg[158][5]  ( .D(n17825), .SI(\mem0[158][4] ), .SE(test_se), 
        .CLK(n1646), .Q(\mem0[158][5] ), .QN(n24331) );
  SDFFX1 \mem0_reg[158][4]  ( .D(n17824), .SI(\mem0[158][3] ), .SE(test_se), 
        .CLK(n1646), .Q(\mem0[158][4] ), .QN(n24332) );
  SDFFX1 \mem0_reg[158][3]  ( .D(n17823), .SI(\mem0[158][2] ), .SE(test_se), 
        .CLK(n1646), .Q(\mem0[158][3] ), .QN(n24333) );
  SDFFX1 \mem0_reg[158][2]  ( .D(n17822), .SI(\mem0[158][1] ), .SE(test_se), 
        .CLK(n1646), .Q(\mem0[158][2] ), .QN(n24334) );
  SDFFX1 \mem0_reg[158][1]  ( .D(n17821), .SI(\mem0[158][0] ), .SE(test_se), 
        .CLK(n1646), .Q(\mem0[158][1] ), .QN(n24335) );
  SDFFX1 \mem0_reg[158][0]  ( .D(n17820), .SI(\mem0[157][7] ), .SE(test_se), 
        .CLK(n1646), .Q(\mem0[158][0] ), .QN(n24336) );
  SDFFX1 \mem0_reg[157][7]  ( .D(n17819), .SI(\mem0[157][6] ), .SE(test_se), 
        .CLK(n1646), .Q(\mem0[157][7] ), .QN(n24337) );
  SDFFX1 \mem0_reg[157][6]  ( .D(n17818), .SI(\mem0[157][5] ), .SE(test_se), 
        .CLK(n1646), .Q(\mem0[157][6] ), .QN(n24338) );
  SDFFX1 \mem0_reg[157][5]  ( .D(n17817), .SI(\mem0[157][4] ), .SE(test_se), 
        .CLK(n1646), .Q(\mem0[157][5] ), .QN(n24339) );
  SDFFX1 \mem0_reg[157][4]  ( .D(n17816), .SI(\mem0[157][3] ), .SE(test_se), 
        .CLK(n1646), .Q(\mem0[157][4] ), .QN(n24340) );
  SDFFX1 \mem0_reg[157][3]  ( .D(n17815), .SI(\mem0[157][2] ), .SE(test_se), 
        .CLK(n1646), .Q(\mem0[157][3] ), .QN(n24341) );
  SDFFX1 \mem0_reg[157][2]  ( .D(n17814), .SI(\mem0[157][1] ), .SE(test_se), 
        .CLK(n1646), .Q(\mem0[157][2] ), .QN(n24342) );
  SDFFX1 \mem0_reg[157][1]  ( .D(n17813), .SI(\mem0[157][0] ), .SE(test_se), 
        .CLK(n1647), .Q(\mem0[157][1] ), .QN(n24343) );
  SDFFX1 \mem0_reg[157][0]  ( .D(n17812), .SI(\mem0[156][7] ), .SE(test_se), 
        .CLK(n1647), .Q(\mem0[157][0] ), .QN(n24344) );
  SDFFX1 \mem0_reg[156][7]  ( .D(n17811), .SI(\mem0[156][6] ), .SE(test_se), 
        .CLK(n1647), .Q(\mem0[156][7] ), .QN(n24345) );
  SDFFX1 \mem0_reg[156][6]  ( .D(n17810), .SI(\mem0[156][5] ), .SE(test_se), 
        .CLK(n1647), .Q(\mem0[156][6] ), .QN(n24346) );
  SDFFX1 \mem0_reg[156][5]  ( .D(n17809), .SI(\mem0[156][4] ), .SE(test_se), 
        .CLK(n1647), .Q(\mem0[156][5] ), .QN(n24347) );
  SDFFX1 \mem0_reg[156][4]  ( .D(n17808), .SI(\mem0[156][3] ), .SE(test_se), 
        .CLK(n1647), .Q(\mem0[156][4] ), .QN(n24348) );
  SDFFX1 \mem0_reg[156][3]  ( .D(n17807), .SI(\mem0[156][2] ), .SE(test_se), 
        .CLK(n1647), .Q(\mem0[156][3] ), .QN(n24349) );
  SDFFX1 \mem0_reg[156][2]  ( .D(n17806), .SI(\mem0[156][1] ), .SE(test_se), 
        .CLK(n1647), .Q(\mem0[156][2] ), .QN(n24350) );
  SDFFX1 \mem0_reg[156][1]  ( .D(n17805), .SI(\mem0[156][0] ), .SE(test_se), 
        .CLK(n1647), .Q(\mem0[156][1] ), .QN(n24351) );
  SDFFX1 \mem0_reg[156][0]  ( .D(n17804), .SI(\mem0[155][7] ), .SE(test_se), 
        .CLK(n1647), .Q(\mem0[156][0] ), .QN(n24352) );
  SDFFX1 \mem0_reg[155][7]  ( .D(n17803), .SI(\mem0[155][6] ), .SE(test_se), 
        .CLK(n1647), .Q(\mem0[155][7] ), .QN(n24353) );
  SDFFX1 \mem0_reg[155][6]  ( .D(n17802), .SI(\mem0[155][5] ), .SE(test_se), 
        .CLK(n1647), .Q(\mem0[155][6] ), .QN(n24354) );
  SDFFX1 \mem0_reg[155][5]  ( .D(n17801), .SI(\mem0[155][4] ), .SE(test_se), 
        .CLK(n1648), .Q(\mem0[155][5] ), .QN(n24355) );
  SDFFX1 \mem0_reg[155][4]  ( .D(n17800), .SI(\mem0[155][3] ), .SE(test_se), 
        .CLK(n1648), .Q(\mem0[155][4] ), .QN(n24356) );
  SDFFX1 \mem0_reg[155][3]  ( .D(n17799), .SI(\mem0[155][2] ), .SE(test_se), 
        .CLK(n1648), .Q(\mem0[155][3] ), .QN(n24357) );
  SDFFX1 \mem0_reg[155][2]  ( .D(n17798), .SI(\mem0[155][1] ), .SE(test_se), 
        .CLK(n1648), .Q(\mem0[155][2] ), .QN(n24358) );
  SDFFX1 \mem0_reg[155][1]  ( .D(n17797), .SI(\mem0[155][0] ), .SE(test_se), 
        .CLK(n1648), .Q(\mem0[155][1] ), .QN(n24359) );
  SDFFX1 \mem0_reg[155][0]  ( .D(n17796), .SI(\mem0[154][7] ), .SE(test_se), 
        .CLK(n1648), .Q(\mem0[155][0] ), .QN(n24360) );
  SDFFX1 \mem0_reg[154][7]  ( .D(n17795), .SI(\mem0[154][6] ), .SE(test_se), 
        .CLK(n1648), .Q(\mem0[154][7] ), .QN(n24361) );
  SDFFX1 \mem0_reg[154][6]  ( .D(n17794), .SI(\mem0[154][5] ), .SE(test_se), 
        .CLK(n1648), .Q(\mem0[154][6] ), .QN(n24362) );
  SDFFX1 \mem0_reg[154][5]  ( .D(n17793), .SI(\mem0[154][4] ), .SE(test_se), 
        .CLK(n1648), .Q(\mem0[154][5] ), .QN(n24363) );
  SDFFX1 \mem0_reg[154][4]  ( .D(n17792), .SI(\mem0[154][3] ), .SE(test_se), 
        .CLK(n1648), .Q(\mem0[154][4] ), .QN(n24364) );
  SDFFX1 \mem0_reg[154][3]  ( .D(n17791), .SI(\mem0[154][2] ), .SE(test_se), 
        .CLK(n1648), .Q(\mem0[154][3] ), .QN(n24365) );
  SDFFX1 \mem0_reg[154][2]  ( .D(n17790), .SI(\mem0[154][1] ), .SE(test_se), 
        .CLK(n1648), .Q(\mem0[154][2] ), .QN(n24366) );
  SDFFX1 \mem0_reg[154][1]  ( .D(n17789), .SI(\mem0[154][0] ), .SE(test_se), 
        .CLK(n1649), .Q(\mem0[154][1] ), .QN(n24367) );
  SDFFX1 \mem0_reg[154][0]  ( .D(n17788), .SI(\mem0[153][7] ), .SE(test_se), 
        .CLK(n1649), .Q(\mem0[154][0] ), .QN(n24368) );
  SDFFX1 \mem0_reg[153][7]  ( .D(n17787), .SI(\mem0[153][6] ), .SE(test_se), 
        .CLK(n1649), .Q(\mem0[153][7] ), .QN(n24369) );
  SDFFX1 \mem0_reg[153][6]  ( .D(n17786), .SI(\mem0[153][5] ), .SE(test_se), 
        .CLK(n1649), .Q(\mem0[153][6] ), .QN(n24370) );
  SDFFX1 \mem0_reg[153][5]  ( .D(n17785), .SI(\mem0[153][4] ), .SE(test_se), 
        .CLK(n1649), .Q(\mem0[153][5] ), .QN(n24371) );
  SDFFX1 \mem0_reg[153][4]  ( .D(n17784), .SI(\mem0[153][3] ), .SE(test_se), 
        .CLK(n1649), .Q(\mem0[153][4] ), .QN(n24372) );
  SDFFX1 \mem0_reg[153][3]  ( .D(n17783), .SI(\mem0[153][2] ), .SE(test_se), 
        .CLK(n1649), .Q(\mem0[153][3] ), .QN(n24373) );
  SDFFX1 \mem0_reg[153][2]  ( .D(n17782), .SI(\mem0[153][1] ), .SE(test_se), 
        .CLK(n1649), .Q(\mem0[153][2] ), .QN(n24374) );
  SDFFX1 \mem0_reg[153][1]  ( .D(n17781), .SI(\mem0[153][0] ), .SE(test_se), 
        .CLK(n1649), .Q(\mem0[153][1] ), .QN(n24375) );
  SDFFX1 \mem0_reg[153][0]  ( .D(n17780), .SI(\mem0[152][7] ), .SE(test_se), 
        .CLK(n1649), .Q(\mem0[153][0] ), .QN(n24376) );
  SDFFX1 \mem0_reg[152][7]  ( .D(n17779), .SI(\mem0[152][6] ), .SE(test_se), 
        .CLK(n1649), .Q(\mem0[152][7] ), .QN(n24377) );
  SDFFX1 \mem0_reg[152][6]  ( .D(n17778), .SI(\mem0[152][5] ), .SE(test_se), 
        .CLK(n1649), .Q(\mem0[152][6] ), .QN(n24378) );
  SDFFX1 \mem0_reg[152][5]  ( .D(n17777), .SI(\mem0[152][4] ), .SE(test_se), 
        .CLK(n1650), .Q(\mem0[152][5] ), .QN(n24379) );
  SDFFX1 \mem0_reg[152][4]  ( .D(n17776), .SI(\mem0[152][3] ), .SE(test_se), 
        .CLK(n1650), .Q(\mem0[152][4] ), .QN(n24380) );
  SDFFX1 \mem0_reg[152][3]  ( .D(n17775), .SI(\mem0[152][2] ), .SE(test_se), 
        .CLK(n1650), .Q(\mem0[152][3] ), .QN(n24381) );
  SDFFX1 \mem0_reg[152][2]  ( .D(n17774), .SI(\mem0[152][1] ), .SE(test_se), 
        .CLK(n1650), .Q(\mem0[152][2] ), .QN(n24382) );
  SDFFX1 \mem0_reg[152][1]  ( .D(n17773), .SI(\mem0[152][0] ), .SE(test_se), 
        .CLK(n1650), .Q(\mem0[152][1] ), .QN(n24383) );
  SDFFX1 \mem0_reg[152][0]  ( .D(n17772), .SI(\mem0[151][7] ), .SE(test_se), 
        .CLK(n1650), .Q(\mem0[152][0] ), .QN(n24384) );
  SDFFX1 \mem0_reg[151][7]  ( .D(n17771), .SI(\mem0[151][6] ), .SE(test_se), 
        .CLK(n1650), .Q(\mem0[151][7] ), .QN(n24385) );
  SDFFX1 \mem0_reg[151][6]  ( .D(n17770), .SI(\mem0[151][5] ), .SE(test_se), 
        .CLK(n1650), .Q(\mem0[151][6] ), .QN(n24386) );
  SDFFX1 \mem0_reg[151][5]  ( .D(n17769), .SI(\mem0[151][4] ), .SE(test_se), 
        .CLK(n1650), .Q(\mem0[151][5] ), .QN(n24387) );
  SDFFX1 \mem0_reg[151][4]  ( .D(n17768), .SI(\mem0[151][3] ), .SE(test_se), 
        .CLK(n1650), .Q(\mem0[151][4] ), .QN(n24388) );
  SDFFX1 \mem0_reg[151][3]  ( .D(n17767), .SI(\mem0[151][2] ), .SE(test_se), 
        .CLK(n1650), .Q(\mem0[151][3] ), .QN(n24389) );
  SDFFX1 \mem0_reg[151][2]  ( .D(n17766), .SI(\mem0[151][1] ), .SE(test_se), 
        .CLK(n1650), .Q(\mem0[151][2] ), .QN(n24390) );
  SDFFX1 \mem0_reg[151][1]  ( .D(n17765), .SI(\mem0[151][0] ), .SE(test_se), 
        .CLK(n1651), .Q(\mem0[151][1] ), .QN(n24391) );
  SDFFX1 \mem0_reg[151][0]  ( .D(n17764), .SI(\mem0[150][7] ), .SE(test_se), 
        .CLK(n1651), .Q(\mem0[151][0] ), .QN(n24392) );
  SDFFX1 \mem0_reg[150][7]  ( .D(n17763), .SI(\mem0[150][6] ), .SE(test_se), 
        .CLK(n1651), .Q(\mem0[150][7] ), .QN(n24393) );
  SDFFX1 \mem0_reg[150][6]  ( .D(n17762), .SI(\mem0[150][5] ), .SE(test_se), 
        .CLK(n1651), .Q(\mem0[150][6] ), .QN(n24394) );
  SDFFX1 \mem0_reg[150][5]  ( .D(n17761), .SI(\mem0[150][4] ), .SE(test_se), 
        .CLK(n1651), .Q(\mem0[150][5] ), .QN(n24395) );
  SDFFX1 \mem0_reg[150][4]  ( .D(n17760), .SI(\mem0[150][3] ), .SE(test_se), 
        .CLK(n1651), .Q(\mem0[150][4] ), .QN(n24396) );
  SDFFX1 \mem0_reg[150][3]  ( .D(n17759), .SI(\mem0[150][2] ), .SE(test_se), 
        .CLK(n1651), .Q(\mem0[150][3] ), .QN(n24397) );
  SDFFX1 \mem0_reg[150][2]  ( .D(n17758), .SI(\mem0[150][1] ), .SE(test_se), 
        .CLK(n1651), .Q(\mem0[150][2] ), .QN(n24398) );
  SDFFX1 \mem0_reg[150][1]  ( .D(n17757), .SI(\mem0[150][0] ), .SE(test_se), 
        .CLK(n1651), .Q(\mem0[150][1] ), .QN(n24399) );
  SDFFX1 \mem0_reg[150][0]  ( .D(n17756), .SI(\mem0[149][7] ), .SE(test_se), 
        .CLK(n1651), .Q(\mem0[150][0] ), .QN(n24400) );
  SDFFX1 \mem0_reg[149][7]  ( .D(n17755), .SI(\mem0[149][6] ), .SE(test_se), 
        .CLK(n1651), .Q(\mem0[149][7] ), .QN(n24401) );
  SDFFX1 \mem0_reg[149][6]  ( .D(n17754), .SI(\mem0[149][5] ), .SE(test_se), 
        .CLK(n1651), .Q(\mem0[149][6] ), .QN(n24402) );
  SDFFX1 \mem0_reg[149][5]  ( .D(n17753), .SI(\mem0[149][4] ), .SE(test_se), 
        .CLK(n1652), .Q(\mem0[149][5] ), .QN(n24403) );
  SDFFX1 \mem0_reg[149][4]  ( .D(n17752), .SI(\mem0[149][3] ), .SE(test_se), 
        .CLK(n1652), .Q(\mem0[149][4] ), .QN(n24404) );
  SDFFX1 \mem0_reg[149][3]  ( .D(n17751), .SI(\mem0[149][2] ), .SE(test_se), 
        .CLK(n1652), .Q(\mem0[149][3] ), .QN(n24405) );
  SDFFX1 \mem0_reg[149][2]  ( .D(n17750), .SI(\mem0[149][1] ), .SE(test_se), 
        .CLK(n1652), .Q(\mem0[149][2] ), .QN(n24406) );
  SDFFX1 \mem0_reg[149][1]  ( .D(n17749), .SI(\mem0[149][0] ), .SE(test_se), 
        .CLK(n1652), .Q(\mem0[149][1] ), .QN(n24407) );
  SDFFX1 \mem0_reg[149][0]  ( .D(n17748), .SI(\mem0[148][7] ), .SE(test_se), 
        .CLK(n1652), .Q(\mem0[149][0] ), .QN(n24408) );
  SDFFX1 \mem0_reg[148][7]  ( .D(n17747), .SI(\mem0[148][6] ), .SE(test_se), 
        .CLK(n1652), .Q(\mem0[148][7] ), .QN(n24409) );
  SDFFX1 \mem0_reg[148][6]  ( .D(n17746), .SI(\mem0[148][5] ), .SE(test_se), 
        .CLK(n1652), .Q(\mem0[148][6] ), .QN(n24410) );
  SDFFX1 \mem0_reg[148][5]  ( .D(n17745), .SI(\mem0[148][4] ), .SE(test_se), 
        .CLK(n1652), .Q(\mem0[148][5] ), .QN(n24411) );
  SDFFX1 \mem0_reg[148][4]  ( .D(n17744), .SI(\mem0[148][3] ), .SE(test_se), 
        .CLK(n1652), .Q(\mem0[148][4] ), .QN(n24412) );
  SDFFX1 \mem0_reg[148][3]  ( .D(n17743), .SI(\mem0[148][2] ), .SE(test_se), 
        .CLK(n1652), .Q(\mem0[148][3] ), .QN(n24413) );
  SDFFX1 \mem0_reg[148][2]  ( .D(n17742), .SI(\mem0[148][1] ), .SE(test_se), 
        .CLK(n1652), .Q(\mem0[148][2] ), .QN(n24414) );
  SDFFX1 \mem0_reg[148][1]  ( .D(n17741), .SI(\mem0[148][0] ), .SE(test_se), 
        .CLK(n1653), .Q(\mem0[148][1] ), .QN(n24415) );
  SDFFX1 \mem0_reg[148][0]  ( .D(n17740), .SI(\mem0[147][7] ), .SE(test_se), 
        .CLK(n1653), .Q(\mem0[148][0] ), .QN(n24416) );
  SDFFX1 \mem0_reg[147][7]  ( .D(n17739), .SI(\mem0[147][6] ), .SE(test_se), 
        .CLK(n1653), .Q(\mem0[147][7] ), .QN(n24417) );
  SDFFX1 \mem0_reg[147][6]  ( .D(n17738), .SI(\mem0[147][5] ), .SE(test_se), 
        .CLK(n1653), .Q(\mem0[147][6] ), .QN(n24418) );
  SDFFX1 \mem0_reg[147][5]  ( .D(n17737), .SI(\mem0[147][4] ), .SE(test_se), 
        .CLK(n1653), .Q(\mem0[147][5] ), .QN(n24419) );
  SDFFX1 \mem0_reg[147][4]  ( .D(n17736), .SI(\mem0[147][3] ), .SE(test_se), 
        .CLK(n1653), .Q(\mem0[147][4] ), .QN(n24420) );
  SDFFX1 \mem0_reg[147][3]  ( .D(n17735), .SI(\mem0[147][2] ), .SE(test_se), 
        .CLK(n1653), .Q(\mem0[147][3] ), .QN(n24421) );
  SDFFX1 \mem0_reg[147][2]  ( .D(n17734), .SI(\mem0[147][1] ), .SE(test_se), 
        .CLK(n1653), .Q(\mem0[147][2] ), .QN(n24422) );
  SDFFX1 \mem0_reg[147][1]  ( .D(n17733), .SI(\mem0[147][0] ), .SE(test_se), 
        .CLK(n1653), .Q(\mem0[147][1] ), .QN(n24423) );
  SDFFX1 \mem0_reg[147][0]  ( .D(n17732), .SI(\mem0[146][7] ), .SE(test_se), 
        .CLK(n1653), .Q(\mem0[147][0] ), .QN(n24424) );
  SDFFX1 \mem0_reg[146][7]  ( .D(n17731), .SI(\mem0[146][6] ), .SE(test_se), 
        .CLK(n1653), .Q(\mem0[146][7] ), .QN(n24425) );
  SDFFX1 \mem0_reg[146][6]  ( .D(n17730), .SI(\mem0[146][5] ), .SE(test_se), 
        .CLK(n1653), .Q(\mem0[146][6] ), .QN(n24426) );
  SDFFX1 \mem0_reg[146][5]  ( .D(n17729), .SI(\mem0[146][4] ), .SE(test_se), 
        .CLK(n1654), .Q(\mem0[146][5] ), .QN(n24427) );
  SDFFX1 \mem0_reg[146][4]  ( .D(n17728), .SI(\mem0[146][3] ), .SE(test_se), 
        .CLK(n1654), .Q(\mem0[146][4] ), .QN(n24428) );
  SDFFX1 \mem0_reg[146][3]  ( .D(n17727), .SI(\mem0[146][2] ), .SE(test_se), 
        .CLK(n1654), .Q(\mem0[146][3] ), .QN(n24429) );
  SDFFX1 \mem0_reg[146][2]  ( .D(n17726), .SI(\mem0[146][1] ), .SE(test_se), 
        .CLK(n1654), .Q(\mem0[146][2] ), .QN(n24430) );
  SDFFX1 \mem0_reg[146][1]  ( .D(n17725), .SI(\mem0[146][0] ), .SE(test_se), 
        .CLK(n1654), .Q(\mem0[146][1] ), .QN(n24431) );
  SDFFX1 \mem0_reg[146][0]  ( .D(n17724), .SI(\mem0[145][7] ), .SE(test_se), 
        .CLK(n1654), .Q(\mem0[146][0] ), .QN(n24432) );
  SDFFX1 \mem0_reg[145][7]  ( .D(n17723), .SI(\mem0[145][6] ), .SE(test_se), 
        .CLK(n1654), .Q(\mem0[145][7] ), .QN(n24433) );
  SDFFX1 \mem0_reg[145][6]  ( .D(n17722), .SI(\mem0[145][5] ), .SE(test_se), 
        .CLK(n1654), .Q(\mem0[145][6] ), .QN(n24434) );
  SDFFX1 \mem0_reg[145][5]  ( .D(n17721), .SI(\mem0[145][4] ), .SE(test_se), 
        .CLK(n1654), .Q(\mem0[145][5] ), .QN(n24435) );
  SDFFX1 \mem0_reg[145][4]  ( .D(n17720), .SI(\mem0[145][3] ), .SE(test_se), 
        .CLK(n1654), .Q(\mem0[145][4] ), .QN(n24436) );
  SDFFX1 \mem0_reg[145][3]  ( .D(n17719), .SI(\mem0[145][2] ), .SE(test_se), 
        .CLK(n1654), .Q(\mem0[145][3] ), .QN(n24437) );
  SDFFX1 \mem0_reg[145][2]  ( .D(n17718), .SI(\mem0[145][1] ), .SE(test_se), 
        .CLK(n1654), .Q(\mem0[145][2] ), .QN(n24438) );
  SDFFX1 \mem0_reg[145][1]  ( .D(n17717), .SI(\mem0[145][0] ), .SE(test_se), 
        .CLK(n1655), .Q(\mem0[145][1] ), .QN(n24439) );
  SDFFX1 \mem0_reg[145][0]  ( .D(n17716), .SI(\mem0[144][7] ), .SE(test_se), 
        .CLK(n1655), .Q(\mem0[145][0] ), .QN(n24440) );
  SDFFX1 \mem0_reg[144][7]  ( .D(n17715), .SI(\mem0[144][6] ), .SE(test_se), 
        .CLK(n1655), .Q(\mem0[144][7] ), .QN(n24441) );
  SDFFX1 \mem0_reg[144][6]  ( .D(n17714), .SI(\mem0[144][5] ), .SE(test_se), 
        .CLK(n1655), .Q(\mem0[144][6] ), .QN(n24442) );
  SDFFX1 \mem0_reg[144][5]  ( .D(n17713), .SI(\mem0[144][4] ), .SE(test_se), 
        .CLK(n1655), .Q(\mem0[144][5] ), .QN(n24443) );
  SDFFX1 \mem0_reg[144][4]  ( .D(n17712), .SI(\mem0[144][3] ), .SE(test_se), 
        .CLK(n1655), .Q(\mem0[144][4] ), .QN(n24444) );
  SDFFX1 \mem0_reg[144][3]  ( .D(n17711), .SI(\mem0[144][2] ), .SE(test_se), 
        .CLK(n1655), .Q(\mem0[144][3] ), .QN(n24445) );
  SDFFX1 \mem0_reg[144][2]  ( .D(n17710), .SI(\mem0[144][1] ), .SE(test_se), 
        .CLK(n1655), .Q(\mem0[144][2] ), .QN(n24446) );
  SDFFX1 \mem0_reg[144][1]  ( .D(n17709), .SI(\mem0[144][0] ), .SE(test_se), 
        .CLK(n1655), .Q(\mem0[144][1] ), .QN(n24447) );
  SDFFX1 \mem0_reg[144][0]  ( .D(n17708), .SI(\mem0[143][7] ), .SE(test_se), 
        .CLK(n1655), .Q(\mem0[144][0] ), .QN(n24448) );
  SDFFX1 \mem0_reg[143][7]  ( .D(n17707), .SI(\mem0[143][6] ), .SE(test_se), 
        .CLK(n1655), .Q(\mem0[143][7] ), .QN(n24449) );
  SDFFX1 \mem0_reg[143][6]  ( .D(n17706), .SI(\mem0[143][5] ), .SE(test_se), 
        .CLK(n1655), .Q(\mem0[143][6] ), .QN(n24450) );
  SDFFX1 \mem0_reg[143][5]  ( .D(n17705), .SI(\mem0[143][4] ), .SE(test_se), 
        .CLK(n1656), .Q(\mem0[143][5] ), .QN(n24451) );
  SDFFX1 \mem0_reg[143][4]  ( .D(n17704), .SI(\mem0[143][3] ), .SE(test_se), 
        .CLK(n1656), .Q(\mem0[143][4] ), .QN(n24452) );
  SDFFX1 \mem0_reg[143][3]  ( .D(n17703), .SI(\mem0[143][2] ), .SE(test_se), 
        .CLK(n1656), .Q(\mem0[143][3] ), .QN(n24453) );
  SDFFX1 \mem0_reg[143][2]  ( .D(n17702), .SI(\mem0[143][1] ), .SE(test_se), 
        .CLK(n1656), .Q(\mem0[143][2] ), .QN(n24454) );
  SDFFX1 \mem0_reg[143][1]  ( .D(n17701), .SI(\mem0[143][0] ), .SE(test_se), 
        .CLK(n1656), .Q(\mem0[143][1] ), .QN(n24455) );
  SDFFX1 \mem0_reg[143][0]  ( .D(n17700), .SI(\mem0[142][7] ), .SE(test_se), 
        .CLK(n1656), .Q(\mem0[143][0] ), .QN(n24456) );
  SDFFX1 \mem0_reg[142][7]  ( .D(n17699), .SI(\mem0[142][6] ), .SE(test_se), 
        .CLK(n1656), .Q(\mem0[142][7] ), .QN(n24457) );
  SDFFX1 \mem0_reg[142][6]  ( .D(n17698), .SI(\mem0[142][5] ), .SE(test_se), 
        .CLK(n1656), .Q(\mem0[142][6] ), .QN(n24458) );
  SDFFX1 \mem0_reg[142][5]  ( .D(n17697), .SI(\mem0[142][4] ), .SE(test_se), 
        .CLK(n1656), .Q(\mem0[142][5] ), .QN(n24459) );
  SDFFX1 \mem0_reg[142][4]  ( .D(n17696), .SI(\mem0[142][3] ), .SE(test_se), 
        .CLK(n1656), .Q(\mem0[142][4] ), .QN(n24460) );
  SDFFX1 \mem0_reg[142][3]  ( .D(n17695), .SI(\mem0[142][2] ), .SE(test_se), 
        .CLK(n1656), .Q(\mem0[142][3] ), .QN(n24461) );
  SDFFX1 \mem0_reg[142][2]  ( .D(n17694), .SI(\mem0[142][1] ), .SE(test_se), 
        .CLK(n1656), .Q(\mem0[142][2] ), .QN(n24462) );
  SDFFX1 \mem0_reg[142][1]  ( .D(n17693), .SI(\mem0[142][0] ), .SE(test_se), 
        .CLK(n1657), .Q(\mem0[142][1] ), .QN(n24463) );
  SDFFX1 \mem0_reg[142][0]  ( .D(n17692), .SI(\mem0[141][7] ), .SE(test_se), 
        .CLK(n1657), .Q(\mem0[142][0] ), .QN(n24464) );
  SDFFX1 \mem0_reg[141][7]  ( .D(n17691), .SI(\mem0[141][6] ), .SE(test_se), 
        .CLK(n1657), .Q(\mem0[141][7] ), .QN(n24465) );
  SDFFX1 \mem0_reg[141][6]  ( .D(n17690), .SI(\mem0[141][5] ), .SE(test_se), 
        .CLK(n1657), .Q(\mem0[141][6] ), .QN(n24466) );
  SDFFX1 \mem0_reg[141][5]  ( .D(n17689), .SI(\mem0[141][4] ), .SE(test_se), 
        .CLK(n1657), .Q(\mem0[141][5] ), .QN(n24467) );
  SDFFX1 \mem0_reg[141][4]  ( .D(n17688), .SI(\mem0[141][3] ), .SE(test_se), 
        .CLK(n1657), .Q(\mem0[141][4] ), .QN(n24468) );
  SDFFX1 \mem0_reg[141][3]  ( .D(n17687), .SI(\mem0[141][2] ), .SE(test_se), 
        .CLK(n1657), .Q(\mem0[141][3] ), .QN(n24469) );
  SDFFX1 \mem0_reg[141][2]  ( .D(n17686), .SI(\mem0[141][1] ), .SE(test_se), 
        .CLK(n1657), .Q(\mem0[141][2] ), .QN(n24470) );
  SDFFX1 \mem0_reg[141][1]  ( .D(n17685), .SI(\mem0[141][0] ), .SE(test_se), 
        .CLK(n1657), .Q(\mem0[141][1] ), .QN(n24471) );
  SDFFX1 \mem0_reg[141][0]  ( .D(n17684), .SI(\mem0[140][7] ), .SE(test_se), 
        .CLK(n1657), .Q(\mem0[141][0] ), .QN(n24472) );
  SDFFX1 \mem0_reg[140][7]  ( .D(n17683), .SI(\mem0[140][6] ), .SE(test_se), 
        .CLK(n1657), .Q(\mem0[140][7] ), .QN(n24473) );
  SDFFX1 \mem0_reg[140][6]  ( .D(n17682), .SI(\mem0[140][5] ), .SE(test_se), 
        .CLK(n1657), .Q(\mem0[140][6] ), .QN(n24474) );
  SDFFX1 \mem0_reg[140][5]  ( .D(n17681), .SI(\mem0[140][4] ), .SE(test_se), 
        .CLK(n1658), .Q(\mem0[140][5] ), .QN(n24475) );
  SDFFX1 \mem0_reg[140][4]  ( .D(n17680), .SI(\mem0[140][3] ), .SE(test_se), 
        .CLK(n1658), .Q(\mem0[140][4] ), .QN(n24476) );
  SDFFX1 \mem0_reg[140][3]  ( .D(n17679), .SI(\mem0[140][2] ), .SE(test_se), 
        .CLK(n1658), .Q(\mem0[140][3] ), .QN(n24477) );
  SDFFX1 \mem0_reg[140][2]  ( .D(n17678), .SI(\mem0[140][1] ), .SE(test_se), 
        .CLK(n1658), .Q(\mem0[140][2] ), .QN(n24478) );
  SDFFX1 \mem0_reg[140][1]  ( .D(n17677), .SI(\mem0[140][0] ), .SE(test_se), 
        .CLK(n1658), .Q(\mem0[140][1] ), .QN(n24479) );
  SDFFX1 \mem0_reg[140][0]  ( .D(n17676), .SI(\mem0[139][7] ), .SE(test_se), 
        .CLK(n1658), .Q(\mem0[140][0] ), .QN(n24480) );
  SDFFX1 \mem0_reg[139][7]  ( .D(n17675), .SI(\mem0[139][6] ), .SE(test_se), 
        .CLK(n1658), .Q(\mem0[139][7] ), .QN(n24481) );
  SDFFX1 \mem0_reg[139][6]  ( .D(n17674), .SI(\mem0[139][5] ), .SE(test_se), 
        .CLK(n1658), .Q(\mem0[139][6] ), .QN(n24482) );
  SDFFX1 \mem0_reg[139][5]  ( .D(n17673), .SI(\mem0[139][4] ), .SE(test_se), 
        .CLK(n1658), .Q(\mem0[139][5] ), .QN(n24483) );
  SDFFX1 \mem0_reg[139][4]  ( .D(n17672), .SI(\mem0[139][3] ), .SE(test_se), 
        .CLK(n1658), .Q(\mem0[139][4] ), .QN(n24484) );
  SDFFX1 \mem0_reg[139][3]  ( .D(n17671), .SI(\mem0[139][2] ), .SE(test_se), 
        .CLK(n1658), .Q(\mem0[139][3] ), .QN(n24485) );
  SDFFX1 \mem0_reg[139][2]  ( .D(n17670), .SI(\mem0[139][1] ), .SE(test_se), 
        .CLK(n1658), .Q(\mem0[139][2] ), .QN(n24486) );
  SDFFX1 \mem0_reg[139][1]  ( .D(n17669), .SI(\mem0[139][0] ), .SE(test_se), 
        .CLK(n1659), .Q(\mem0[139][1] ), .QN(n24487) );
  SDFFX1 \mem0_reg[139][0]  ( .D(n17668), .SI(\mem0[138][7] ), .SE(test_se), 
        .CLK(n1659), .Q(\mem0[139][0] ), .QN(n24488) );
  SDFFX1 \mem0_reg[138][7]  ( .D(n17667), .SI(\mem0[138][6] ), .SE(test_se), 
        .CLK(n1659), .Q(\mem0[138][7] ), .QN(n24489) );
  SDFFX1 \mem0_reg[138][6]  ( .D(n17666), .SI(\mem0[138][5] ), .SE(test_se), 
        .CLK(n1659), .Q(\mem0[138][6] ), .QN(n24490) );
  SDFFX1 \mem0_reg[138][5]  ( .D(n17665), .SI(\mem0[138][4] ), .SE(test_se), 
        .CLK(n1659), .Q(\mem0[138][5] ), .QN(n24491) );
  SDFFX1 \mem0_reg[138][4]  ( .D(n17664), .SI(\mem0[138][3] ), .SE(test_se), 
        .CLK(n1659), .Q(\mem0[138][4] ), .QN(n24492) );
  SDFFX1 \mem0_reg[138][3]  ( .D(n17663), .SI(\mem0[138][2] ), .SE(test_se), 
        .CLK(n1659), .Q(\mem0[138][3] ), .QN(n24493) );
  SDFFX1 \mem0_reg[138][2]  ( .D(n17662), .SI(\mem0[138][1] ), .SE(test_se), 
        .CLK(n1659), .Q(\mem0[138][2] ), .QN(n24494) );
  SDFFX1 \mem0_reg[138][1]  ( .D(n17661), .SI(\mem0[138][0] ), .SE(test_se), 
        .CLK(n1659), .Q(\mem0[138][1] ), .QN(n24495) );
  SDFFX1 \mem0_reg[138][0]  ( .D(n17660), .SI(\mem0[137][7] ), .SE(test_se), 
        .CLK(n1659), .Q(\mem0[138][0] ), .QN(n24496) );
  SDFFX1 \mem0_reg[137][7]  ( .D(n17659), .SI(\mem0[137][6] ), .SE(test_se), 
        .CLK(n1659), .Q(\mem0[137][7] ), .QN(n24497) );
  SDFFX1 \mem0_reg[137][6]  ( .D(n17658), .SI(\mem0[137][5] ), .SE(test_se), 
        .CLK(n1659), .Q(\mem0[137][6] ), .QN(n24498) );
  SDFFX1 \mem0_reg[137][5]  ( .D(n17657), .SI(\mem0[137][4] ), .SE(test_se), 
        .CLK(n1660), .Q(\mem0[137][5] ), .QN(n24499) );
  SDFFX1 \mem0_reg[137][4]  ( .D(n17656), .SI(\mem0[137][3] ), .SE(test_se), 
        .CLK(n1660), .Q(\mem0[137][4] ), .QN(n24500) );
  SDFFX1 \mem0_reg[137][3]  ( .D(n17655), .SI(\mem0[137][2] ), .SE(test_se), 
        .CLK(n1660), .Q(\mem0[137][3] ), .QN(n24501) );
  SDFFX1 \mem0_reg[137][2]  ( .D(n17654), .SI(\mem0[137][1] ), .SE(test_se), 
        .CLK(n1660), .Q(\mem0[137][2] ), .QN(n24502) );
  SDFFX1 \mem0_reg[137][1]  ( .D(n17653), .SI(\mem0[137][0] ), .SE(test_se), 
        .CLK(n1660), .Q(\mem0[137][1] ), .QN(n24503) );
  SDFFX1 \mem0_reg[137][0]  ( .D(n17652), .SI(\mem0[136][7] ), .SE(test_se), 
        .CLK(n1660), .Q(\mem0[137][0] ), .QN(n24504) );
  SDFFX1 \mem0_reg[136][7]  ( .D(n17651), .SI(\mem0[136][6] ), .SE(test_se), 
        .CLK(n1660), .Q(\mem0[136][7] ), .QN(n24505) );
  SDFFX1 \mem0_reg[136][6]  ( .D(n17650), .SI(\mem0[136][5] ), .SE(test_se), 
        .CLK(n1660), .Q(\mem0[136][6] ), .QN(n24506) );
  SDFFX1 \mem0_reg[136][5]  ( .D(n17649), .SI(\mem0[136][4] ), .SE(test_se), 
        .CLK(n1660), .Q(\mem0[136][5] ), .QN(n24507) );
  SDFFX1 \mem0_reg[136][4]  ( .D(n17648), .SI(\mem0[136][3] ), .SE(test_se), 
        .CLK(n1660), .Q(\mem0[136][4] ), .QN(n24508) );
  SDFFX1 \mem0_reg[136][3]  ( .D(n17647), .SI(\mem0[136][2] ), .SE(test_se), 
        .CLK(n1660), .Q(\mem0[136][3] ), .QN(n24509) );
  SDFFX1 \mem0_reg[136][2]  ( .D(n17646), .SI(\mem0[136][1] ), .SE(test_se), 
        .CLK(n1660), .Q(\mem0[136][2] ), .QN(n24510) );
  SDFFX1 \mem0_reg[136][1]  ( .D(n17645), .SI(\mem0[136][0] ), .SE(test_se), 
        .CLK(n1661), .Q(\mem0[136][1] ), .QN(n24511) );
  SDFFX1 \mem0_reg[136][0]  ( .D(n17644), .SI(\mem0[135][7] ), .SE(test_se), 
        .CLK(n1661), .Q(\mem0[136][0] ), .QN(n24512) );
  SDFFX1 \mem0_reg[135][7]  ( .D(n17643), .SI(\mem0[135][6] ), .SE(test_se), 
        .CLK(n1661), .Q(\mem0[135][7] ), .QN(n24513) );
  SDFFX1 \mem0_reg[135][6]  ( .D(n17642), .SI(\mem0[135][5] ), .SE(test_se), 
        .CLK(n1661), .Q(\mem0[135][6] ), .QN(n24514) );
  SDFFX1 \mem0_reg[135][5]  ( .D(n17641), .SI(\mem0[135][4] ), .SE(test_se), 
        .CLK(n1661), .Q(\mem0[135][5] ), .QN(n24515) );
  SDFFX1 \mem0_reg[135][4]  ( .D(n17640), .SI(\mem0[135][3] ), .SE(test_se), 
        .CLK(n1661), .Q(\mem0[135][4] ), .QN(n24516) );
  SDFFX1 \mem0_reg[135][3]  ( .D(n17639), .SI(\mem0[135][2] ), .SE(test_se), 
        .CLK(n1661), .Q(\mem0[135][3] ), .QN(n24517) );
  SDFFX1 \mem0_reg[135][2]  ( .D(n17638), .SI(\mem0[135][1] ), .SE(test_se), 
        .CLK(n1661), .Q(\mem0[135][2] ), .QN(n24518) );
  SDFFX1 \mem0_reg[135][1]  ( .D(n17637), .SI(\mem0[135][0] ), .SE(test_se), 
        .CLK(n1661), .Q(\mem0[135][1] ), .QN(n24519) );
  SDFFX1 \mem0_reg[135][0]  ( .D(n17636), .SI(\mem0[134][7] ), .SE(test_se), 
        .CLK(n1661), .Q(\mem0[135][0] ), .QN(n24520) );
  SDFFX1 \mem0_reg[134][7]  ( .D(n17635), .SI(\mem0[134][6] ), .SE(test_se), 
        .CLK(n1661), .Q(\mem0[134][7] ), .QN(n24521) );
  SDFFX1 \mem0_reg[134][6]  ( .D(n17634), .SI(\mem0[134][5] ), .SE(test_se), 
        .CLK(n1661), .Q(\mem0[134][6] ), .QN(n24522) );
  SDFFX1 \mem0_reg[134][5]  ( .D(n17633), .SI(\mem0[134][4] ), .SE(test_se), 
        .CLK(n1662), .Q(\mem0[134][5] ), .QN(n24523) );
  SDFFX1 \mem0_reg[134][4]  ( .D(n17632), .SI(\mem0[134][3] ), .SE(test_se), 
        .CLK(n1662), .Q(\mem0[134][4] ), .QN(n24524) );
  SDFFX1 \mem0_reg[134][3]  ( .D(n17631), .SI(\mem0[134][2] ), .SE(test_se), 
        .CLK(n1662), .Q(\mem0[134][3] ), .QN(n24525) );
  SDFFX1 \mem0_reg[134][2]  ( .D(n17630), .SI(\mem0[134][1] ), .SE(test_se), 
        .CLK(n1662), .Q(\mem0[134][2] ), .QN(n24526) );
  SDFFX1 \mem0_reg[134][1]  ( .D(n17629), .SI(\mem0[134][0] ), .SE(test_se), 
        .CLK(n1662), .Q(\mem0[134][1] ), .QN(n24527) );
  SDFFX1 \mem0_reg[134][0]  ( .D(n17628), .SI(\mem0[133][7] ), .SE(test_se), 
        .CLK(n1662), .Q(\mem0[134][0] ), .QN(n24528) );
  SDFFX1 \mem0_reg[133][7]  ( .D(n17627), .SI(\mem0[133][6] ), .SE(test_se), 
        .CLK(n1662), .Q(\mem0[133][7] ), .QN(n24529) );
  SDFFX1 \mem0_reg[133][6]  ( .D(n17626), .SI(\mem0[133][5] ), .SE(test_se), 
        .CLK(n1662), .Q(\mem0[133][6] ), .QN(n24530) );
  SDFFX1 \mem0_reg[133][5]  ( .D(n17625), .SI(\mem0[133][4] ), .SE(test_se), 
        .CLK(n1662), .Q(\mem0[133][5] ), .QN(n24531) );
  SDFFX1 \mem0_reg[133][4]  ( .D(n17624), .SI(\mem0[133][3] ), .SE(test_se), 
        .CLK(n1662), .Q(\mem0[133][4] ), .QN(n24532) );
  SDFFX1 \mem0_reg[133][3]  ( .D(n17623), .SI(\mem0[133][2] ), .SE(test_se), 
        .CLK(n1662), .Q(\mem0[133][3] ), .QN(n24533) );
  SDFFX1 \mem0_reg[133][2]  ( .D(n17622), .SI(\mem0[133][1] ), .SE(test_se), 
        .CLK(n1662), .Q(\mem0[133][2] ), .QN(n24534) );
  SDFFX1 \mem0_reg[133][1]  ( .D(n17621), .SI(\mem0[133][0] ), .SE(test_se), 
        .CLK(n1663), .Q(\mem0[133][1] ), .QN(n24535) );
  SDFFX1 \mem0_reg[133][0]  ( .D(n17620), .SI(\mem0[132][7] ), .SE(test_se), 
        .CLK(n1663), .Q(\mem0[133][0] ), .QN(n24536) );
  SDFFX1 \mem0_reg[132][7]  ( .D(n17619), .SI(\mem0[132][6] ), .SE(test_se), 
        .CLK(n1663), .Q(\mem0[132][7] ), .QN(n24537) );
  SDFFX1 \mem0_reg[132][6]  ( .D(n17618), .SI(\mem0[132][5] ), .SE(test_se), 
        .CLK(n1663), .Q(\mem0[132][6] ), .QN(n24538) );
  SDFFX1 \mem0_reg[132][5]  ( .D(n17617), .SI(\mem0[132][4] ), .SE(test_se), 
        .CLK(n1663), .Q(\mem0[132][5] ), .QN(n24539) );
  SDFFX1 \mem0_reg[132][4]  ( .D(n17616), .SI(\mem0[132][3] ), .SE(test_se), 
        .CLK(n1663), .Q(\mem0[132][4] ), .QN(n24540) );
  SDFFX1 \mem0_reg[132][3]  ( .D(n17615), .SI(\mem0[132][2] ), .SE(test_se), 
        .CLK(n1663), .Q(\mem0[132][3] ), .QN(n24541) );
  SDFFX1 \mem0_reg[132][2]  ( .D(n17614), .SI(\mem0[132][1] ), .SE(test_se), 
        .CLK(n1663), .Q(\mem0[132][2] ), .QN(n24542) );
  SDFFX1 \mem0_reg[132][1]  ( .D(n17613), .SI(\mem0[132][0] ), .SE(test_se), 
        .CLK(n1663), .Q(\mem0[132][1] ), .QN(n24543) );
  SDFFX1 \mem0_reg[132][0]  ( .D(n17612), .SI(\mem0[131][7] ), .SE(test_se), 
        .CLK(n1663), .Q(\mem0[132][0] ), .QN(n24544) );
  SDFFX1 \mem0_reg[131][7]  ( .D(n17611), .SI(\mem0[131][6] ), .SE(test_se), 
        .CLK(n1663), .Q(\mem0[131][7] ), .QN(n24545) );
  SDFFX1 \mem0_reg[131][6]  ( .D(n17610), .SI(\mem0[131][5] ), .SE(test_se), 
        .CLK(n1663), .Q(\mem0[131][6] ), .QN(n24546) );
  SDFFX1 \mem0_reg[131][5]  ( .D(n17609), .SI(\mem0[131][4] ), .SE(test_se), 
        .CLK(n1664), .Q(\mem0[131][5] ), .QN(n24547) );
  SDFFX1 \mem0_reg[131][4]  ( .D(n17608), .SI(\mem0[131][3] ), .SE(test_se), 
        .CLK(n1664), .Q(\mem0[131][4] ), .QN(n24548) );
  SDFFX1 \mem0_reg[131][3]  ( .D(n17607), .SI(\mem0[131][2] ), .SE(test_se), 
        .CLK(n1664), .Q(\mem0[131][3] ), .QN(n24549) );
  SDFFX1 \mem0_reg[131][2]  ( .D(n17606), .SI(\mem0[131][1] ), .SE(test_se), 
        .CLK(n1664), .Q(\mem0[131][2] ), .QN(n24550) );
  SDFFX1 \mem0_reg[131][1]  ( .D(n17605), .SI(\mem0[131][0] ), .SE(test_se), 
        .CLK(n1664), .Q(\mem0[131][1] ), .QN(n24551) );
  SDFFX1 \mem0_reg[131][0]  ( .D(n17604), .SI(\mem0[130][7] ), .SE(test_se), 
        .CLK(n1664), .Q(\mem0[131][0] ), .QN(n24552) );
  SDFFX1 \mem0_reg[130][7]  ( .D(n17603), .SI(\mem0[130][6] ), .SE(test_se), 
        .CLK(n1664), .Q(\mem0[130][7] ), .QN(n24553) );
  SDFFX1 \mem0_reg[130][6]  ( .D(n17602), .SI(\mem0[130][5] ), .SE(test_se), 
        .CLK(n1664), .Q(\mem0[130][6] ), .QN(n24554) );
  SDFFX1 \mem0_reg[130][5]  ( .D(n17601), .SI(\mem0[130][4] ), .SE(test_se), 
        .CLK(n1664), .Q(\mem0[130][5] ), .QN(n24555) );
  SDFFX1 \mem0_reg[130][4]  ( .D(n17600), .SI(\mem0[130][3] ), .SE(test_se), 
        .CLK(n1664), .Q(\mem0[130][4] ), .QN(n24556) );
  SDFFX1 \mem0_reg[130][3]  ( .D(n17599), .SI(\mem0[130][2] ), .SE(test_se), 
        .CLK(n1664), .Q(\mem0[130][3] ), .QN(n24557) );
  SDFFX1 \mem0_reg[130][2]  ( .D(n17598), .SI(\mem0[130][1] ), .SE(test_se), 
        .CLK(n1664), .Q(\mem0[130][2] ), .QN(n24558) );
  SDFFX1 \mem0_reg[130][1]  ( .D(n17597), .SI(\mem0[130][0] ), .SE(test_se), 
        .CLK(n1665), .Q(\mem0[130][1] ), .QN(n24559) );
  SDFFX1 \mem0_reg[130][0]  ( .D(n17596), .SI(\mem0[129][7] ), .SE(test_se), 
        .CLK(n1665), .Q(\mem0[130][0] ), .QN(n24560) );
  SDFFX1 \mem0_reg[129][7]  ( .D(n17595), .SI(\mem0[129][6] ), .SE(test_se), 
        .CLK(n1665), .Q(\mem0[129][7] ), .QN(n24561) );
  SDFFX1 \mem0_reg[129][6]  ( .D(n17594), .SI(\mem0[129][5] ), .SE(test_se), 
        .CLK(n1665), .Q(\mem0[129][6] ), .QN(n24562) );
  SDFFX1 \mem0_reg[129][5]  ( .D(n17593), .SI(\mem0[129][4] ), .SE(test_se), 
        .CLK(n1665), .Q(\mem0[129][5] ), .QN(n24563) );
  SDFFX1 \mem0_reg[129][4]  ( .D(n17592), .SI(\mem0[129][3] ), .SE(test_se), 
        .CLK(n1665), .Q(\mem0[129][4] ), .QN(n24564) );
  SDFFX1 \mem0_reg[129][3]  ( .D(n17591), .SI(\mem0[129][2] ), .SE(test_se), 
        .CLK(n1665), .Q(\mem0[129][3] ), .QN(n24565) );
  SDFFX1 \mem0_reg[129][2]  ( .D(n17590), .SI(\mem0[129][1] ), .SE(test_se), 
        .CLK(n1665), .Q(\mem0[129][2] ), .QN(n24566) );
  SDFFX1 \mem0_reg[129][1]  ( .D(n17589), .SI(\mem0[129][0] ), .SE(test_se), 
        .CLK(n1665), .Q(\mem0[129][1] ), .QN(n24567) );
  SDFFX1 \mem0_reg[129][0]  ( .D(n17588), .SI(\mem0[128][7] ), .SE(test_se), 
        .CLK(n1665), .Q(\mem0[129][0] ), .QN(n24568) );
  SDFFX1 \mem0_reg[128][7]  ( .D(n17587), .SI(\mem0[128][6] ), .SE(test_se), 
        .CLK(n1665), .Q(\mem0[128][7] ), .QN(n24569) );
  SDFFX1 \mem0_reg[128][6]  ( .D(n17586), .SI(\mem0[128][5] ), .SE(test_se), 
        .CLK(n1665), .Q(\mem0[128][6] ), .QN(n24570) );
  SDFFX1 \mem0_reg[128][5]  ( .D(n17585), .SI(\mem0[128][4] ), .SE(test_se), 
        .CLK(n1666), .Q(\mem0[128][5] ), .QN(n24571) );
  SDFFX1 \mem0_reg[128][4]  ( .D(n17584), .SI(\mem0[128][3] ), .SE(test_se), 
        .CLK(n1666), .Q(\mem0[128][4] ), .QN(n24572) );
  SDFFX1 \mem0_reg[128][3]  ( .D(n17583), .SI(\mem0[128][2] ), .SE(test_se), 
        .CLK(n1666), .Q(\mem0[128][3] ), .QN(n24573) );
  SDFFX1 \mem0_reg[128][2]  ( .D(n17582), .SI(\mem0[128][1] ), .SE(test_se), 
        .CLK(n1666), .Q(\mem0[128][2] ), .QN(n24574) );
  SDFFX1 \mem0_reg[128][1]  ( .D(n17581), .SI(\mem0[128][0] ), .SE(test_se), 
        .CLK(n1666), .Q(\mem0[128][1] ), .QN(n24575) );
  SDFFX1 \mem0_reg[128][0]  ( .D(n17580), .SI(\mem0[127][7] ), .SE(test_se), 
        .CLK(n1666), .Q(\mem0[128][0] ), .QN(n24576) );
  SDFFX1 \mem0_reg[127][7]  ( .D(n17579), .SI(\mem0[127][6] ), .SE(test_se), 
        .CLK(n1666), .Q(\mem0[127][7] ), .QN(n24577) );
  SDFFX1 \mem0_reg[127][6]  ( .D(n17578), .SI(\mem0[127][5] ), .SE(test_se), 
        .CLK(n1666), .Q(\mem0[127][6] ), .QN(n24578) );
  SDFFX1 \mem0_reg[127][5]  ( .D(n17577), .SI(\mem0[127][4] ), .SE(test_se), 
        .CLK(n1666), .Q(\mem0[127][5] ), .QN(n24579) );
  SDFFX1 \mem0_reg[127][4]  ( .D(n17576), .SI(\mem0[127][3] ), .SE(test_se), 
        .CLK(n1666), .Q(\mem0[127][4] ), .QN(n24580) );
  SDFFX1 \mem0_reg[127][3]  ( .D(n17575), .SI(\mem0[127][2] ), .SE(test_se), 
        .CLK(n1666), .Q(\mem0[127][3] ), .QN(n24581) );
  SDFFX1 \mem0_reg[127][2]  ( .D(n17574), .SI(\mem0[127][1] ), .SE(test_se), 
        .CLK(n1666), .Q(\mem0[127][2] ), .QN(n24582) );
  SDFFX1 \mem0_reg[127][1]  ( .D(n17573), .SI(\mem0[127][0] ), .SE(test_se), 
        .CLK(n1667), .Q(\mem0[127][1] ), .QN(n24583) );
  SDFFX1 \mem0_reg[127][0]  ( .D(n17572), .SI(\mem0[126][7] ), .SE(test_se), 
        .CLK(n1667), .Q(\mem0[127][0] ), .QN(n24584) );
  SDFFX1 \mem0_reg[126][7]  ( .D(n17571), .SI(\mem0[126][6] ), .SE(test_se), 
        .CLK(n1667), .Q(\mem0[126][7] ), .QN(n24585) );
  SDFFX1 \mem0_reg[126][6]  ( .D(n17570), .SI(\mem0[126][5] ), .SE(test_se), 
        .CLK(n1667), .Q(\mem0[126][6] ), .QN(n24586) );
  SDFFX1 \mem0_reg[126][5]  ( .D(n17569), .SI(\mem0[126][4] ), .SE(test_se), 
        .CLK(n1667), .Q(\mem0[126][5] ), .QN(n24587) );
  SDFFX1 \mem0_reg[126][4]  ( .D(n17568), .SI(\mem0[126][3] ), .SE(test_se), 
        .CLK(n1667), .Q(\mem0[126][4] ), .QN(n24588) );
  SDFFX1 \mem0_reg[126][3]  ( .D(n17567), .SI(\mem0[126][2] ), .SE(test_se), 
        .CLK(n1667), .Q(\mem0[126][3] ), .QN(n24589) );
  SDFFX1 \mem0_reg[126][2]  ( .D(n17566), .SI(\mem0[126][1] ), .SE(test_se), 
        .CLK(n1667), .Q(\mem0[126][2] ), .QN(n24590) );
  SDFFX1 \mem0_reg[126][1]  ( .D(n17565), .SI(\mem0[126][0] ), .SE(test_se), 
        .CLK(n1667), .Q(\mem0[126][1] ), .QN(n24591) );
  SDFFX1 \mem0_reg[126][0]  ( .D(n17564), .SI(\mem0[125][7] ), .SE(test_se), 
        .CLK(n1667), .Q(\mem0[126][0] ), .QN(n24592) );
  SDFFX1 \mem0_reg[125][7]  ( .D(n17563), .SI(\mem0[125][6] ), .SE(test_se), 
        .CLK(n1667), .Q(\mem0[125][7] ), .QN(n24593) );
  SDFFX1 \mem0_reg[125][6]  ( .D(n17562), .SI(\mem0[125][5] ), .SE(test_se), 
        .CLK(n1667), .Q(\mem0[125][6] ), .QN(n24594) );
  SDFFX1 \mem0_reg[125][5]  ( .D(n17561), .SI(\mem0[125][4] ), .SE(test_se), 
        .CLK(n1668), .Q(\mem0[125][5] ), .QN(n24595) );
  SDFFX1 \mem0_reg[125][4]  ( .D(n17560), .SI(\mem0[125][3] ), .SE(test_se), 
        .CLK(n1668), .Q(\mem0[125][4] ), .QN(n24596) );
  SDFFX1 \mem0_reg[125][3]  ( .D(n17559), .SI(\mem0[125][2] ), .SE(test_se), 
        .CLK(n1668), .Q(\mem0[125][3] ), .QN(n24597) );
  SDFFX1 \mem0_reg[125][2]  ( .D(n17558), .SI(\mem0[125][1] ), .SE(test_se), 
        .CLK(n1668), .Q(\mem0[125][2] ), .QN(n24598) );
  SDFFX1 \mem0_reg[125][1]  ( .D(n17557), .SI(\mem0[125][0] ), .SE(test_se), 
        .CLK(n1668), .Q(\mem0[125][1] ), .QN(n24599) );
  SDFFX1 \mem0_reg[125][0]  ( .D(n17556), .SI(\mem0[124][7] ), .SE(test_se), 
        .CLK(n1668), .Q(\mem0[125][0] ), .QN(n24600) );
  SDFFX1 \mem0_reg[124][7]  ( .D(n17555), .SI(\mem0[124][6] ), .SE(test_se), 
        .CLK(n1668), .Q(\mem0[124][7] ), .QN(n24601) );
  SDFFX1 \mem0_reg[124][6]  ( .D(n17554), .SI(\mem0[124][5] ), .SE(test_se), 
        .CLK(n1668), .Q(\mem0[124][6] ), .QN(n24602) );
  SDFFX1 \mem0_reg[124][5]  ( .D(n17553), .SI(\mem0[124][4] ), .SE(test_se), 
        .CLK(n1668), .Q(\mem0[124][5] ), .QN(n24603) );
  SDFFX1 \mem0_reg[124][4]  ( .D(n17552), .SI(\mem0[124][3] ), .SE(test_se), 
        .CLK(n1668), .Q(\mem0[124][4] ), .QN(n24604) );
  SDFFX1 \mem0_reg[124][3]  ( .D(n17551), .SI(\mem0[124][2] ), .SE(test_se), 
        .CLK(n1668), .Q(\mem0[124][3] ), .QN(n24605) );
  SDFFX1 \mem0_reg[124][2]  ( .D(n17550), .SI(\mem0[124][1] ), .SE(test_se), 
        .CLK(n1668), .Q(\mem0[124][2] ), .QN(n24606) );
  SDFFX1 \mem0_reg[124][1]  ( .D(n17549), .SI(\mem0[124][0] ), .SE(test_se), 
        .CLK(n1669), .Q(\mem0[124][1] ), .QN(n24607) );
  SDFFX1 \mem0_reg[124][0]  ( .D(n17548), .SI(\mem0[123][7] ), .SE(test_se), 
        .CLK(n1669), .Q(\mem0[124][0] ), .QN(n24608) );
  SDFFX1 \mem0_reg[123][7]  ( .D(n17547), .SI(\mem0[123][6] ), .SE(test_se), 
        .CLK(n1669), .Q(\mem0[123][7] ), .QN(n24609) );
  SDFFX1 \mem0_reg[123][6]  ( .D(n17546), .SI(\mem0[123][5] ), .SE(test_se), 
        .CLK(n1669), .Q(\mem0[123][6] ), .QN(n24610) );
  SDFFX1 \mem0_reg[123][5]  ( .D(n17545), .SI(\mem0[123][4] ), .SE(test_se), 
        .CLK(n1669), .Q(\mem0[123][5] ), .QN(n24611) );
  SDFFX1 \mem0_reg[123][4]  ( .D(n17544), .SI(\mem0[123][3] ), .SE(test_se), 
        .CLK(n1669), .Q(\mem0[123][4] ), .QN(n24612) );
  SDFFX1 \mem0_reg[123][3]  ( .D(n17543), .SI(\mem0[123][2] ), .SE(test_se), 
        .CLK(n1669), .Q(\mem0[123][3] ), .QN(n24613) );
  SDFFX1 \mem0_reg[123][2]  ( .D(n17542), .SI(\mem0[123][1] ), .SE(test_se), 
        .CLK(n1669), .Q(\mem0[123][2] ), .QN(n24614) );
  SDFFX1 \mem0_reg[123][1]  ( .D(n17541), .SI(\mem0[123][0] ), .SE(test_se), 
        .CLK(n1669), .Q(\mem0[123][1] ), .QN(n24615) );
  SDFFX1 \mem0_reg[123][0]  ( .D(n17540), .SI(\mem0[122][7] ), .SE(test_se), 
        .CLK(n1669), .Q(\mem0[123][0] ), .QN(n24616) );
  SDFFX1 \mem0_reg[122][7]  ( .D(n17539), .SI(\mem0[122][6] ), .SE(test_se), 
        .CLK(n1669), .Q(\mem0[122][7] ), .QN(n24617) );
  SDFFX1 \mem0_reg[122][6]  ( .D(n17538), .SI(\mem0[122][5] ), .SE(test_se), 
        .CLK(n1669), .Q(\mem0[122][6] ), .QN(n24618) );
  SDFFX1 \mem0_reg[122][5]  ( .D(n17537), .SI(\mem0[122][4] ), .SE(test_se), 
        .CLK(n1670), .Q(\mem0[122][5] ), .QN(n24619) );
  SDFFX1 \mem0_reg[122][4]  ( .D(n17536), .SI(\mem0[122][3] ), .SE(test_se), 
        .CLK(n1670), .Q(\mem0[122][4] ), .QN(n24620) );
  SDFFX1 \mem0_reg[122][3]  ( .D(n17535), .SI(\mem0[122][2] ), .SE(test_se), 
        .CLK(n1670), .Q(\mem0[122][3] ), .QN(n24621) );
  SDFFX1 \mem0_reg[122][2]  ( .D(n17534), .SI(\mem0[122][1] ), .SE(test_se), 
        .CLK(n1670), .Q(\mem0[122][2] ), .QN(n24622) );
  SDFFX1 \mem0_reg[122][1]  ( .D(n17533), .SI(\mem0[122][0] ), .SE(test_se), 
        .CLK(n1670), .Q(\mem0[122][1] ), .QN(n24623) );
  SDFFX1 \mem0_reg[122][0]  ( .D(n17532), .SI(\mem0[121][7] ), .SE(test_se), 
        .CLK(n1670), .Q(\mem0[122][0] ), .QN(n24624) );
  SDFFX1 \mem0_reg[121][7]  ( .D(n17531), .SI(\mem0[121][6] ), .SE(test_se), 
        .CLK(n1670), .Q(\mem0[121][7] ), .QN(n24625) );
  SDFFX1 \mem0_reg[121][6]  ( .D(n17530), .SI(\mem0[121][5] ), .SE(test_se), 
        .CLK(n1670), .Q(\mem0[121][6] ), .QN(n24626) );
  SDFFX1 \mem0_reg[121][5]  ( .D(n17529), .SI(\mem0[121][4] ), .SE(test_se), 
        .CLK(n1670), .Q(\mem0[121][5] ), .QN(n24627) );
  SDFFX1 \mem0_reg[121][4]  ( .D(n17528), .SI(\mem0[121][3] ), .SE(test_se), 
        .CLK(n1670), .Q(\mem0[121][4] ), .QN(n24628) );
  SDFFX1 \mem0_reg[121][3]  ( .D(n17527), .SI(\mem0[121][2] ), .SE(test_se), 
        .CLK(n1670), .Q(\mem0[121][3] ), .QN(n24629) );
  SDFFX1 \mem0_reg[121][2]  ( .D(n17526), .SI(\mem0[121][1] ), .SE(test_se), 
        .CLK(n1670), .Q(\mem0[121][2] ), .QN(n24630) );
  SDFFX1 \mem0_reg[121][1]  ( .D(n17525), .SI(\mem0[121][0] ), .SE(test_se), 
        .CLK(n1671), .Q(\mem0[121][1] ), .QN(n24631) );
  SDFFX1 \mem0_reg[121][0]  ( .D(n17524), .SI(\mem0[120][7] ), .SE(test_se), 
        .CLK(n1671), .Q(\mem0[121][0] ), .QN(n24632) );
  SDFFX1 \mem0_reg[120][7]  ( .D(n17523), .SI(\mem0[120][6] ), .SE(test_se), 
        .CLK(n1671), .Q(\mem0[120][7] ), .QN(n24633) );
  SDFFX1 \mem0_reg[120][6]  ( .D(n17522), .SI(\mem0[120][5] ), .SE(test_se), 
        .CLK(n1671), .Q(\mem0[120][6] ), .QN(n24634) );
  SDFFX1 \mem0_reg[120][5]  ( .D(n17521), .SI(\mem0[120][4] ), .SE(test_se), 
        .CLK(n1671), .Q(\mem0[120][5] ), .QN(n24635) );
  SDFFX1 \mem0_reg[120][4]  ( .D(n17520), .SI(\mem0[120][3] ), .SE(test_se), 
        .CLK(n1671), .Q(\mem0[120][4] ), .QN(n24636) );
  SDFFX1 \mem0_reg[120][3]  ( .D(n17519), .SI(\mem0[120][2] ), .SE(test_se), 
        .CLK(n1671), .Q(\mem0[120][3] ), .QN(n24637) );
  SDFFX1 \mem0_reg[120][2]  ( .D(n17518), .SI(\mem0[120][1] ), .SE(test_se), 
        .CLK(n1671), .Q(\mem0[120][2] ), .QN(n24638) );
  SDFFX1 \mem0_reg[120][1]  ( .D(n17517), .SI(\mem0[120][0] ), .SE(test_se), 
        .CLK(n1671), .Q(\mem0[120][1] ), .QN(n24639) );
  SDFFX1 \mem0_reg[120][0]  ( .D(n17516), .SI(\mem0[119][7] ), .SE(test_se), 
        .CLK(n1671), .Q(\mem0[120][0] ), .QN(n24640) );
  SDFFX1 \mem0_reg[119][7]  ( .D(n17515), .SI(\mem0[119][6] ), .SE(test_se), 
        .CLK(n1671), .Q(\mem0[119][7] ), .QN(n24641) );
  SDFFX1 \mem0_reg[119][6]  ( .D(n17514), .SI(\mem0[119][5] ), .SE(test_se), 
        .CLK(n1671), .Q(\mem0[119][6] ), .QN(n24642) );
  SDFFX1 \mem0_reg[119][5]  ( .D(n17513), .SI(\mem0[119][4] ), .SE(test_se), 
        .CLK(n1672), .Q(\mem0[119][5] ), .QN(n24643) );
  SDFFX1 \mem0_reg[119][4]  ( .D(n17512), .SI(\mem0[119][3] ), .SE(test_se), 
        .CLK(n1672), .Q(\mem0[119][4] ), .QN(n24644) );
  SDFFX1 \mem0_reg[119][3]  ( .D(n17511), .SI(\mem0[119][2] ), .SE(test_se), 
        .CLK(n1672), .Q(\mem0[119][3] ), .QN(n24645) );
  SDFFX1 \mem0_reg[119][2]  ( .D(n17510), .SI(\mem0[119][1] ), .SE(test_se), 
        .CLK(n1672), .Q(\mem0[119][2] ), .QN(n24646) );
  SDFFX1 \mem0_reg[119][1]  ( .D(n17509), .SI(\mem0[119][0] ), .SE(test_se), 
        .CLK(n1672), .Q(\mem0[119][1] ), .QN(n24647) );
  SDFFX1 \mem0_reg[119][0]  ( .D(n17508), .SI(\mem0[118][7] ), .SE(test_se), 
        .CLK(n1672), .Q(\mem0[119][0] ), .QN(n24648) );
  SDFFX1 \mem0_reg[118][7]  ( .D(n17507), .SI(\mem0[118][6] ), .SE(test_se), 
        .CLK(n1672), .Q(\mem0[118][7] ), .QN(n24649) );
  SDFFX1 \mem0_reg[118][6]  ( .D(n17506), .SI(\mem0[118][5] ), .SE(test_se), 
        .CLK(n1672), .Q(\mem0[118][6] ), .QN(n24650) );
  SDFFX1 \mem0_reg[118][5]  ( .D(n17505), .SI(\mem0[118][4] ), .SE(test_se), 
        .CLK(n1672), .Q(\mem0[118][5] ), .QN(n24651) );
  SDFFX1 \mem0_reg[118][4]  ( .D(n17504), .SI(\mem0[118][3] ), .SE(test_se), 
        .CLK(n1672), .Q(\mem0[118][4] ), .QN(n24652) );
  SDFFX1 \mem0_reg[118][3]  ( .D(n17503), .SI(\mem0[118][2] ), .SE(test_se), 
        .CLK(n1672), .Q(\mem0[118][3] ), .QN(n24653) );
  SDFFX1 \mem0_reg[118][2]  ( .D(n17502), .SI(\mem0[118][1] ), .SE(test_se), 
        .CLK(n1672), .Q(\mem0[118][2] ), .QN(n24654) );
  SDFFX1 \mem0_reg[118][1]  ( .D(n17501), .SI(\mem0[118][0] ), .SE(test_se), 
        .CLK(n1673), .Q(\mem0[118][1] ), .QN(n24655) );
  SDFFX1 \mem0_reg[118][0]  ( .D(n17500), .SI(\mem0[117][7] ), .SE(test_se), 
        .CLK(n1673), .Q(\mem0[118][0] ), .QN(n24656) );
  SDFFX1 \mem0_reg[117][7]  ( .D(n17499), .SI(\mem0[117][6] ), .SE(test_se), 
        .CLK(n1673), .Q(\mem0[117][7] ), .QN(n24657) );
  SDFFX1 \mem0_reg[117][6]  ( .D(n17498), .SI(\mem0[117][5] ), .SE(test_se), 
        .CLK(n1673), .Q(\mem0[117][6] ), .QN(n24658) );
  SDFFX1 \mem0_reg[117][5]  ( .D(n17497), .SI(\mem0[117][4] ), .SE(test_se), 
        .CLK(n1673), .Q(\mem0[117][5] ), .QN(n24659) );
  SDFFX1 \mem0_reg[117][4]  ( .D(n17496), .SI(\mem0[117][3] ), .SE(test_se), 
        .CLK(n1673), .Q(\mem0[117][4] ), .QN(n24660) );
  SDFFX1 \mem0_reg[117][3]  ( .D(n17495), .SI(\mem0[117][2] ), .SE(test_se), 
        .CLK(n1673), .Q(\mem0[117][3] ), .QN(n24661) );
  SDFFX1 \mem0_reg[117][2]  ( .D(n17494), .SI(\mem0[117][1] ), .SE(test_se), 
        .CLK(n1673), .Q(\mem0[117][2] ), .QN(n24662) );
  SDFFX1 \mem0_reg[117][1]  ( .D(n17493), .SI(\mem0[117][0] ), .SE(test_se), 
        .CLK(n1673), .Q(\mem0[117][1] ), .QN(n24663) );
  SDFFX1 \mem0_reg[117][0]  ( .D(n17492), .SI(\mem0[116][7] ), .SE(test_se), 
        .CLK(n1673), .Q(\mem0[117][0] ), .QN(n24664) );
  SDFFX1 \mem0_reg[116][7]  ( .D(n17491), .SI(\mem0[116][6] ), .SE(test_se), 
        .CLK(n1673), .Q(\mem0[116][7] ), .QN(n24665) );
  SDFFX1 \mem0_reg[116][6]  ( .D(n17490), .SI(\mem0[116][5] ), .SE(test_se), 
        .CLK(n1673), .Q(\mem0[116][6] ), .QN(n24666) );
  SDFFX1 \mem0_reg[116][5]  ( .D(n17489), .SI(\mem0[116][4] ), .SE(test_se), 
        .CLK(n1674), .Q(\mem0[116][5] ), .QN(n24667) );
  SDFFX1 \mem0_reg[116][4]  ( .D(n17488), .SI(\mem0[116][3] ), .SE(test_se), 
        .CLK(n1674), .Q(\mem0[116][4] ), .QN(n24668) );
  SDFFX1 \mem0_reg[116][3]  ( .D(n17487), .SI(\mem0[116][2] ), .SE(test_se), 
        .CLK(n1674), .Q(\mem0[116][3] ), .QN(n24669) );
  SDFFX1 \mem0_reg[116][2]  ( .D(n17486), .SI(\mem0[116][1] ), .SE(test_se), 
        .CLK(n1674), .Q(\mem0[116][2] ), .QN(n24670) );
  SDFFX1 \mem0_reg[116][1]  ( .D(n17485), .SI(\mem0[116][0] ), .SE(test_se), 
        .CLK(n1674), .Q(\mem0[116][1] ), .QN(n24671) );
  SDFFX1 \mem0_reg[116][0]  ( .D(n17484), .SI(\mem0[115][7] ), .SE(test_se), 
        .CLK(n1674), .Q(\mem0[116][0] ), .QN(n24672) );
  SDFFX1 \mem0_reg[115][7]  ( .D(n17483), .SI(\mem0[115][6] ), .SE(test_se), 
        .CLK(n1674), .Q(\mem0[115][7] ), .QN(n24673) );
  SDFFX1 \mem0_reg[115][6]  ( .D(n17482), .SI(\mem0[115][5] ), .SE(test_se), 
        .CLK(n1674), .Q(\mem0[115][6] ), .QN(n24674) );
  SDFFX1 \mem0_reg[115][5]  ( .D(n17481), .SI(\mem0[115][4] ), .SE(test_se), 
        .CLK(n1674), .Q(\mem0[115][5] ), .QN(n24675) );
  SDFFX1 \mem0_reg[115][4]  ( .D(n17480), .SI(\mem0[115][3] ), .SE(test_se), 
        .CLK(n1674), .Q(\mem0[115][4] ), .QN(n24676) );
  SDFFX1 \mem0_reg[115][3]  ( .D(n17479), .SI(\mem0[115][2] ), .SE(test_se), 
        .CLK(n1674), .Q(\mem0[115][3] ), .QN(n24677) );
  SDFFX1 \mem0_reg[115][2]  ( .D(n17478), .SI(\mem0[115][1] ), .SE(test_se), 
        .CLK(n1674), .Q(\mem0[115][2] ), .QN(n24678) );
  SDFFX1 \mem0_reg[115][1]  ( .D(n17477), .SI(\mem0[115][0] ), .SE(test_se), 
        .CLK(n1675), .Q(\mem0[115][1] ), .QN(n24679) );
  SDFFX1 \mem0_reg[115][0]  ( .D(n17476), .SI(\mem0[114][7] ), .SE(test_se), 
        .CLK(n1675), .Q(\mem0[115][0] ), .QN(n24680) );
  SDFFX1 \mem0_reg[114][7]  ( .D(n17475), .SI(\mem0[114][6] ), .SE(test_se), 
        .CLK(n1675), .Q(\mem0[114][7] ), .QN(n24681) );
  SDFFX1 \mem0_reg[114][6]  ( .D(n17474), .SI(\mem0[114][5] ), .SE(test_se), 
        .CLK(n1675), .Q(\mem0[114][6] ), .QN(n24682) );
  SDFFX1 \mem0_reg[114][5]  ( .D(n17473), .SI(\mem0[114][4] ), .SE(test_se), 
        .CLK(n1675), .Q(\mem0[114][5] ), .QN(n24683) );
  SDFFX1 \mem0_reg[114][4]  ( .D(n17472), .SI(\mem0[114][3] ), .SE(test_se), 
        .CLK(n1675), .Q(\mem0[114][4] ), .QN(n24684) );
  SDFFX1 \mem0_reg[114][3]  ( .D(n17471), .SI(\mem0[114][2] ), .SE(test_se), 
        .CLK(n1675), .Q(\mem0[114][3] ), .QN(n24685) );
  SDFFX1 \mem0_reg[114][2]  ( .D(n17470), .SI(\mem0[114][1] ), .SE(test_se), 
        .CLK(n1675), .Q(\mem0[114][2] ), .QN(n24686) );
  SDFFX1 \mem0_reg[114][1]  ( .D(n17469), .SI(\mem0[114][0] ), .SE(test_se), 
        .CLK(n1675), .Q(\mem0[114][1] ), .QN(n24687) );
  SDFFX1 \mem0_reg[114][0]  ( .D(n17468), .SI(\mem0[113][7] ), .SE(test_se), 
        .CLK(n1675), .Q(\mem0[114][0] ), .QN(n24688) );
  SDFFX1 \mem0_reg[113][7]  ( .D(n17467), .SI(\mem0[113][6] ), .SE(test_se), 
        .CLK(n1675), .Q(\mem0[113][7] ), .QN(n24689) );
  SDFFX1 \mem0_reg[113][6]  ( .D(n17466), .SI(\mem0[113][5] ), .SE(test_se), 
        .CLK(n1675), .Q(\mem0[113][6] ), .QN(n24690) );
  SDFFX1 \mem0_reg[113][5]  ( .D(n17465), .SI(\mem0[113][4] ), .SE(test_se), 
        .CLK(n1676), .Q(\mem0[113][5] ), .QN(n24691) );
  SDFFX1 \mem0_reg[113][4]  ( .D(n17464), .SI(\mem0[113][3] ), .SE(test_se), 
        .CLK(n1676), .Q(\mem0[113][4] ), .QN(n24692) );
  SDFFX1 \mem0_reg[113][3]  ( .D(n17463), .SI(\mem0[113][2] ), .SE(test_se), 
        .CLK(n1676), .Q(\mem0[113][3] ), .QN(n24693) );
  SDFFX1 \mem0_reg[113][2]  ( .D(n17462), .SI(\mem0[113][1] ), .SE(test_se), 
        .CLK(n1676), .Q(\mem0[113][2] ), .QN(n24694) );
  SDFFX1 \mem0_reg[113][1]  ( .D(n17461), .SI(\mem0[113][0] ), .SE(test_se), 
        .CLK(n1676), .Q(\mem0[113][1] ), .QN(n24695) );
  SDFFX1 \mem0_reg[113][0]  ( .D(n17460), .SI(\mem0[112][7] ), .SE(test_se), 
        .CLK(n1676), .Q(\mem0[113][0] ), .QN(n24696) );
  SDFFX1 \mem0_reg[112][7]  ( .D(n17459), .SI(\mem0[112][6] ), .SE(test_se), 
        .CLK(n1676), .Q(\mem0[112][7] ), .QN(n24697) );
  SDFFX1 \mem0_reg[112][6]  ( .D(n17458), .SI(\mem0[112][5] ), .SE(test_se), 
        .CLK(n1676), .Q(\mem0[112][6] ), .QN(n24698) );
  SDFFX1 \mem0_reg[112][5]  ( .D(n17457), .SI(\mem0[112][4] ), .SE(test_se), 
        .CLK(n1676), .Q(\mem0[112][5] ), .QN(n24699) );
  SDFFX1 \mem0_reg[112][4]  ( .D(n17456), .SI(\mem0[112][3] ), .SE(test_se), 
        .CLK(n1676), .Q(\mem0[112][4] ), .QN(n24700) );
  SDFFX1 \mem0_reg[112][3]  ( .D(n17455), .SI(\mem0[112][2] ), .SE(test_se), 
        .CLK(n1676), .Q(\mem0[112][3] ), .QN(n24701) );
  SDFFX1 \mem0_reg[112][2]  ( .D(n17454), .SI(\mem0[112][1] ), .SE(test_se), 
        .CLK(n1676), .Q(\mem0[112][2] ), .QN(n24702) );
  SDFFX1 \mem0_reg[112][1]  ( .D(n17453), .SI(\mem0[112][0] ), .SE(test_se), 
        .CLK(n1677), .Q(\mem0[112][1] ), .QN(n24703) );
  SDFFX1 \mem0_reg[112][0]  ( .D(n17452), .SI(\mem0[111][7] ), .SE(test_se), 
        .CLK(n1677), .Q(\mem0[112][0] ), .QN(n24704) );
  SDFFX1 \mem0_reg[111][7]  ( .D(n17451), .SI(\mem0[111][6] ), .SE(test_se), 
        .CLK(n1677), .Q(\mem0[111][7] ), .QN(n24705) );
  SDFFX1 \mem0_reg[111][6]  ( .D(n17450), .SI(\mem0[111][5] ), .SE(test_se), 
        .CLK(n1677), .Q(\mem0[111][6] ), .QN(n24706) );
  SDFFX1 \mem0_reg[111][5]  ( .D(n17449), .SI(\mem0[111][4] ), .SE(test_se), 
        .CLK(n1677), .Q(\mem0[111][5] ), .QN(n24707) );
  SDFFX1 \mem0_reg[111][4]  ( .D(n17448), .SI(\mem0[111][3] ), .SE(test_se), 
        .CLK(n1677), .Q(\mem0[111][4] ), .QN(n24708) );
  SDFFX1 \mem0_reg[111][3]  ( .D(n17447), .SI(\mem0[111][2] ), .SE(test_se), 
        .CLK(n1677), .Q(\mem0[111][3] ), .QN(n24709) );
  SDFFX1 \mem0_reg[111][2]  ( .D(n17446), .SI(\mem0[111][1] ), .SE(test_se), 
        .CLK(n1677), .Q(\mem0[111][2] ), .QN(n24710) );
  SDFFX1 \mem0_reg[111][1]  ( .D(n17445), .SI(\mem0[111][0] ), .SE(test_se), 
        .CLK(n1677), .Q(\mem0[111][1] ), .QN(n24711) );
  SDFFX1 \mem0_reg[111][0]  ( .D(n17444), .SI(\mem0[110][7] ), .SE(test_se), 
        .CLK(n1677), .Q(\mem0[111][0] ), .QN(n24712) );
  SDFFX1 \mem0_reg[110][7]  ( .D(n17443), .SI(\mem0[110][6] ), .SE(test_se), 
        .CLK(n1677), .Q(\mem0[110][7] ), .QN(n24713) );
  SDFFX1 \mem0_reg[110][6]  ( .D(n17442), .SI(\mem0[110][5] ), .SE(test_se), 
        .CLK(n1677), .Q(\mem0[110][6] ), .QN(n24714) );
  SDFFX1 \mem0_reg[110][5]  ( .D(n17441), .SI(\mem0[110][4] ), .SE(test_se), 
        .CLK(n1678), .Q(\mem0[110][5] ), .QN(n24715) );
  SDFFX1 \mem0_reg[110][4]  ( .D(n17440), .SI(\mem0[110][3] ), .SE(test_se), 
        .CLK(n1678), .Q(\mem0[110][4] ), .QN(n24716) );
  SDFFX1 \mem0_reg[110][3]  ( .D(n17439), .SI(\mem0[110][2] ), .SE(test_se), 
        .CLK(n1678), .Q(\mem0[110][3] ), .QN(n24717) );
  SDFFX1 \mem0_reg[110][2]  ( .D(n17438), .SI(\mem0[110][1] ), .SE(test_se), 
        .CLK(n1678), .Q(\mem0[110][2] ), .QN(n24718) );
  SDFFX1 \mem0_reg[110][1]  ( .D(n17437), .SI(\mem0[110][0] ), .SE(test_se), 
        .CLK(n1678), .Q(\mem0[110][1] ), .QN(n24719) );
  SDFFX1 \mem0_reg[110][0]  ( .D(n17436), .SI(\mem0[109][7] ), .SE(test_se), 
        .CLK(n1678), .Q(\mem0[110][0] ), .QN(n24720) );
  SDFFX1 \mem0_reg[109][7]  ( .D(n17435), .SI(\mem0[109][6] ), .SE(test_se), 
        .CLK(n1678), .Q(\mem0[109][7] ), .QN(n24721) );
  SDFFX1 \mem0_reg[109][6]  ( .D(n17434), .SI(\mem0[109][5] ), .SE(test_se), 
        .CLK(n1678), .Q(\mem0[109][6] ), .QN(n24722) );
  SDFFX1 \mem0_reg[109][5]  ( .D(n17433), .SI(\mem0[109][4] ), .SE(test_se), 
        .CLK(n1678), .Q(\mem0[109][5] ), .QN(n24723) );
  SDFFX1 \mem0_reg[109][4]  ( .D(n17432), .SI(\mem0[109][3] ), .SE(test_se), 
        .CLK(n1678), .Q(\mem0[109][4] ), .QN(n24724) );
  SDFFX1 \mem0_reg[109][3]  ( .D(n17431), .SI(\mem0[109][2] ), .SE(test_se), 
        .CLK(n1678), .Q(\mem0[109][3] ), .QN(n24725) );
  SDFFX1 \mem0_reg[109][2]  ( .D(n17430), .SI(\mem0[109][1] ), .SE(test_se), 
        .CLK(n1678), .Q(\mem0[109][2] ), .QN(n24726) );
  SDFFX1 \mem0_reg[109][1]  ( .D(n17429), .SI(\mem0[109][0] ), .SE(test_se), 
        .CLK(n1679), .Q(\mem0[109][1] ), .QN(n24727) );
  SDFFX1 \mem0_reg[109][0]  ( .D(n17428), .SI(\mem0[108][7] ), .SE(test_se), 
        .CLK(n1679), .Q(\mem0[109][0] ), .QN(n24728) );
  SDFFX1 \mem0_reg[108][7]  ( .D(n17427), .SI(\mem0[108][6] ), .SE(test_se), 
        .CLK(n1679), .Q(\mem0[108][7] ), .QN(n24729) );
  SDFFX1 \mem0_reg[108][6]  ( .D(n17426), .SI(\mem0[108][5] ), .SE(test_se), 
        .CLK(n1679), .Q(\mem0[108][6] ), .QN(n24730) );
  SDFFX1 \mem0_reg[108][5]  ( .D(n17425), .SI(\mem0[108][4] ), .SE(test_se), 
        .CLK(n1679), .Q(\mem0[108][5] ), .QN(n24731) );
  SDFFX1 \mem0_reg[108][4]  ( .D(n17424), .SI(\mem0[108][3] ), .SE(test_se), 
        .CLK(n1679), .Q(\mem0[108][4] ), .QN(n24732) );
  SDFFX1 \mem0_reg[108][3]  ( .D(n17423), .SI(\mem0[108][2] ), .SE(test_se), 
        .CLK(n1679), .Q(\mem0[108][3] ), .QN(n24733) );
  SDFFX1 \mem0_reg[108][2]  ( .D(n17422), .SI(\mem0[108][1] ), .SE(test_se), 
        .CLK(n1679), .Q(\mem0[108][2] ), .QN(n24734) );
  SDFFX1 \mem0_reg[108][1]  ( .D(n17421), .SI(\mem0[108][0] ), .SE(test_se), 
        .CLK(n1679), .Q(\mem0[108][1] ), .QN(n24735) );
  SDFFX1 \mem0_reg[108][0]  ( .D(n17420), .SI(\mem0[107][7] ), .SE(test_se), 
        .CLK(n1679), .Q(\mem0[108][0] ), .QN(n24736) );
  SDFFX1 \mem0_reg[107][7]  ( .D(n17419), .SI(\mem0[107][6] ), .SE(test_se), 
        .CLK(n1679), .Q(\mem0[107][7] ), .QN(n24737) );
  SDFFX1 \mem0_reg[107][6]  ( .D(n17418), .SI(\mem0[107][5] ), .SE(test_se), 
        .CLK(n1679), .Q(\mem0[107][6] ), .QN(n24738) );
  SDFFX1 \mem0_reg[107][5]  ( .D(n17417), .SI(\mem0[107][4] ), .SE(test_se), 
        .CLK(n1680), .Q(\mem0[107][5] ), .QN(n24739) );
  SDFFX1 \mem0_reg[107][4]  ( .D(n17416), .SI(\mem0[107][3] ), .SE(test_se), 
        .CLK(n1680), .Q(\mem0[107][4] ), .QN(n24740) );
  SDFFX1 \mem0_reg[107][3]  ( .D(n17415), .SI(\mem0[107][2] ), .SE(test_se), 
        .CLK(n1680), .Q(\mem0[107][3] ), .QN(n24741) );
  SDFFX1 \mem0_reg[107][2]  ( .D(n17414), .SI(\mem0[107][1] ), .SE(test_se), 
        .CLK(n1680), .Q(\mem0[107][2] ), .QN(n24742) );
  SDFFX1 \mem0_reg[107][1]  ( .D(n17413), .SI(\mem0[107][0] ), .SE(test_se), 
        .CLK(n1680), .Q(\mem0[107][1] ), .QN(n24743) );
  SDFFX1 \mem0_reg[107][0]  ( .D(n17412), .SI(\mem0[106][7] ), .SE(test_se), 
        .CLK(n1680), .Q(\mem0[107][0] ), .QN(n24744) );
  SDFFX1 \mem0_reg[106][7]  ( .D(n17411), .SI(\mem0[106][6] ), .SE(test_se), 
        .CLK(n1680), .Q(\mem0[106][7] ), .QN(n24745) );
  SDFFX1 \mem0_reg[106][6]  ( .D(n17410), .SI(\mem0[106][5] ), .SE(test_se), 
        .CLK(n1680), .Q(\mem0[106][6] ), .QN(n24746) );
  SDFFX1 \mem0_reg[106][5]  ( .D(n17409), .SI(\mem0[106][4] ), .SE(test_se), 
        .CLK(n1680), .Q(\mem0[106][5] ), .QN(n24747) );
  SDFFX1 \mem0_reg[106][4]  ( .D(n17408), .SI(\mem0[106][3] ), .SE(test_se), 
        .CLK(n1680), .Q(\mem0[106][4] ), .QN(n24748) );
  SDFFX1 \mem0_reg[106][3]  ( .D(n17407), .SI(\mem0[106][2] ), .SE(test_se), 
        .CLK(n1680), .Q(\mem0[106][3] ), .QN(n24749) );
  SDFFX1 \mem0_reg[106][2]  ( .D(n17406), .SI(\mem0[106][1] ), .SE(test_se), 
        .CLK(n1680), .Q(\mem0[106][2] ), .QN(n24750) );
  SDFFX1 \mem0_reg[106][1]  ( .D(n17405), .SI(\mem0[106][0] ), .SE(test_se), 
        .CLK(n1681), .Q(\mem0[106][1] ), .QN(n24751) );
  SDFFX1 \mem0_reg[106][0]  ( .D(n17404), .SI(\mem0[105][7] ), .SE(test_se), 
        .CLK(n1681), .Q(\mem0[106][0] ), .QN(n24752) );
  SDFFX1 \mem0_reg[105][7]  ( .D(n17403), .SI(\mem0[105][6] ), .SE(test_se), 
        .CLK(n1681), .Q(\mem0[105][7] ), .QN(n24753) );
  SDFFX1 \mem0_reg[105][6]  ( .D(n17402), .SI(\mem0[105][5] ), .SE(test_se), 
        .CLK(n1681), .Q(\mem0[105][6] ), .QN(n24754) );
  SDFFX1 \mem0_reg[105][5]  ( .D(n17401), .SI(\mem0[105][4] ), .SE(test_se), 
        .CLK(n1681), .Q(\mem0[105][5] ), .QN(n24755) );
  SDFFX1 \mem0_reg[105][4]  ( .D(n17400), .SI(\mem0[105][3] ), .SE(test_se), 
        .CLK(n1681), .Q(\mem0[105][4] ), .QN(n24756) );
  SDFFX1 \mem0_reg[105][3]  ( .D(n17399), .SI(\mem0[105][2] ), .SE(test_se), 
        .CLK(n1681), .Q(\mem0[105][3] ), .QN(n24757) );
  SDFFX1 \mem0_reg[105][2]  ( .D(n17398), .SI(\mem0[105][1] ), .SE(test_se), 
        .CLK(n1681), .Q(\mem0[105][2] ), .QN(n24758) );
  SDFFX1 \mem0_reg[105][1]  ( .D(n17397), .SI(\mem0[105][0] ), .SE(test_se), 
        .CLK(n1681), .Q(\mem0[105][1] ), .QN(n24759) );
  SDFFX1 \mem0_reg[105][0]  ( .D(n17396), .SI(\mem0[104][7] ), .SE(test_se), 
        .CLK(n1681), .Q(\mem0[105][0] ), .QN(n24760) );
  SDFFX1 \mem0_reg[104][7]  ( .D(n17395), .SI(\mem0[104][6] ), .SE(test_se), 
        .CLK(n1681), .Q(\mem0[104][7] ), .QN(n24761) );
  SDFFX1 \mem0_reg[104][6]  ( .D(n17394), .SI(\mem0[104][5] ), .SE(test_se), 
        .CLK(n1681), .Q(\mem0[104][6] ), .QN(n24762) );
  SDFFX1 \mem0_reg[104][5]  ( .D(n17393), .SI(\mem0[104][4] ), .SE(test_se), 
        .CLK(n1682), .Q(\mem0[104][5] ), .QN(n24763) );
  SDFFX1 \mem0_reg[104][4]  ( .D(n17392), .SI(\mem0[104][3] ), .SE(test_se), 
        .CLK(n1682), .Q(\mem0[104][4] ), .QN(n24764) );
  SDFFX1 \mem0_reg[104][3]  ( .D(n17391), .SI(\mem0[104][2] ), .SE(test_se), 
        .CLK(n1682), .Q(\mem0[104][3] ), .QN(n24765) );
  SDFFX1 \mem0_reg[104][2]  ( .D(n17390), .SI(\mem0[104][1] ), .SE(test_se), 
        .CLK(n1682), .Q(\mem0[104][2] ), .QN(n24766) );
  SDFFX1 \mem0_reg[104][1]  ( .D(n17389), .SI(\mem0[104][0] ), .SE(test_se), 
        .CLK(n1682), .Q(\mem0[104][1] ), .QN(n24767) );
  SDFFX1 \mem0_reg[104][0]  ( .D(n17388), .SI(\mem0[103][7] ), .SE(test_se), 
        .CLK(n1682), .Q(\mem0[104][0] ), .QN(n24768) );
  SDFFX1 \mem0_reg[103][7]  ( .D(n17387), .SI(\mem0[103][6] ), .SE(test_se), 
        .CLK(n1682), .Q(\mem0[103][7] ), .QN(n24769) );
  SDFFX1 \mem0_reg[103][6]  ( .D(n17386), .SI(\mem0[103][5] ), .SE(test_se), 
        .CLK(n1682), .Q(\mem0[103][6] ), .QN(n24770) );
  SDFFX1 \mem0_reg[103][5]  ( .D(n17385), .SI(\mem0[103][4] ), .SE(test_se), 
        .CLK(n1682), .Q(\mem0[103][5] ), .QN(n24771) );
  SDFFX1 \mem0_reg[103][4]  ( .D(n17384), .SI(\mem0[103][3] ), .SE(test_se), 
        .CLK(n1682), .Q(\mem0[103][4] ), .QN(n24772) );
  SDFFX1 \mem0_reg[103][3]  ( .D(n17383), .SI(\mem0[103][2] ), .SE(test_se), 
        .CLK(n1682), .Q(\mem0[103][3] ), .QN(n24773) );
  SDFFX1 \mem0_reg[103][2]  ( .D(n17382), .SI(\mem0[103][1] ), .SE(test_se), 
        .CLK(n1682), .Q(\mem0[103][2] ), .QN(n24774) );
  SDFFX1 \mem0_reg[103][1]  ( .D(n17381), .SI(\mem0[103][0] ), .SE(test_se), 
        .CLK(n1683), .Q(\mem0[103][1] ), .QN(n24775) );
  SDFFX1 \mem0_reg[103][0]  ( .D(n17380), .SI(\mem0[102][7] ), .SE(test_se), 
        .CLK(n1683), .Q(\mem0[103][0] ), .QN(n24776) );
  SDFFX1 \mem0_reg[102][7]  ( .D(n17379), .SI(\mem0[102][6] ), .SE(test_se), 
        .CLK(n1683), .Q(\mem0[102][7] ), .QN(n24777) );
  SDFFX1 \mem0_reg[102][6]  ( .D(n17378), .SI(\mem0[102][5] ), .SE(test_se), 
        .CLK(n1683), .Q(\mem0[102][6] ), .QN(n24778) );
  SDFFX1 \mem0_reg[102][5]  ( .D(n17377), .SI(\mem0[102][4] ), .SE(test_se), 
        .CLK(n1683), .Q(\mem0[102][5] ), .QN(n24779) );
  SDFFX1 \mem0_reg[102][4]  ( .D(n17376), .SI(\mem0[102][3] ), .SE(test_se), 
        .CLK(n1683), .Q(\mem0[102][4] ), .QN(n24780) );
  SDFFX1 \mem0_reg[102][3]  ( .D(n17375), .SI(\mem0[102][2] ), .SE(test_se), 
        .CLK(n1683), .Q(\mem0[102][3] ), .QN(n24781) );
  SDFFX1 \mem0_reg[102][2]  ( .D(n17374), .SI(\mem0[102][1] ), .SE(test_se), 
        .CLK(n1683), .Q(\mem0[102][2] ), .QN(n24782) );
  SDFFX1 \mem0_reg[102][1]  ( .D(n17373), .SI(\mem0[102][0] ), .SE(test_se), 
        .CLK(n1683), .Q(\mem0[102][1] ), .QN(n24783) );
  SDFFX1 \mem0_reg[102][0]  ( .D(n17372), .SI(\mem0[101][7] ), .SE(test_se), 
        .CLK(n1683), .Q(\mem0[102][0] ), .QN(n24784) );
  SDFFX1 \mem0_reg[101][7]  ( .D(n17371), .SI(\mem0[101][6] ), .SE(test_se), 
        .CLK(n1683), .Q(\mem0[101][7] ), .QN(n24785) );
  SDFFX1 \mem0_reg[101][6]  ( .D(n17370), .SI(\mem0[101][5] ), .SE(test_se), 
        .CLK(n1683), .Q(\mem0[101][6] ), .QN(n24786) );
  SDFFX1 \mem0_reg[101][5]  ( .D(n17369), .SI(\mem0[101][4] ), .SE(test_se), 
        .CLK(n1684), .Q(\mem0[101][5] ), .QN(n24787) );
  SDFFX1 \mem0_reg[101][4]  ( .D(n17368), .SI(\mem0[101][3] ), .SE(test_se), 
        .CLK(n1684), .Q(\mem0[101][4] ), .QN(n24788) );
  SDFFX1 \mem0_reg[101][3]  ( .D(n17367), .SI(\mem0[101][2] ), .SE(test_se), 
        .CLK(n1684), .Q(\mem0[101][3] ), .QN(n24789) );
  SDFFX1 \mem0_reg[101][2]  ( .D(n17366), .SI(\mem0[101][1] ), .SE(test_se), 
        .CLK(n1684), .Q(\mem0[101][2] ), .QN(n24790) );
  SDFFX1 \mem0_reg[101][1]  ( .D(n17365), .SI(\mem0[101][0] ), .SE(test_se), 
        .CLK(n1684), .Q(\mem0[101][1] ), .QN(n24791) );
  SDFFX1 \mem0_reg[101][0]  ( .D(n17364), .SI(\mem0[100][7] ), .SE(test_se), 
        .CLK(n1684), .Q(\mem0[101][0] ), .QN(n24792) );
  SDFFX1 \mem0_reg[100][7]  ( .D(n17363), .SI(\mem0[100][6] ), .SE(test_se), 
        .CLK(n1684), .Q(\mem0[100][7] ), .QN(n24793) );
  SDFFX1 \mem0_reg[100][6]  ( .D(n17362), .SI(\mem0[100][5] ), .SE(test_se), 
        .CLK(n1684), .Q(\mem0[100][6] ), .QN(n24794) );
  SDFFX1 \mem0_reg[100][5]  ( .D(n17361), .SI(\mem0[100][4] ), .SE(test_se), 
        .CLK(n1684), .Q(\mem0[100][5] ), .QN(n24795) );
  SDFFX1 \mem0_reg[100][4]  ( .D(n17360), .SI(\mem0[100][3] ), .SE(test_se), 
        .CLK(n1684), .Q(\mem0[100][4] ), .QN(n24796) );
  SDFFX1 \mem0_reg[100][3]  ( .D(n17359), .SI(\mem0[100][2] ), .SE(test_se), 
        .CLK(n1684), .Q(\mem0[100][3] ), .QN(n24797) );
  SDFFX1 \mem0_reg[100][2]  ( .D(n17358), .SI(\mem0[100][1] ), .SE(test_se), 
        .CLK(n1684), .Q(\mem0[100][2] ), .QN(n24798) );
  SDFFX1 \mem0_reg[100][1]  ( .D(n17357), .SI(\mem0[100][0] ), .SE(test_se), 
        .CLK(n1685), .Q(\mem0[100][1] ), .QN(n24799) );
  SDFFX1 \mem0_reg[100][0]  ( .D(n17356), .SI(\mem0[99][7] ), .SE(test_se), 
        .CLK(n1685), .Q(\mem0[100][0] ), .QN(n24800) );
  SDFFX1 \mem0_reg[99][7]  ( .D(n17355), .SI(\mem0[99][6] ), .SE(test_se), 
        .CLK(n1685), .Q(\mem0[99][7] ), .QN(n24801) );
  SDFFX1 \mem0_reg[99][6]  ( .D(n17354), .SI(\mem0[99][5] ), .SE(test_se), 
        .CLK(n1685), .Q(\mem0[99][6] ), .QN(n24802) );
  SDFFX1 \mem0_reg[99][5]  ( .D(n17353), .SI(\mem0[99][4] ), .SE(test_se), 
        .CLK(n1685), .Q(\mem0[99][5] ), .QN(n24803) );
  SDFFX1 \mem0_reg[99][4]  ( .D(n17352), .SI(\mem0[99][3] ), .SE(test_se), 
        .CLK(n1685), .Q(\mem0[99][4] ), .QN(n24804) );
  SDFFX1 \mem0_reg[99][3]  ( .D(n17351), .SI(\mem0[99][2] ), .SE(test_se), 
        .CLK(n1685), .Q(\mem0[99][3] ), .QN(n24805) );
  SDFFX1 \mem0_reg[99][2]  ( .D(n17350), .SI(\mem0[99][1] ), .SE(test_se), 
        .CLK(n1685), .Q(\mem0[99][2] ), .QN(n24806) );
  SDFFX1 \mem0_reg[99][1]  ( .D(n17349), .SI(\mem0[99][0] ), .SE(test_se), 
        .CLK(n1685), .Q(\mem0[99][1] ), .QN(n24807) );
  SDFFX1 \mem0_reg[99][0]  ( .D(n17348), .SI(\mem0[98][7] ), .SE(test_se), 
        .CLK(n1685), .Q(\mem0[99][0] ), .QN(n24808) );
  SDFFX1 \mem0_reg[98][7]  ( .D(n17347), .SI(\mem0[98][6] ), .SE(test_se), 
        .CLK(n1685), .Q(\mem0[98][7] ), .QN(n24809) );
  SDFFX1 \mem0_reg[98][6]  ( .D(n17346), .SI(\mem0[98][5] ), .SE(test_se), 
        .CLK(n1685), .Q(\mem0[98][6] ), .QN(n24810) );
  SDFFX1 \mem0_reg[98][5]  ( .D(n17345), .SI(\mem0[98][4] ), .SE(test_se), 
        .CLK(n1686), .Q(\mem0[98][5] ), .QN(n24811) );
  SDFFX1 \mem0_reg[98][4]  ( .D(n17344), .SI(\mem0[98][3] ), .SE(test_se), 
        .CLK(n1686), .Q(\mem0[98][4] ), .QN(n24812) );
  SDFFX1 \mem0_reg[98][3]  ( .D(n17343), .SI(\mem0[98][2] ), .SE(test_se), 
        .CLK(n1686), .Q(\mem0[98][3] ), .QN(n24813) );
  SDFFX1 \mem0_reg[98][2]  ( .D(n17342), .SI(\mem0[98][1] ), .SE(test_se), 
        .CLK(n1686), .Q(\mem0[98][2] ), .QN(n24814) );
  SDFFX1 \mem0_reg[98][1]  ( .D(n17341), .SI(\mem0[98][0] ), .SE(test_se), 
        .CLK(n1686), .Q(\mem0[98][1] ), .QN(n24815) );
  SDFFX1 \mem0_reg[98][0]  ( .D(n17340), .SI(\mem0[97][7] ), .SE(test_se), 
        .CLK(n1686), .Q(\mem0[98][0] ), .QN(n24816) );
  SDFFX1 \mem0_reg[97][7]  ( .D(n17339), .SI(\mem0[97][6] ), .SE(test_se), 
        .CLK(n1686), .Q(\mem0[97][7] ), .QN(n24817) );
  SDFFX1 \mem0_reg[97][6]  ( .D(n17338), .SI(\mem0[97][5] ), .SE(test_se), 
        .CLK(n1686), .Q(\mem0[97][6] ), .QN(n24818) );
  SDFFX1 \mem0_reg[97][5]  ( .D(n17337), .SI(\mem0[97][4] ), .SE(test_se), 
        .CLK(n1686), .Q(\mem0[97][5] ), .QN(n24819) );
  SDFFX1 \mem0_reg[97][4]  ( .D(n17336), .SI(\mem0[97][3] ), .SE(test_se), 
        .CLK(n1686), .Q(\mem0[97][4] ), .QN(n24820) );
  SDFFX1 \mem0_reg[97][3]  ( .D(n17335), .SI(\mem0[97][2] ), .SE(test_se), 
        .CLK(n1686), .Q(\mem0[97][3] ), .QN(n24821) );
  SDFFX1 \mem0_reg[97][2]  ( .D(n17334), .SI(\mem0[97][1] ), .SE(test_se), 
        .CLK(n1686), .Q(\mem0[97][2] ), .QN(n24822) );
  SDFFX1 \mem0_reg[97][1]  ( .D(n17333), .SI(\mem0[97][0] ), .SE(test_se), 
        .CLK(n1687), .Q(\mem0[97][1] ), .QN(n24823) );
  SDFFX1 \mem0_reg[97][0]  ( .D(n17332), .SI(\mem0[96][7] ), .SE(test_se), 
        .CLK(n1687), .Q(\mem0[97][0] ), .QN(n24824) );
  SDFFX1 \mem0_reg[96][7]  ( .D(n17331), .SI(\mem0[96][6] ), .SE(test_se), 
        .CLK(n1687), .Q(\mem0[96][7] ), .QN(n24825) );
  SDFFX1 \mem0_reg[96][6]  ( .D(n17330), .SI(\mem0[96][5] ), .SE(test_se), 
        .CLK(n1687), .Q(\mem0[96][6] ), .QN(n24826) );
  SDFFX1 \mem0_reg[96][5]  ( .D(n17329), .SI(\mem0[96][4] ), .SE(test_se), 
        .CLK(n1687), .Q(\mem0[96][5] ), .QN(n24827) );
  SDFFX1 \mem0_reg[96][4]  ( .D(n17328), .SI(\mem0[96][3] ), .SE(test_se), 
        .CLK(n1687), .Q(\mem0[96][4] ), .QN(n24828) );
  SDFFX1 \mem0_reg[96][3]  ( .D(n17327), .SI(\mem0[96][2] ), .SE(test_se), 
        .CLK(n1687), .Q(\mem0[96][3] ), .QN(n24829) );
  SDFFX1 \mem0_reg[96][2]  ( .D(n17326), .SI(\mem0[96][1] ), .SE(test_se), 
        .CLK(n1687), .Q(\mem0[96][2] ), .QN(n24830) );
  SDFFX1 \mem0_reg[96][1]  ( .D(n17325), .SI(\mem0[96][0] ), .SE(test_se), 
        .CLK(n1687), .Q(\mem0[96][1] ), .QN(n24831) );
  SDFFX1 \mem0_reg[96][0]  ( .D(n17324), .SI(\mem0[95][7] ), .SE(test_se), 
        .CLK(n1687), .Q(\mem0[96][0] ), .QN(n24832) );
  SDFFX1 \mem0_reg[95][7]  ( .D(n17323), .SI(\mem0[95][6] ), .SE(test_se), 
        .CLK(n1687), .Q(\mem0[95][7] ), .QN(n24833) );
  SDFFX1 \mem0_reg[95][6]  ( .D(n17322), .SI(\mem0[95][5] ), .SE(test_se), 
        .CLK(n1687), .Q(\mem0[95][6] ), .QN(n24834) );
  SDFFX1 \mem0_reg[95][5]  ( .D(n17321), .SI(\mem0[95][4] ), .SE(test_se), 
        .CLK(n1688), .Q(\mem0[95][5] ), .QN(n24835) );
  SDFFX1 \mem0_reg[95][4]  ( .D(n17320), .SI(\mem0[95][3] ), .SE(test_se), 
        .CLK(n1688), .Q(\mem0[95][4] ), .QN(n24836) );
  SDFFX1 \mem0_reg[95][3]  ( .D(n17319), .SI(\mem0[95][2] ), .SE(test_se), 
        .CLK(n1688), .Q(\mem0[95][3] ), .QN(n24837) );
  SDFFX1 \mem0_reg[95][2]  ( .D(n17318), .SI(\mem0[95][1] ), .SE(test_se), 
        .CLK(n1688), .Q(\mem0[95][2] ), .QN(n24838) );
  SDFFX1 \mem0_reg[95][1]  ( .D(n17317), .SI(\mem0[95][0] ), .SE(test_se), 
        .CLK(n1688), .Q(\mem0[95][1] ), .QN(n24839) );
  SDFFX1 \mem0_reg[95][0]  ( .D(n17316), .SI(\mem0[94][7] ), .SE(test_se), 
        .CLK(n1688), .Q(\mem0[95][0] ), .QN(n24840) );
  SDFFX1 \mem0_reg[94][7]  ( .D(n17315), .SI(\mem0[94][6] ), .SE(test_se), 
        .CLK(n1688), .Q(\mem0[94][7] ), .QN(n24841) );
  SDFFX1 \mem0_reg[94][6]  ( .D(n17314), .SI(\mem0[94][5] ), .SE(test_se), 
        .CLK(n1688), .Q(\mem0[94][6] ), .QN(n24842) );
  SDFFX1 \mem0_reg[94][5]  ( .D(n17313), .SI(\mem0[94][4] ), .SE(test_se), 
        .CLK(n1688), .Q(\mem0[94][5] ), .QN(n24843) );
  SDFFX1 \mem0_reg[94][4]  ( .D(n17312), .SI(\mem0[94][3] ), .SE(test_se), 
        .CLK(n1688), .Q(\mem0[94][4] ), .QN(n24844) );
  SDFFX1 \mem0_reg[94][3]  ( .D(n17311), .SI(\mem0[94][2] ), .SE(test_se), 
        .CLK(n1688), .Q(\mem0[94][3] ), .QN(n24845) );
  SDFFX1 \mem0_reg[94][2]  ( .D(n17310), .SI(\mem0[94][1] ), .SE(test_se), 
        .CLK(n1688), .Q(\mem0[94][2] ), .QN(n24846) );
  SDFFX1 \mem0_reg[94][1]  ( .D(n17309), .SI(\mem0[94][0] ), .SE(test_se), 
        .CLK(n1689), .Q(\mem0[94][1] ), .QN(n24847) );
  SDFFX1 \mem0_reg[94][0]  ( .D(n17308), .SI(\mem0[93][7] ), .SE(test_se), 
        .CLK(n1689), .Q(\mem0[94][0] ), .QN(n24848) );
  SDFFX1 \mem0_reg[93][7]  ( .D(n17307), .SI(\mem0[93][6] ), .SE(test_se), 
        .CLK(n1689), .Q(\mem0[93][7] ), .QN(n24849) );
  SDFFX1 \mem0_reg[93][6]  ( .D(n17306), .SI(\mem0[93][5] ), .SE(test_se), 
        .CLK(n1689), .Q(\mem0[93][6] ), .QN(n24850) );
  SDFFX1 \mem0_reg[93][5]  ( .D(n17305), .SI(\mem0[93][4] ), .SE(test_se), 
        .CLK(n1689), .Q(\mem0[93][5] ), .QN(n24851) );
  SDFFX1 \mem0_reg[93][4]  ( .D(n17304), .SI(\mem0[93][3] ), .SE(test_se), 
        .CLK(n1689), .Q(\mem0[93][4] ), .QN(n24852) );
  SDFFX1 \mem0_reg[93][3]  ( .D(n17303), .SI(\mem0[93][2] ), .SE(test_se), 
        .CLK(n1689), .Q(\mem0[93][3] ), .QN(n24853) );
  SDFFX1 \mem0_reg[93][2]  ( .D(n17302), .SI(\mem0[93][1] ), .SE(test_se), 
        .CLK(n1689), .Q(\mem0[93][2] ), .QN(n24854) );
  SDFFX1 \mem0_reg[93][1]  ( .D(n17301), .SI(\mem0[93][0] ), .SE(test_se), 
        .CLK(n1689), .Q(\mem0[93][1] ), .QN(n24855) );
  SDFFX1 \mem0_reg[93][0]  ( .D(n17300), .SI(\mem0[92][7] ), .SE(test_se), 
        .CLK(n1689), .Q(\mem0[93][0] ), .QN(n24856) );
  SDFFX1 \mem0_reg[92][7]  ( .D(n17299), .SI(\mem0[92][6] ), .SE(test_se), 
        .CLK(n1689), .Q(\mem0[92][7] ), .QN(n24857) );
  SDFFX1 \mem0_reg[92][6]  ( .D(n17298), .SI(\mem0[92][5] ), .SE(test_se), 
        .CLK(n1689), .Q(\mem0[92][6] ), .QN(n24858) );
  SDFFX1 \mem0_reg[92][5]  ( .D(n17297), .SI(\mem0[92][4] ), .SE(test_se), 
        .CLK(n1690), .Q(\mem0[92][5] ), .QN(n24859) );
  SDFFX1 \mem0_reg[92][4]  ( .D(n17296), .SI(\mem0[92][3] ), .SE(test_se), 
        .CLK(n1690), .Q(\mem0[92][4] ), .QN(n24860) );
  SDFFX1 \mem0_reg[92][3]  ( .D(n17295), .SI(\mem0[92][2] ), .SE(test_se), 
        .CLK(n1690), .Q(\mem0[92][3] ), .QN(n24861) );
  SDFFX1 \mem0_reg[92][2]  ( .D(n17294), .SI(\mem0[92][1] ), .SE(test_se), 
        .CLK(n1690), .Q(\mem0[92][2] ), .QN(n24862) );
  SDFFX1 \mem0_reg[92][1]  ( .D(n17293), .SI(\mem0[92][0] ), .SE(test_se), 
        .CLK(n1690), .Q(\mem0[92][1] ), .QN(n24863) );
  SDFFX1 \mem0_reg[92][0]  ( .D(n17292), .SI(\mem0[91][7] ), .SE(test_se), 
        .CLK(n1690), .Q(\mem0[92][0] ), .QN(n24864) );
  SDFFX1 \mem0_reg[91][7]  ( .D(n17291), .SI(\mem0[91][6] ), .SE(test_se), 
        .CLK(n1690), .Q(\mem0[91][7] ), .QN(n24865) );
  SDFFX1 \mem0_reg[91][6]  ( .D(n17290), .SI(\mem0[91][5] ), .SE(test_se), 
        .CLK(n1690), .Q(\mem0[91][6] ), .QN(n24866) );
  SDFFX1 \mem0_reg[91][5]  ( .D(n17289), .SI(\mem0[91][4] ), .SE(test_se), 
        .CLK(n1690), .Q(\mem0[91][5] ), .QN(n24867) );
  SDFFX1 \mem0_reg[91][4]  ( .D(n17288), .SI(\mem0[91][3] ), .SE(test_se), 
        .CLK(n1690), .Q(\mem0[91][4] ), .QN(n24868) );
  SDFFX1 \mem0_reg[91][3]  ( .D(n17287), .SI(\mem0[91][2] ), .SE(test_se), 
        .CLK(n1690), .Q(\mem0[91][3] ), .QN(n24869) );
  SDFFX1 \mem0_reg[91][2]  ( .D(n17286), .SI(\mem0[91][1] ), .SE(test_se), 
        .CLK(n1690), .Q(\mem0[91][2] ), .QN(n24870) );
  SDFFX1 \mem0_reg[91][1]  ( .D(n17285), .SI(\mem0[91][0] ), .SE(test_se), 
        .CLK(n1691), .Q(\mem0[91][1] ), .QN(n24871) );
  SDFFX1 \mem0_reg[91][0]  ( .D(n17284), .SI(\mem0[90][7] ), .SE(test_se), 
        .CLK(n1691), .Q(\mem0[91][0] ), .QN(n24872) );
  SDFFX1 \mem0_reg[90][7]  ( .D(n17283), .SI(\mem0[90][6] ), .SE(test_se), 
        .CLK(n1691), .Q(\mem0[90][7] ), .QN(n24873) );
  SDFFX1 \mem0_reg[90][6]  ( .D(n17282), .SI(\mem0[90][5] ), .SE(test_se), 
        .CLK(n1691), .Q(\mem0[90][6] ), .QN(n24874) );
  SDFFX1 \mem0_reg[90][5]  ( .D(n17281), .SI(\mem0[90][4] ), .SE(test_se), 
        .CLK(n1691), .Q(\mem0[90][5] ), .QN(n24875) );
  SDFFX1 \mem0_reg[90][4]  ( .D(n17280), .SI(\mem0[90][3] ), .SE(test_se), 
        .CLK(n1691), .Q(\mem0[90][4] ), .QN(n24876) );
  SDFFX1 \mem0_reg[90][3]  ( .D(n17279), .SI(\mem0[90][2] ), .SE(test_se), 
        .CLK(n1691), .Q(\mem0[90][3] ), .QN(n24877) );
  SDFFX1 \mem0_reg[90][2]  ( .D(n17278), .SI(\mem0[90][1] ), .SE(test_se), 
        .CLK(n1691), .Q(\mem0[90][2] ), .QN(n24878) );
  SDFFX1 \mem0_reg[90][1]  ( .D(n17277), .SI(\mem0[90][0] ), .SE(test_se), 
        .CLK(n1691), .Q(\mem0[90][1] ), .QN(n24879) );
  SDFFX1 \mem0_reg[90][0]  ( .D(n17276), .SI(\mem0[89][7] ), .SE(test_se), 
        .CLK(n1691), .Q(\mem0[90][0] ), .QN(n24880) );
  SDFFX1 \mem0_reg[89][7]  ( .D(n17275), .SI(\mem0[89][6] ), .SE(test_se), 
        .CLK(n1691), .Q(\mem0[89][7] ), .QN(n24881) );
  SDFFX1 \mem0_reg[89][6]  ( .D(n17274), .SI(\mem0[89][5] ), .SE(test_se), 
        .CLK(n1691), .Q(\mem0[89][6] ), .QN(n24882) );
  SDFFX1 \mem0_reg[89][5]  ( .D(n17273), .SI(\mem0[89][4] ), .SE(test_se), 
        .CLK(n1692), .Q(\mem0[89][5] ), .QN(n24883) );
  SDFFX1 \mem0_reg[89][4]  ( .D(n17272), .SI(\mem0[89][3] ), .SE(test_se), 
        .CLK(n1692), .Q(\mem0[89][4] ), .QN(n24884) );
  SDFFX1 \mem0_reg[89][3]  ( .D(n17271), .SI(\mem0[89][2] ), .SE(test_se), 
        .CLK(n1692), .Q(\mem0[89][3] ), .QN(n24885) );
  SDFFX1 \mem0_reg[89][2]  ( .D(n17270), .SI(\mem0[89][1] ), .SE(test_se), 
        .CLK(n1692), .Q(\mem0[89][2] ), .QN(n24886) );
  SDFFX1 \mem0_reg[89][1]  ( .D(n17269), .SI(\mem0[89][0] ), .SE(test_se), 
        .CLK(n1692), .Q(\mem0[89][1] ), .QN(n24887) );
  SDFFX1 \mem0_reg[89][0]  ( .D(n17268), .SI(\mem0[88][7] ), .SE(test_se), 
        .CLK(n1692), .Q(\mem0[89][0] ), .QN(n24888) );
  SDFFX1 \mem0_reg[88][7]  ( .D(n17267), .SI(\mem0[88][6] ), .SE(test_se), 
        .CLK(n1692), .Q(\mem0[88][7] ), .QN(n24889) );
  SDFFX1 \mem0_reg[88][6]  ( .D(n17266), .SI(\mem0[88][5] ), .SE(test_se), 
        .CLK(n1692), .Q(\mem0[88][6] ), .QN(n24890) );
  SDFFX1 \mem0_reg[88][5]  ( .D(n17265), .SI(\mem0[88][4] ), .SE(test_se), 
        .CLK(n1692), .Q(\mem0[88][5] ), .QN(n24891) );
  SDFFX1 \mem0_reg[88][4]  ( .D(n17264), .SI(\mem0[88][3] ), .SE(test_se), 
        .CLK(n1692), .Q(\mem0[88][4] ), .QN(n24892) );
  SDFFX1 \mem0_reg[88][3]  ( .D(n17263), .SI(\mem0[88][2] ), .SE(test_se), 
        .CLK(n1692), .Q(\mem0[88][3] ), .QN(n24893) );
  SDFFX1 \mem0_reg[88][2]  ( .D(n17262), .SI(\mem0[88][1] ), .SE(test_se), 
        .CLK(n1692), .Q(\mem0[88][2] ), .QN(n24894) );
  SDFFX1 \mem0_reg[88][1]  ( .D(n17261), .SI(\mem0[88][0] ), .SE(test_se), 
        .CLK(n1693), .Q(\mem0[88][1] ), .QN(n24895) );
  SDFFX1 \mem0_reg[88][0]  ( .D(n17260), .SI(\mem0[87][7] ), .SE(test_se), 
        .CLK(n1693), .Q(\mem0[88][0] ), .QN(n24896) );
  SDFFX1 \mem0_reg[87][7]  ( .D(n17259), .SI(\mem0[87][6] ), .SE(test_se), 
        .CLK(n1693), .Q(\mem0[87][7] ), .QN(n24897) );
  SDFFX1 \mem0_reg[87][6]  ( .D(n17258), .SI(\mem0[87][5] ), .SE(test_se), 
        .CLK(n1693), .Q(\mem0[87][6] ), .QN(n24898) );
  SDFFX1 \mem0_reg[87][5]  ( .D(n17257), .SI(\mem0[87][4] ), .SE(test_se), 
        .CLK(n1693), .Q(\mem0[87][5] ), .QN(n24899) );
  SDFFX1 \mem0_reg[87][4]  ( .D(n17256), .SI(\mem0[87][3] ), .SE(test_se), 
        .CLK(n1693), .Q(\mem0[87][4] ), .QN(n24900) );
  SDFFX1 \mem0_reg[87][3]  ( .D(n17255), .SI(\mem0[87][2] ), .SE(test_se), 
        .CLK(n1693), .Q(\mem0[87][3] ), .QN(n24901) );
  SDFFX1 \mem0_reg[87][2]  ( .D(n17254), .SI(\mem0[87][1] ), .SE(test_se), 
        .CLK(n1693), .Q(\mem0[87][2] ), .QN(n24902) );
  SDFFX1 \mem0_reg[87][1]  ( .D(n17253), .SI(\mem0[87][0] ), .SE(test_se), 
        .CLK(n1693), .Q(\mem0[87][1] ), .QN(n24903) );
  SDFFX1 \mem0_reg[87][0]  ( .D(n17252), .SI(\mem0[86][7] ), .SE(test_se), 
        .CLK(n1693), .Q(\mem0[87][0] ), .QN(n24904) );
  SDFFX1 \mem0_reg[86][7]  ( .D(n17251), .SI(\mem0[86][6] ), .SE(test_se), 
        .CLK(n1693), .Q(\mem0[86][7] ), .QN(n24905) );
  SDFFX1 \mem0_reg[86][6]  ( .D(n17250), .SI(\mem0[86][5] ), .SE(test_se), 
        .CLK(n1693), .Q(\mem0[86][6] ), .QN(n24906) );
  SDFFX1 \mem0_reg[86][5]  ( .D(n17249), .SI(\mem0[86][4] ), .SE(test_se), 
        .CLK(n1694), .Q(\mem0[86][5] ), .QN(n24907) );
  SDFFX1 \mem0_reg[86][4]  ( .D(n17248), .SI(\mem0[86][3] ), .SE(test_se), 
        .CLK(n1694), .Q(\mem0[86][4] ), .QN(n24908) );
  SDFFX1 \mem0_reg[86][3]  ( .D(n17247), .SI(\mem0[86][2] ), .SE(test_se), 
        .CLK(n1694), .Q(\mem0[86][3] ), .QN(n24909) );
  SDFFX1 \mem0_reg[86][2]  ( .D(n17246), .SI(\mem0[86][1] ), .SE(test_se), 
        .CLK(n1694), .Q(\mem0[86][2] ), .QN(n24910) );
  SDFFX1 \mem0_reg[86][1]  ( .D(n17245), .SI(\mem0[86][0] ), .SE(test_se), 
        .CLK(n1694), .Q(\mem0[86][1] ), .QN(n24911) );
  SDFFX1 \mem0_reg[86][0]  ( .D(n17244), .SI(\mem0[85][7] ), .SE(test_se), 
        .CLK(n1694), .Q(\mem0[86][0] ), .QN(n24912) );
  SDFFX1 \mem0_reg[85][7]  ( .D(n17243), .SI(\mem0[85][6] ), .SE(test_se), 
        .CLK(n1694), .Q(\mem0[85][7] ), .QN(n24913) );
  SDFFX1 \mem0_reg[85][6]  ( .D(n17242), .SI(\mem0[85][5] ), .SE(test_se), 
        .CLK(n1694), .Q(\mem0[85][6] ), .QN(n24914) );
  SDFFX1 \mem0_reg[85][5]  ( .D(n17241), .SI(\mem0[85][4] ), .SE(test_se), 
        .CLK(n1694), .Q(\mem0[85][5] ), .QN(n24915) );
  SDFFX1 \mem0_reg[85][4]  ( .D(n17240), .SI(\mem0[85][3] ), .SE(test_se), 
        .CLK(n1694), .Q(\mem0[85][4] ), .QN(n24916) );
  SDFFX1 \mem0_reg[85][3]  ( .D(n17239), .SI(\mem0[85][2] ), .SE(test_se), 
        .CLK(n1694), .Q(\mem0[85][3] ), .QN(n24917) );
  SDFFX1 \mem0_reg[85][2]  ( .D(n17238), .SI(\mem0[85][1] ), .SE(test_se), 
        .CLK(n1694), .Q(\mem0[85][2] ), .QN(n24918) );
  SDFFX1 \mem0_reg[85][1]  ( .D(n17237), .SI(\mem0[85][0] ), .SE(test_se), 
        .CLK(n1695), .Q(\mem0[85][1] ), .QN(n24919) );
  SDFFX1 \mem0_reg[85][0]  ( .D(n17236), .SI(\mem0[84][7] ), .SE(test_se), 
        .CLK(n1695), .Q(\mem0[85][0] ), .QN(n24920) );
  SDFFX1 \mem0_reg[84][7]  ( .D(n17235), .SI(\mem0[84][6] ), .SE(test_se), 
        .CLK(n1695), .Q(\mem0[84][7] ), .QN(n24921) );
  SDFFX1 \mem0_reg[84][6]  ( .D(n17234), .SI(\mem0[84][5] ), .SE(test_se), 
        .CLK(n1695), .Q(\mem0[84][6] ), .QN(n24922) );
  SDFFX1 \mem0_reg[84][5]  ( .D(n17233), .SI(\mem0[84][4] ), .SE(test_se), 
        .CLK(n1695), .Q(\mem0[84][5] ), .QN(n24923) );
  SDFFX1 \mem0_reg[84][4]  ( .D(n17232), .SI(\mem0[84][3] ), .SE(test_se), 
        .CLK(n1695), .Q(\mem0[84][4] ), .QN(n24924) );
  SDFFX1 \mem0_reg[84][3]  ( .D(n17231), .SI(\mem0[84][2] ), .SE(test_se), 
        .CLK(n1695), .Q(\mem0[84][3] ), .QN(n24925) );
  SDFFX1 \mem0_reg[84][2]  ( .D(n17230), .SI(\mem0[84][1] ), .SE(test_se), 
        .CLK(n1695), .Q(\mem0[84][2] ), .QN(n24926) );
  SDFFX1 \mem0_reg[84][1]  ( .D(n17229), .SI(\mem0[84][0] ), .SE(test_se), 
        .CLK(n1695), .Q(\mem0[84][1] ), .QN(n24927) );
  SDFFX1 \mem0_reg[84][0]  ( .D(n17228), .SI(\mem0[83][7] ), .SE(test_se), 
        .CLK(n1695), .Q(\mem0[84][0] ), .QN(n24928) );
  SDFFX1 \mem0_reg[83][7]  ( .D(n17227), .SI(\mem0[83][6] ), .SE(test_se), 
        .CLK(n1695), .Q(\mem0[83][7] ), .QN(n24929) );
  SDFFX1 \mem0_reg[83][6]  ( .D(n17226), .SI(\mem0[83][5] ), .SE(test_se), 
        .CLK(n1695), .Q(\mem0[83][6] ), .QN(n24930) );
  SDFFX1 \mem0_reg[83][5]  ( .D(n17225), .SI(\mem0[83][4] ), .SE(test_se), 
        .CLK(n1696), .Q(\mem0[83][5] ), .QN(n24931) );
  SDFFX1 \mem0_reg[83][4]  ( .D(n17224), .SI(\mem0[83][3] ), .SE(test_se), 
        .CLK(n1696), .Q(\mem0[83][4] ), .QN(n24932) );
  SDFFX1 \mem0_reg[83][3]  ( .D(n17223), .SI(\mem0[83][2] ), .SE(test_se), 
        .CLK(n1696), .Q(\mem0[83][3] ), .QN(n24933) );
  SDFFX1 \mem0_reg[83][2]  ( .D(n17222), .SI(\mem0[83][1] ), .SE(test_se), 
        .CLK(n1696), .Q(\mem0[83][2] ), .QN(n24934) );
  SDFFX1 \mem0_reg[83][1]  ( .D(n17221), .SI(\mem0[83][0] ), .SE(test_se), 
        .CLK(n1696), .Q(\mem0[83][1] ), .QN(n24935) );
  SDFFX1 \mem0_reg[83][0]  ( .D(n17220), .SI(\mem0[82][7] ), .SE(test_se), 
        .CLK(n1696), .Q(\mem0[83][0] ), .QN(n24936) );
  SDFFX1 \mem0_reg[82][7]  ( .D(n17219), .SI(\mem0[82][6] ), .SE(test_se), 
        .CLK(n1696), .Q(\mem0[82][7] ), .QN(n24937) );
  SDFFX1 \mem0_reg[82][6]  ( .D(n17218), .SI(\mem0[82][5] ), .SE(test_se), 
        .CLK(n1696), .Q(\mem0[82][6] ), .QN(n24938) );
  SDFFX1 \mem0_reg[82][5]  ( .D(n17217), .SI(\mem0[82][4] ), .SE(test_se), 
        .CLK(n1696), .Q(\mem0[82][5] ), .QN(n24939) );
  SDFFX1 \mem0_reg[82][4]  ( .D(n17216), .SI(\mem0[82][3] ), .SE(test_se), 
        .CLK(n1696), .Q(\mem0[82][4] ), .QN(n24940) );
  SDFFX1 \mem0_reg[82][3]  ( .D(n17215), .SI(\mem0[82][2] ), .SE(test_se), 
        .CLK(n1696), .Q(\mem0[82][3] ), .QN(n24941) );
  SDFFX1 \mem0_reg[82][2]  ( .D(n17214), .SI(\mem0[82][1] ), .SE(test_se), 
        .CLK(n1696), .Q(\mem0[82][2] ), .QN(n24942) );
  SDFFX1 \mem0_reg[82][1]  ( .D(n17213), .SI(\mem0[82][0] ), .SE(test_se), 
        .CLK(n1697), .Q(\mem0[82][1] ), .QN(n24943) );
  SDFFX1 \mem0_reg[82][0]  ( .D(n17212), .SI(\mem0[81][7] ), .SE(test_se), 
        .CLK(n1697), .Q(\mem0[82][0] ), .QN(n24944) );
  SDFFX1 \mem0_reg[81][7]  ( .D(n17211), .SI(\mem0[81][6] ), .SE(test_se), 
        .CLK(n1697), .Q(\mem0[81][7] ), .QN(n24945) );
  SDFFX1 \mem0_reg[81][6]  ( .D(n17210), .SI(\mem0[81][5] ), .SE(test_se), 
        .CLK(n1697), .Q(\mem0[81][6] ), .QN(n24946) );
  SDFFX1 \mem0_reg[81][5]  ( .D(n17209), .SI(\mem0[81][4] ), .SE(test_se), 
        .CLK(n1697), .Q(\mem0[81][5] ), .QN(n24947) );
  SDFFX1 \mem0_reg[81][4]  ( .D(n17208), .SI(\mem0[81][3] ), .SE(test_se), 
        .CLK(n1697), .Q(\mem0[81][4] ), .QN(n24948) );
  SDFFX1 \mem0_reg[81][3]  ( .D(n17207), .SI(\mem0[81][2] ), .SE(test_se), 
        .CLK(n1697), .Q(\mem0[81][3] ), .QN(n24949) );
  SDFFX1 \mem0_reg[81][2]  ( .D(n17206), .SI(\mem0[81][1] ), .SE(test_se), 
        .CLK(n1697), .Q(\mem0[81][2] ), .QN(n24950) );
  SDFFX1 \mem0_reg[81][1]  ( .D(n17205), .SI(\mem0[81][0] ), .SE(test_se), 
        .CLK(n1697), .Q(\mem0[81][1] ), .QN(n24951) );
  SDFFX1 \mem0_reg[81][0]  ( .D(n17204), .SI(\mem0[80][7] ), .SE(test_se), 
        .CLK(n1697), .Q(\mem0[81][0] ), .QN(n24952) );
  SDFFX1 \mem0_reg[80][7]  ( .D(n17203), .SI(\mem0[80][6] ), .SE(test_se), 
        .CLK(n1697), .Q(\mem0[80][7] ), .QN(n24953) );
  SDFFX1 \mem0_reg[80][6]  ( .D(n17202), .SI(\mem0[80][5] ), .SE(test_se), 
        .CLK(n1697), .Q(\mem0[80][6] ), .QN(n24954) );
  SDFFX1 \mem0_reg[80][5]  ( .D(n17201), .SI(\mem0[80][4] ), .SE(test_se), 
        .CLK(n1698), .Q(\mem0[80][5] ), .QN(n24955) );
  SDFFX1 \mem0_reg[80][4]  ( .D(n17200), .SI(\mem0[80][3] ), .SE(test_se), 
        .CLK(n1698), .Q(\mem0[80][4] ), .QN(n24956) );
  SDFFX1 \mem0_reg[80][3]  ( .D(n17199), .SI(\mem0[80][2] ), .SE(test_se), 
        .CLK(n1698), .Q(\mem0[80][3] ), .QN(n24957) );
  SDFFX1 \mem0_reg[80][2]  ( .D(n17198), .SI(\mem0[80][1] ), .SE(test_se), 
        .CLK(n1698), .Q(\mem0[80][2] ), .QN(n24958) );
  SDFFX1 \mem0_reg[80][1]  ( .D(n17197), .SI(\mem0[80][0] ), .SE(test_se), 
        .CLK(n1698), .Q(\mem0[80][1] ), .QN(n24959) );
  SDFFX1 \mem0_reg[80][0]  ( .D(n17196), .SI(\mem0[79][7] ), .SE(test_se), 
        .CLK(n1698), .Q(\mem0[80][0] ), .QN(n24960) );
  SDFFX1 \mem0_reg[79][7]  ( .D(n17195), .SI(\mem0[79][6] ), .SE(test_se), 
        .CLK(n1698), .Q(\mem0[79][7] ), .QN(n24961) );
  SDFFX1 \mem0_reg[79][6]  ( .D(n17194), .SI(\mem0[79][5] ), .SE(test_se), 
        .CLK(n1698), .Q(\mem0[79][6] ), .QN(n24962) );
  SDFFX1 \mem0_reg[79][5]  ( .D(n17193), .SI(\mem0[79][4] ), .SE(test_se), 
        .CLK(n1698), .Q(\mem0[79][5] ), .QN(n24963) );
  SDFFX1 \mem0_reg[79][4]  ( .D(n17192), .SI(\mem0[79][3] ), .SE(test_se), 
        .CLK(n1698), .Q(\mem0[79][4] ), .QN(n24964) );
  SDFFX1 \mem0_reg[79][3]  ( .D(n17191), .SI(\mem0[79][2] ), .SE(test_se), 
        .CLK(n1698), .Q(\mem0[79][3] ), .QN(n24965) );
  SDFFX1 \mem0_reg[79][2]  ( .D(n17190), .SI(\mem0[79][1] ), .SE(test_se), 
        .CLK(n1698), .Q(\mem0[79][2] ), .QN(n24966) );
  SDFFX1 \mem0_reg[79][1]  ( .D(n17189), .SI(\mem0[79][0] ), .SE(test_se), 
        .CLK(n1699), .Q(\mem0[79][1] ), .QN(n24967) );
  SDFFX1 \mem0_reg[79][0]  ( .D(n17188), .SI(\mem0[78][7] ), .SE(test_se), 
        .CLK(n1699), .Q(\mem0[79][0] ), .QN(n24968) );
  SDFFX1 \mem0_reg[78][7]  ( .D(n17187), .SI(\mem0[78][6] ), .SE(test_se), 
        .CLK(n1699), .Q(\mem0[78][7] ), .QN(n24969) );
  SDFFX1 \mem0_reg[78][6]  ( .D(n17186), .SI(\mem0[78][5] ), .SE(test_se), 
        .CLK(n1699), .Q(\mem0[78][6] ), .QN(n24970) );
  SDFFX1 \mem0_reg[78][5]  ( .D(n17185), .SI(\mem0[78][4] ), .SE(test_se), 
        .CLK(n1699), .Q(\mem0[78][5] ), .QN(n24971) );
  SDFFX1 \mem0_reg[78][4]  ( .D(n17184), .SI(\mem0[78][3] ), .SE(test_se), 
        .CLK(n1699), .Q(\mem0[78][4] ), .QN(n24972) );
  SDFFX1 \mem0_reg[78][3]  ( .D(n17183), .SI(\mem0[78][2] ), .SE(test_se), 
        .CLK(n1699), .Q(\mem0[78][3] ), .QN(n24973) );
  SDFFX1 \mem0_reg[78][2]  ( .D(n17182), .SI(\mem0[78][1] ), .SE(test_se), 
        .CLK(n1699), .Q(\mem0[78][2] ), .QN(n24974) );
  SDFFX1 \mem0_reg[78][1]  ( .D(n17181), .SI(\mem0[78][0] ), .SE(test_se), 
        .CLK(n1699), .Q(\mem0[78][1] ), .QN(n24975) );
  SDFFX1 \mem0_reg[78][0]  ( .D(n17180), .SI(\mem0[77][7] ), .SE(test_se), 
        .CLK(n1699), .Q(\mem0[78][0] ), .QN(n24976) );
  SDFFX1 \mem0_reg[77][7]  ( .D(n17179), .SI(\mem0[77][6] ), .SE(test_se), 
        .CLK(n1699), .Q(\mem0[77][7] ), .QN(n24977) );
  SDFFX1 \mem0_reg[77][6]  ( .D(n17178), .SI(\mem0[77][5] ), .SE(test_se), 
        .CLK(n1699), .Q(\mem0[77][6] ), .QN(n24978) );
  SDFFX1 \mem0_reg[77][5]  ( .D(n17177), .SI(\mem0[77][4] ), .SE(test_se), 
        .CLK(n1700), .Q(\mem0[77][5] ), .QN(n24979) );
  SDFFX1 \mem0_reg[77][4]  ( .D(n17176), .SI(\mem0[77][3] ), .SE(test_se), 
        .CLK(n1700), .Q(\mem0[77][4] ), .QN(n24980) );
  SDFFX1 \mem0_reg[77][3]  ( .D(n17175), .SI(\mem0[77][2] ), .SE(test_se), 
        .CLK(n1700), .Q(\mem0[77][3] ), .QN(n24981) );
  SDFFX1 \mem0_reg[77][2]  ( .D(n17174), .SI(\mem0[77][1] ), .SE(test_se), 
        .CLK(n1700), .Q(\mem0[77][2] ), .QN(n24982) );
  SDFFX1 \mem0_reg[77][1]  ( .D(n17173), .SI(\mem0[77][0] ), .SE(test_se), 
        .CLK(n1700), .Q(\mem0[77][1] ), .QN(n24983) );
  SDFFX1 \mem0_reg[77][0]  ( .D(n17172), .SI(\mem0[76][7] ), .SE(test_se), 
        .CLK(n1700), .Q(\mem0[77][0] ), .QN(n24984) );
  SDFFX1 \mem0_reg[76][7]  ( .D(n17171), .SI(\mem0[76][6] ), .SE(test_se), 
        .CLK(n1700), .Q(\mem0[76][7] ), .QN(n24985) );
  SDFFX1 \mem0_reg[76][6]  ( .D(n17170), .SI(\mem0[76][5] ), .SE(test_se), 
        .CLK(n1700), .Q(\mem0[76][6] ), .QN(n24986) );
  SDFFX1 \mem0_reg[76][5]  ( .D(n17169), .SI(\mem0[76][4] ), .SE(test_se), 
        .CLK(n1700), .Q(\mem0[76][5] ), .QN(n24987) );
  SDFFX1 \mem0_reg[76][4]  ( .D(n17168), .SI(\mem0[76][3] ), .SE(test_se), 
        .CLK(n1700), .Q(\mem0[76][4] ), .QN(n24988) );
  SDFFX1 \mem0_reg[76][3]  ( .D(n17167), .SI(\mem0[76][2] ), .SE(test_se), 
        .CLK(n1700), .Q(\mem0[76][3] ), .QN(n24989) );
  SDFFX1 \mem0_reg[76][2]  ( .D(n17166), .SI(\mem0[76][1] ), .SE(test_se), 
        .CLK(n1700), .Q(\mem0[76][2] ), .QN(n24990) );
  SDFFX1 \mem0_reg[76][1]  ( .D(n17165), .SI(\mem0[76][0] ), .SE(test_se), 
        .CLK(n1701), .Q(\mem0[76][1] ), .QN(n24991) );
  SDFFX1 \mem0_reg[76][0]  ( .D(n17164), .SI(\mem0[75][7] ), .SE(test_se), 
        .CLK(n1701), .Q(\mem0[76][0] ), .QN(n24992) );
  SDFFX1 \mem0_reg[75][7]  ( .D(n17163), .SI(\mem0[75][6] ), .SE(test_se), 
        .CLK(n1701), .Q(\mem0[75][7] ), .QN(n24993) );
  SDFFX1 \mem0_reg[75][6]  ( .D(n17162), .SI(\mem0[75][5] ), .SE(test_se), 
        .CLK(n1701), .Q(\mem0[75][6] ), .QN(n24994) );
  SDFFX1 \mem0_reg[75][5]  ( .D(n17161), .SI(\mem0[75][4] ), .SE(test_se), 
        .CLK(n1701), .Q(\mem0[75][5] ), .QN(n24995) );
  SDFFX1 \mem0_reg[75][4]  ( .D(n17160), .SI(\mem0[75][3] ), .SE(test_se), 
        .CLK(n1701), .Q(\mem0[75][4] ), .QN(n24996) );
  SDFFX1 \mem0_reg[75][3]  ( .D(n17159), .SI(\mem0[75][2] ), .SE(test_se), 
        .CLK(n1701), .Q(\mem0[75][3] ), .QN(n24997) );
  SDFFX1 \mem0_reg[75][2]  ( .D(n17158), .SI(\mem0[75][1] ), .SE(test_se), 
        .CLK(n1701), .Q(\mem0[75][2] ), .QN(n24998) );
  SDFFX1 \mem0_reg[75][1]  ( .D(n17157), .SI(\mem0[75][0] ), .SE(test_se), 
        .CLK(n1701), .Q(\mem0[75][1] ), .QN(n24999) );
  SDFFX1 \mem0_reg[75][0]  ( .D(n17156), .SI(\mem0[74][7] ), .SE(test_se), 
        .CLK(n1701), .Q(\mem0[75][0] ), .QN(n25000) );
  SDFFX1 \mem0_reg[74][7]  ( .D(n17155), .SI(\mem0[74][6] ), .SE(test_se), 
        .CLK(n1701), .Q(\mem0[74][7] ), .QN(n25001) );
  SDFFX1 \mem0_reg[74][6]  ( .D(n17154), .SI(\mem0[74][5] ), .SE(test_se), 
        .CLK(n1701), .Q(\mem0[74][6] ), .QN(n25002) );
  SDFFX1 \mem0_reg[74][5]  ( .D(n17153), .SI(\mem0[74][4] ), .SE(test_se), 
        .CLK(n1702), .Q(\mem0[74][5] ), .QN(n25003) );
  SDFFX1 \mem0_reg[74][4]  ( .D(n17152), .SI(\mem0[74][3] ), .SE(test_se), 
        .CLK(n1702), .Q(\mem0[74][4] ), .QN(n25004) );
  SDFFX1 \mem0_reg[74][3]  ( .D(n17151), .SI(\mem0[74][2] ), .SE(test_se), 
        .CLK(n1702), .Q(\mem0[74][3] ), .QN(n25005) );
  SDFFX1 \mem0_reg[74][2]  ( .D(n17150), .SI(\mem0[74][1] ), .SE(test_se), 
        .CLK(n1702), .Q(\mem0[74][2] ), .QN(n25006) );
  SDFFX1 \mem0_reg[74][1]  ( .D(n17149), .SI(\mem0[74][0] ), .SE(test_se), 
        .CLK(n1702), .Q(\mem0[74][1] ), .QN(n25007) );
  SDFFX1 \mem0_reg[74][0]  ( .D(n17148), .SI(\mem0[73][7] ), .SE(test_se), 
        .CLK(n1702), .Q(\mem0[74][0] ), .QN(n25008) );
  SDFFX1 \mem0_reg[73][7]  ( .D(n17147), .SI(\mem0[73][6] ), .SE(test_se), 
        .CLK(n1702), .Q(\mem0[73][7] ), .QN(n25009) );
  SDFFX1 \mem0_reg[73][6]  ( .D(n17146), .SI(\mem0[73][5] ), .SE(test_se), 
        .CLK(n1702), .Q(\mem0[73][6] ), .QN(n25010) );
  SDFFX1 \mem0_reg[73][5]  ( .D(n17145), .SI(\mem0[73][4] ), .SE(test_se), 
        .CLK(n1702), .Q(\mem0[73][5] ), .QN(n25011) );
  SDFFX1 \mem0_reg[73][4]  ( .D(n17144), .SI(\mem0[73][3] ), .SE(test_se), 
        .CLK(n1702), .Q(\mem0[73][4] ), .QN(n25012) );
  SDFFX1 \mem0_reg[73][3]  ( .D(n17143), .SI(\mem0[73][2] ), .SE(test_se), 
        .CLK(n1702), .Q(\mem0[73][3] ), .QN(n25013) );
  SDFFX1 \mem0_reg[73][2]  ( .D(n17142), .SI(\mem0[73][1] ), .SE(test_se), 
        .CLK(n1702), .Q(\mem0[73][2] ), .QN(n25014) );
  SDFFX1 \mem0_reg[73][1]  ( .D(n17141), .SI(\mem0[73][0] ), .SE(test_se), 
        .CLK(n1703), .Q(\mem0[73][1] ), .QN(n25015) );
  SDFFX1 \mem0_reg[73][0]  ( .D(n17140), .SI(\mem0[72][7] ), .SE(test_se), 
        .CLK(n1703), .Q(\mem0[73][0] ), .QN(n25016) );
  SDFFX1 \mem0_reg[72][7]  ( .D(n17139), .SI(\mem0[72][6] ), .SE(test_se), 
        .CLK(n1703), .Q(\mem0[72][7] ), .QN(n25017) );
  SDFFX1 \mem0_reg[72][6]  ( .D(n17138), .SI(\mem0[72][5] ), .SE(test_se), 
        .CLK(n1703), .Q(\mem0[72][6] ), .QN(n25018) );
  SDFFX1 \mem0_reg[72][5]  ( .D(n17137), .SI(\mem0[72][4] ), .SE(test_se), 
        .CLK(n1703), .Q(\mem0[72][5] ), .QN(n25019) );
  SDFFX1 \mem0_reg[72][4]  ( .D(n17136), .SI(\mem0[72][3] ), .SE(test_se), 
        .CLK(n1703), .Q(\mem0[72][4] ), .QN(n25020) );
  SDFFX1 \mem0_reg[72][3]  ( .D(n17135), .SI(\mem0[72][2] ), .SE(test_se), 
        .CLK(n1703), .Q(\mem0[72][3] ), .QN(n25021) );
  SDFFX1 \mem0_reg[72][2]  ( .D(n17134), .SI(\mem0[72][1] ), .SE(test_se), 
        .CLK(n1703), .Q(\mem0[72][2] ), .QN(n25022) );
  SDFFX1 \mem0_reg[72][1]  ( .D(n17133), .SI(\mem0[72][0] ), .SE(test_se), 
        .CLK(n1703), .Q(\mem0[72][1] ), .QN(n25023) );
  SDFFX1 \mem0_reg[72][0]  ( .D(n17132), .SI(\mem0[71][7] ), .SE(test_se), 
        .CLK(n1703), .Q(\mem0[72][0] ), .QN(n25024) );
  SDFFX1 \mem0_reg[71][7]  ( .D(n17131), .SI(\mem0[71][6] ), .SE(test_se), 
        .CLK(n1703), .Q(\mem0[71][7] ), .QN(n25025) );
  SDFFX1 \mem0_reg[71][6]  ( .D(n17130), .SI(\mem0[71][5] ), .SE(test_se), 
        .CLK(n1703), .Q(\mem0[71][6] ), .QN(n25026) );
  SDFFX1 \mem0_reg[71][5]  ( .D(n17129), .SI(\mem0[71][4] ), .SE(test_se), 
        .CLK(n1704), .Q(\mem0[71][5] ), .QN(n25027) );
  SDFFX1 \mem0_reg[71][4]  ( .D(n17128), .SI(\mem0[71][3] ), .SE(test_se), 
        .CLK(n1704), .Q(\mem0[71][4] ), .QN(n25028) );
  SDFFX1 \mem0_reg[71][3]  ( .D(n17127), .SI(\mem0[71][2] ), .SE(test_se), 
        .CLK(n1704), .Q(\mem0[71][3] ), .QN(n25029) );
  SDFFX1 \mem0_reg[71][2]  ( .D(n17126), .SI(\mem0[71][1] ), .SE(test_se), 
        .CLK(n1704), .Q(\mem0[71][2] ), .QN(n25030) );
  SDFFX1 \mem0_reg[71][1]  ( .D(n17125), .SI(\mem0[71][0] ), .SE(test_se), 
        .CLK(n1704), .Q(\mem0[71][1] ), .QN(n25031) );
  SDFFX1 \mem0_reg[71][0]  ( .D(n17124), .SI(\mem0[70][7] ), .SE(test_se), 
        .CLK(n1704), .Q(\mem0[71][0] ), .QN(n25032) );
  SDFFX1 \mem0_reg[70][7]  ( .D(n17123), .SI(\mem0[70][6] ), .SE(test_se), 
        .CLK(n1704), .Q(\mem0[70][7] ), .QN(n25033) );
  SDFFX1 \mem0_reg[70][6]  ( .D(n17122), .SI(\mem0[70][5] ), .SE(test_se), 
        .CLK(n1704), .Q(\mem0[70][6] ), .QN(n25034) );
  SDFFX1 \mem0_reg[70][5]  ( .D(n17121), .SI(\mem0[70][4] ), .SE(test_se), 
        .CLK(n1704), .Q(\mem0[70][5] ), .QN(n25035) );
  SDFFX1 \mem0_reg[70][4]  ( .D(n17120), .SI(\mem0[70][3] ), .SE(test_se), 
        .CLK(n1704), .Q(\mem0[70][4] ), .QN(n25036) );
  SDFFX1 \mem0_reg[70][3]  ( .D(n17119), .SI(\mem0[70][2] ), .SE(test_se), 
        .CLK(n1704), .Q(\mem0[70][3] ), .QN(n25037) );
  SDFFX1 \mem0_reg[70][2]  ( .D(n17118), .SI(\mem0[70][1] ), .SE(test_se), 
        .CLK(n1704), .Q(\mem0[70][2] ), .QN(n25038) );
  SDFFX1 \mem0_reg[70][1]  ( .D(n17117), .SI(\mem0[70][0] ), .SE(test_se), 
        .CLK(n1705), .Q(\mem0[70][1] ), .QN(n25039) );
  SDFFX1 \mem0_reg[70][0]  ( .D(n17116), .SI(\mem0[69][7] ), .SE(test_se), 
        .CLK(n1705), .Q(\mem0[70][0] ), .QN(n25040) );
  SDFFX1 \mem0_reg[69][7]  ( .D(n17115), .SI(\mem0[69][6] ), .SE(test_se), 
        .CLK(n1705), .Q(\mem0[69][7] ), .QN(n25041) );
  SDFFX1 \mem0_reg[69][6]  ( .D(n17114), .SI(\mem0[69][5] ), .SE(test_se), 
        .CLK(n1705), .Q(\mem0[69][6] ), .QN(n25042) );
  SDFFX1 \mem0_reg[69][5]  ( .D(n17113), .SI(\mem0[69][4] ), .SE(test_se), 
        .CLK(n1705), .Q(\mem0[69][5] ), .QN(n25043) );
  SDFFX1 \mem0_reg[69][4]  ( .D(n17112), .SI(\mem0[69][3] ), .SE(test_se), 
        .CLK(n1705), .Q(\mem0[69][4] ), .QN(n25044) );
  SDFFX1 \mem0_reg[69][3]  ( .D(n17111), .SI(\mem0[69][2] ), .SE(test_se), 
        .CLK(n1705), .Q(\mem0[69][3] ), .QN(n25045) );
  SDFFX1 \mem0_reg[69][2]  ( .D(n17110), .SI(\mem0[69][1] ), .SE(test_se), 
        .CLK(n1705), .Q(\mem0[69][2] ), .QN(n25046) );
  SDFFX1 \mem0_reg[69][1]  ( .D(n17109), .SI(\mem0[69][0] ), .SE(test_se), 
        .CLK(n1705), .Q(\mem0[69][1] ), .QN(n25047) );
  SDFFX1 \mem0_reg[69][0]  ( .D(n17108), .SI(\mem0[68][7] ), .SE(test_se), 
        .CLK(n1705), .Q(\mem0[69][0] ), .QN(n25048) );
  SDFFX1 \mem0_reg[68][7]  ( .D(n17107), .SI(\mem0[68][6] ), .SE(test_se), 
        .CLK(n1705), .Q(\mem0[68][7] ), .QN(n25049) );
  SDFFX1 \mem0_reg[68][6]  ( .D(n17106), .SI(\mem0[68][5] ), .SE(test_se), 
        .CLK(n1705), .Q(\mem0[68][6] ), .QN(n25050) );
  SDFFX1 \mem0_reg[68][5]  ( .D(n17105), .SI(\mem0[68][4] ), .SE(test_se), 
        .CLK(n1706), .Q(\mem0[68][5] ), .QN(n25051) );
  SDFFX1 \mem0_reg[68][4]  ( .D(n17104), .SI(\mem0[68][3] ), .SE(test_se), 
        .CLK(n1706), .Q(\mem0[68][4] ), .QN(n25052) );
  SDFFX1 \mem0_reg[68][3]  ( .D(n17103), .SI(\mem0[68][2] ), .SE(test_se), 
        .CLK(n1706), .Q(\mem0[68][3] ), .QN(n25053) );
  SDFFX1 \mem0_reg[68][2]  ( .D(n17102), .SI(\mem0[68][1] ), .SE(test_se), 
        .CLK(n1706), .Q(\mem0[68][2] ), .QN(n25054) );
  SDFFX1 \mem0_reg[68][1]  ( .D(n17101), .SI(\mem0[68][0] ), .SE(test_se), 
        .CLK(n1706), .Q(\mem0[68][1] ), .QN(n25055) );
  SDFFX1 \mem0_reg[68][0]  ( .D(n17100), .SI(\mem0[67][7] ), .SE(test_se), 
        .CLK(n1706), .Q(\mem0[68][0] ), .QN(n25056) );
  SDFFX1 \mem0_reg[67][7]  ( .D(n17099), .SI(\mem0[67][6] ), .SE(test_se), 
        .CLK(n1706), .Q(\mem0[67][7] ), .QN(n25057) );
  SDFFX1 \mem0_reg[67][6]  ( .D(n17098), .SI(\mem0[67][5] ), .SE(test_se), 
        .CLK(n1706), .Q(\mem0[67][6] ), .QN(n25058) );
  SDFFX1 \mem0_reg[67][5]  ( .D(n17097), .SI(\mem0[67][4] ), .SE(test_se), 
        .CLK(n1706), .Q(\mem0[67][5] ), .QN(n25059) );
  SDFFX1 \mem0_reg[67][4]  ( .D(n17096), .SI(\mem0[67][3] ), .SE(test_se), 
        .CLK(n1706), .Q(\mem0[67][4] ), .QN(n25060) );
  SDFFX1 \mem0_reg[67][3]  ( .D(n17095), .SI(\mem0[67][2] ), .SE(test_se), 
        .CLK(n1706), .Q(\mem0[67][3] ), .QN(n25061) );
  SDFFX1 \mem0_reg[67][2]  ( .D(n17094), .SI(\mem0[67][1] ), .SE(test_se), 
        .CLK(n1706), .Q(\mem0[67][2] ), .QN(n25062) );
  SDFFX1 \mem0_reg[67][1]  ( .D(n17093), .SI(\mem0[67][0] ), .SE(test_se), 
        .CLK(n1707), .Q(\mem0[67][1] ), .QN(n25063) );
  SDFFX1 \mem0_reg[67][0]  ( .D(n17092), .SI(\mem0[66][7] ), .SE(test_se), 
        .CLK(n1707), .Q(\mem0[67][0] ), .QN(n25064) );
  SDFFX1 \mem0_reg[66][7]  ( .D(n17091), .SI(\mem0[66][6] ), .SE(test_se), 
        .CLK(n1707), .Q(\mem0[66][7] ), .QN(n25065) );
  SDFFX1 \mem0_reg[66][6]  ( .D(n17090), .SI(\mem0[66][5] ), .SE(test_se), 
        .CLK(n1707), .Q(\mem0[66][6] ), .QN(n25066) );
  SDFFX1 \mem0_reg[66][5]  ( .D(n17089), .SI(\mem0[66][4] ), .SE(test_se), 
        .CLK(n1707), .Q(\mem0[66][5] ), .QN(n25067) );
  SDFFX1 \mem0_reg[66][4]  ( .D(n17088), .SI(\mem0[66][3] ), .SE(test_se), 
        .CLK(n1707), .Q(\mem0[66][4] ), .QN(n25068) );
  SDFFX1 \mem0_reg[66][3]  ( .D(n17087), .SI(\mem0[66][2] ), .SE(test_se), 
        .CLK(n1707), .Q(\mem0[66][3] ), .QN(n25069) );
  SDFFX1 \mem0_reg[66][2]  ( .D(n17086), .SI(\mem0[66][1] ), .SE(test_se), 
        .CLK(n1707), .Q(\mem0[66][2] ), .QN(n25070) );
  SDFFX1 \mem0_reg[66][1]  ( .D(n17085), .SI(\mem0[66][0] ), .SE(test_se), 
        .CLK(n1707), .Q(\mem0[66][1] ), .QN(n25071) );
  SDFFX1 \mem0_reg[66][0]  ( .D(n17084), .SI(\mem0[65][7] ), .SE(test_se), 
        .CLK(n1707), .Q(\mem0[66][0] ), .QN(n25072) );
  SDFFX1 \mem0_reg[65][7]  ( .D(n17083), .SI(\mem0[65][6] ), .SE(test_se), 
        .CLK(n1707), .Q(\mem0[65][7] ), .QN(n25073) );
  SDFFX1 \mem0_reg[65][6]  ( .D(n17082), .SI(\mem0[65][5] ), .SE(test_se), 
        .CLK(n1707), .Q(\mem0[65][6] ), .QN(n25074) );
  SDFFX1 \mem0_reg[65][5]  ( .D(n17081), .SI(\mem0[65][4] ), .SE(test_se), 
        .CLK(n1708), .Q(\mem0[65][5] ), .QN(n25075) );
  SDFFX1 \mem0_reg[65][4]  ( .D(n17080), .SI(\mem0[65][3] ), .SE(test_se), 
        .CLK(n1708), .Q(\mem0[65][4] ), .QN(n25076) );
  SDFFX1 \mem0_reg[65][3]  ( .D(n17079), .SI(\mem0[65][2] ), .SE(test_se), 
        .CLK(n1708), .Q(\mem0[65][3] ), .QN(n25077) );
  SDFFX1 \mem0_reg[65][2]  ( .D(n17078), .SI(\mem0[65][1] ), .SE(test_se), 
        .CLK(n1708), .Q(\mem0[65][2] ), .QN(n25078) );
  SDFFX1 \mem0_reg[65][1]  ( .D(n17077), .SI(\mem0[65][0] ), .SE(test_se), 
        .CLK(n1708), .Q(\mem0[65][1] ), .QN(n25079) );
  SDFFX1 \mem0_reg[65][0]  ( .D(n17076), .SI(\mem0[64][7] ), .SE(test_se), 
        .CLK(n1708), .Q(\mem0[65][0] ), .QN(n25080) );
  SDFFX1 \mem0_reg[64][7]  ( .D(n17075), .SI(\mem0[64][6] ), .SE(test_se), 
        .CLK(n1708), .Q(\mem0[64][7] ), .QN(n25081) );
  SDFFX1 \mem0_reg[64][6]  ( .D(n17074), .SI(\mem0[64][5] ), .SE(test_se), 
        .CLK(n1708), .Q(\mem0[64][6] ), .QN(n25082) );
  SDFFX1 \mem0_reg[64][5]  ( .D(n17073), .SI(\mem0[64][4] ), .SE(test_se), 
        .CLK(n1708), .Q(\mem0[64][5] ), .QN(n25083) );
  SDFFX1 \mem0_reg[64][4]  ( .D(n17072), .SI(\mem0[64][3] ), .SE(test_se), 
        .CLK(n1708), .Q(\mem0[64][4] ), .QN(n25084) );
  SDFFX1 \mem0_reg[64][3]  ( .D(n17071), .SI(\mem0[64][2] ), .SE(test_se), 
        .CLK(n1708), .Q(\mem0[64][3] ), .QN(n25085) );
  SDFFX1 \mem0_reg[64][2]  ( .D(n17070), .SI(\mem0[64][1] ), .SE(test_se), 
        .CLK(n1708), .Q(\mem0[64][2] ), .QN(n25086) );
  SDFFX1 \mem0_reg[64][1]  ( .D(n17069), .SI(\mem0[64][0] ), .SE(test_se), 
        .CLK(n1709), .Q(\mem0[64][1] ), .QN(n25087) );
  SDFFX1 \mem0_reg[64][0]  ( .D(n17068), .SI(\mem0[63][7] ), .SE(test_se), 
        .CLK(n1709), .Q(\mem0[64][0] ), .QN(n25088) );
  SDFFX1 \mem0_reg[63][7]  ( .D(n17067), .SI(\mem0[63][6] ), .SE(test_se), 
        .CLK(n1709), .Q(\mem0[63][7] ), .QN(n25089) );
  SDFFX1 \mem0_reg[63][6]  ( .D(n17066), .SI(\mem0[63][5] ), .SE(test_se), 
        .CLK(n1709), .Q(\mem0[63][6] ), .QN(n25090) );
  SDFFX1 \mem0_reg[63][5]  ( .D(n17065), .SI(\mem0[63][4] ), .SE(test_se), 
        .CLK(n1709), .Q(\mem0[63][5] ), .QN(n25091) );
  SDFFX1 \mem0_reg[63][4]  ( .D(n17064), .SI(\mem0[63][3] ), .SE(test_se), 
        .CLK(n1709), .Q(\mem0[63][4] ), .QN(n25092) );
  SDFFX1 \mem0_reg[63][3]  ( .D(n17063), .SI(\mem0[63][2] ), .SE(test_se), 
        .CLK(n1709), .Q(\mem0[63][3] ), .QN(n25093) );
  SDFFX1 \mem0_reg[63][2]  ( .D(n17062), .SI(\mem0[63][1] ), .SE(test_se), 
        .CLK(n1709), .Q(\mem0[63][2] ), .QN(n25094) );
  SDFFX1 \mem0_reg[63][1]  ( .D(n17061), .SI(\mem0[63][0] ), .SE(test_se), 
        .CLK(n1709), .Q(\mem0[63][1] ), .QN(n25095) );
  SDFFX1 \mem0_reg[63][0]  ( .D(n17060), .SI(\mem0[62][7] ), .SE(test_se), 
        .CLK(n1709), .Q(\mem0[63][0] ), .QN(n25096) );
  SDFFX1 \mem0_reg[62][7]  ( .D(n17059), .SI(\mem0[62][6] ), .SE(test_se), 
        .CLK(n1709), .Q(\mem0[62][7] ), .QN(n25097) );
  SDFFX1 \mem0_reg[62][6]  ( .D(n17058), .SI(\mem0[62][5] ), .SE(test_se), 
        .CLK(n1709), .Q(\mem0[62][6] ), .QN(n25098) );
  SDFFX1 \mem0_reg[62][5]  ( .D(n17057), .SI(\mem0[62][4] ), .SE(test_se), 
        .CLK(n1710), .Q(\mem0[62][5] ), .QN(n25099) );
  SDFFX1 \mem0_reg[62][4]  ( .D(n17056), .SI(\mem0[62][3] ), .SE(test_se), 
        .CLK(n1710), .Q(\mem0[62][4] ), .QN(n25100) );
  SDFFX1 \mem0_reg[62][3]  ( .D(n17055), .SI(\mem0[62][2] ), .SE(test_se), 
        .CLK(n1710), .Q(\mem0[62][3] ), .QN(n25101) );
  SDFFX1 \mem0_reg[62][2]  ( .D(n17054), .SI(\mem0[62][1] ), .SE(test_se), 
        .CLK(n1710), .Q(\mem0[62][2] ), .QN(n25102) );
  SDFFX1 \mem0_reg[62][1]  ( .D(n17053), .SI(\mem0[62][0] ), .SE(test_se), 
        .CLK(n1710), .Q(\mem0[62][1] ), .QN(n25103) );
  SDFFX1 \mem0_reg[62][0]  ( .D(n17052), .SI(\mem0[61][7] ), .SE(test_se), 
        .CLK(n1710), .Q(\mem0[62][0] ), .QN(n25104) );
  SDFFX1 \mem0_reg[61][7]  ( .D(n17051), .SI(\mem0[61][6] ), .SE(test_se), 
        .CLK(n1710), .Q(\mem0[61][7] ), .QN(n25105) );
  SDFFX1 \mem0_reg[61][6]  ( .D(n17050), .SI(\mem0[61][5] ), .SE(test_se), 
        .CLK(n1710), .Q(\mem0[61][6] ), .QN(n25106) );
  SDFFX1 \mem0_reg[61][5]  ( .D(n17049), .SI(\mem0[61][4] ), .SE(test_se), 
        .CLK(n1710), .Q(\mem0[61][5] ), .QN(n25107) );
  SDFFX1 \mem0_reg[61][4]  ( .D(n17048), .SI(\mem0[61][3] ), .SE(test_se), 
        .CLK(n1710), .Q(\mem0[61][4] ), .QN(n25108) );
  SDFFX1 \mem0_reg[61][3]  ( .D(n17047), .SI(\mem0[61][2] ), .SE(test_se), 
        .CLK(n1710), .Q(\mem0[61][3] ), .QN(n25109) );
  SDFFX1 \mem0_reg[61][2]  ( .D(n17046), .SI(\mem0[61][1] ), .SE(test_se), 
        .CLK(n1710), .Q(\mem0[61][2] ), .QN(n25110) );
  SDFFX1 \mem0_reg[61][1]  ( .D(n17045), .SI(\mem0[61][0] ), .SE(test_se), 
        .CLK(n1711), .Q(\mem0[61][1] ), .QN(n25111) );
  SDFFX1 \mem0_reg[61][0]  ( .D(n17044), .SI(\mem0[60][7] ), .SE(test_se), 
        .CLK(n1711), .Q(\mem0[61][0] ), .QN(n25112) );
  SDFFX1 \mem0_reg[60][7]  ( .D(n17043), .SI(\mem0[60][6] ), .SE(test_se), 
        .CLK(n1711), .Q(\mem0[60][7] ), .QN(n25113) );
  SDFFX1 \mem0_reg[60][6]  ( .D(n17042), .SI(\mem0[60][5] ), .SE(test_se), 
        .CLK(n1711), .Q(\mem0[60][6] ), .QN(n25114) );
  SDFFX1 \mem0_reg[60][5]  ( .D(n17041), .SI(\mem0[60][4] ), .SE(test_se), 
        .CLK(n1711), .Q(\mem0[60][5] ), .QN(n25115) );
  SDFFX1 \mem0_reg[60][4]  ( .D(n17040), .SI(\mem0[60][3] ), .SE(test_se), 
        .CLK(n1711), .Q(\mem0[60][4] ), .QN(n25116) );
  SDFFX1 \mem0_reg[60][3]  ( .D(n17039), .SI(\mem0[60][2] ), .SE(test_se), 
        .CLK(n1711), .Q(\mem0[60][3] ), .QN(n25117) );
  SDFFX1 \mem0_reg[60][2]  ( .D(n17038), .SI(\mem0[60][1] ), .SE(test_se), 
        .CLK(n1711), .Q(\mem0[60][2] ), .QN(n25118) );
  SDFFX1 \mem0_reg[60][1]  ( .D(n17037), .SI(\mem0[60][0] ), .SE(test_se), 
        .CLK(n1711), .Q(\mem0[60][1] ), .QN(n25119) );
  SDFFX1 \mem0_reg[60][0]  ( .D(n17036), .SI(\mem0[59][7] ), .SE(test_se), 
        .CLK(n1711), .Q(\mem0[60][0] ), .QN(n25120) );
  SDFFX1 \mem0_reg[59][7]  ( .D(n17035), .SI(\mem0[59][6] ), .SE(test_se), 
        .CLK(n1711), .Q(\mem0[59][7] ), .QN(n25121) );
  SDFFX1 \mem0_reg[59][6]  ( .D(n17034), .SI(\mem0[59][5] ), .SE(test_se), 
        .CLK(n1711), .Q(\mem0[59][6] ), .QN(n25122) );
  SDFFX1 \mem0_reg[59][5]  ( .D(n17033), .SI(\mem0[59][4] ), .SE(test_se), 
        .CLK(n1712), .Q(\mem0[59][5] ), .QN(n25123) );
  SDFFX1 \mem0_reg[59][4]  ( .D(n17032), .SI(\mem0[59][3] ), .SE(test_se), 
        .CLK(n1712), .Q(\mem0[59][4] ), .QN(n25124) );
  SDFFX1 \mem0_reg[59][3]  ( .D(n17031), .SI(\mem0[59][2] ), .SE(test_se), 
        .CLK(n1712), .Q(\mem0[59][3] ), .QN(n25125) );
  SDFFX1 \mem0_reg[59][2]  ( .D(n17030), .SI(\mem0[59][1] ), .SE(test_se), 
        .CLK(n1712), .Q(\mem0[59][2] ), .QN(n25126) );
  SDFFX1 \mem0_reg[59][1]  ( .D(n17029), .SI(\mem0[59][0] ), .SE(test_se), 
        .CLK(n1712), .Q(\mem0[59][1] ), .QN(n25127) );
  SDFFX1 \mem0_reg[59][0]  ( .D(n17028), .SI(\mem0[58][7] ), .SE(test_se), 
        .CLK(n1712), .Q(\mem0[59][0] ), .QN(n25128) );
  SDFFX1 \mem0_reg[58][7]  ( .D(n17027), .SI(\mem0[58][6] ), .SE(test_se), 
        .CLK(n1712), .Q(\mem0[58][7] ), .QN(n25129) );
  SDFFX1 \mem0_reg[58][6]  ( .D(n17026), .SI(\mem0[58][5] ), .SE(test_se), 
        .CLK(n1712), .Q(\mem0[58][6] ), .QN(n25130) );
  SDFFX1 \mem0_reg[58][5]  ( .D(n17025), .SI(\mem0[58][4] ), .SE(test_se), 
        .CLK(n1712), .Q(\mem0[58][5] ), .QN(n25131) );
  SDFFX1 \mem0_reg[58][4]  ( .D(n17024), .SI(\mem0[58][3] ), .SE(test_se), 
        .CLK(n1712), .Q(\mem0[58][4] ), .QN(n25132) );
  SDFFX1 \mem0_reg[58][3]  ( .D(n17023), .SI(\mem0[58][2] ), .SE(test_se), 
        .CLK(n1712), .Q(\mem0[58][3] ), .QN(n25133) );
  SDFFX1 \mem0_reg[58][2]  ( .D(n17022), .SI(\mem0[58][1] ), .SE(test_se), 
        .CLK(n1712), .Q(\mem0[58][2] ), .QN(n25134) );
  SDFFX1 \mem0_reg[58][1]  ( .D(n17021), .SI(\mem0[58][0] ), .SE(test_se), 
        .CLK(n1713), .Q(\mem0[58][1] ), .QN(n25135) );
  SDFFX1 \mem0_reg[58][0]  ( .D(n17020), .SI(\mem0[57][7] ), .SE(test_se), 
        .CLK(n1713), .Q(\mem0[58][0] ), .QN(n25136) );
  SDFFX1 \mem0_reg[57][7]  ( .D(n17019), .SI(\mem0[57][6] ), .SE(test_se), 
        .CLK(n1713), .Q(\mem0[57][7] ), .QN(n25137) );
  SDFFX1 \mem0_reg[57][6]  ( .D(n17018), .SI(\mem0[57][5] ), .SE(test_se), 
        .CLK(n1713), .Q(\mem0[57][6] ), .QN(n25138) );
  SDFFX1 \mem0_reg[57][5]  ( .D(n17017), .SI(\mem0[57][4] ), .SE(test_se), 
        .CLK(n1713), .Q(\mem0[57][5] ), .QN(n25139) );
  SDFFX1 \mem0_reg[57][4]  ( .D(n17016), .SI(\mem0[57][3] ), .SE(test_se), 
        .CLK(n1713), .Q(\mem0[57][4] ), .QN(n25140) );
  SDFFX1 \mem0_reg[57][3]  ( .D(n17015), .SI(\mem0[57][2] ), .SE(test_se), 
        .CLK(n1713), .Q(\mem0[57][3] ), .QN(n25141) );
  SDFFX1 \mem0_reg[57][2]  ( .D(n17014), .SI(\mem0[57][1] ), .SE(test_se), 
        .CLK(n1713), .Q(\mem0[57][2] ), .QN(n25142) );
  SDFFX1 \mem0_reg[57][1]  ( .D(n17013), .SI(\mem0[57][0] ), .SE(test_se), 
        .CLK(n1713), .Q(\mem0[57][1] ), .QN(n25143) );
  SDFFX1 \mem0_reg[57][0]  ( .D(n17012), .SI(\mem0[56][7] ), .SE(test_se), 
        .CLK(n1713), .Q(\mem0[57][0] ), .QN(n25144) );
  SDFFX1 \mem0_reg[56][7]  ( .D(n17011), .SI(\mem0[56][6] ), .SE(test_se), 
        .CLK(n1713), .Q(\mem0[56][7] ), .QN(n25145) );
  SDFFX1 \mem0_reg[56][6]  ( .D(n17010), .SI(\mem0[56][5] ), .SE(test_se), 
        .CLK(n1713), .Q(\mem0[56][6] ), .QN(n25146) );
  SDFFX1 \mem0_reg[56][5]  ( .D(n17009), .SI(\mem0[56][4] ), .SE(test_se), 
        .CLK(n1714), .Q(\mem0[56][5] ), .QN(n25147) );
  SDFFX1 \mem0_reg[56][4]  ( .D(n17008), .SI(\mem0[56][3] ), .SE(test_se), 
        .CLK(n1714), .Q(\mem0[56][4] ), .QN(n25148) );
  SDFFX1 \mem0_reg[56][3]  ( .D(n17007), .SI(\mem0[56][2] ), .SE(test_se), 
        .CLK(n1714), .Q(\mem0[56][3] ), .QN(n25149) );
  SDFFX1 \mem0_reg[56][2]  ( .D(n17006), .SI(\mem0[56][1] ), .SE(test_se), 
        .CLK(n1714), .Q(\mem0[56][2] ), .QN(n25150) );
  SDFFX1 \mem0_reg[56][1]  ( .D(n17005), .SI(\mem0[56][0] ), .SE(test_se), 
        .CLK(n1714), .Q(\mem0[56][1] ), .QN(n25151) );
  SDFFX1 \mem0_reg[56][0]  ( .D(n17004), .SI(\mem0[55][7] ), .SE(test_se), 
        .CLK(n1714), .Q(\mem0[56][0] ), .QN(n25152) );
  SDFFX1 \mem0_reg[55][7]  ( .D(n17003), .SI(\mem0[55][6] ), .SE(test_se), 
        .CLK(n1714), .Q(\mem0[55][7] ), .QN(n25153) );
  SDFFX1 \mem0_reg[55][6]  ( .D(n17002), .SI(\mem0[55][5] ), .SE(test_se), 
        .CLK(n1714), .Q(\mem0[55][6] ), .QN(n25154) );
  SDFFX1 \mem0_reg[55][5]  ( .D(n17001), .SI(\mem0[55][4] ), .SE(test_se), 
        .CLK(n1714), .Q(\mem0[55][5] ), .QN(n25155) );
  SDFFX1 \mem0_reg[55][4]  ( .D(n17000), .SI(\mem0[55][3] ), .SE(test_se), 
        .CLK(n1714), .Q(\mem0[55][4] ), .QN(n25156) );
  SDFFX1 \mem0_reg[55][3]  ( .D(n16999), .SI(\mem0[55][2] ), .SE(test_se), 
        .CLK(n1714), .Q(\mem0[55][3] ), .QN(n25157) );
  SDFFX1 \mem0_reg[55][2]  ( .D(n16998), .SI(\mem0[55][1] ), .SE(test_se), 
        .CLK(n1714), .Q(\mem0[55][2] ), .QN(n25158) );
  SDFFX1 \mem0_reg[55][1]  ( .D(n16997), .SI(\mem0[55][0] ), .SE(test_se), 
        .CLK(n1715), .Q(\mem0[55][1] ), .QN(n25159) );
  SDFFX1 \mem0_reg[55][0]  ( .D(n16996), .SI(\mem0[54][7] ), .SE(test_se), 
        .CLK(n1715), .Q(\mem0[55][0] ), .QN(n25160) );
  SDFFX1 \mem0_reg[54][7]  ( .D(n16995), .SI(\mem0[54][6] ), .SE(test_se), 
        .CLK(n1715), .Q(\mem0[54][7] ), .QN(n25161) );
  SDFFX1 \mem0_reg[54][6]  ( .D(n16994), .SI(\mem0[54][5] ), .SE(test_se), 
        .CLK(n1715), .Q(\mem0[54][6] ), .QN(n25162) );
  SDFFX1 \mem0_reg[54][5]  ( .D(n16993), .SI(\mem0[54][4] ), .SE(test_se), 
        .CLK(n1715), .Q(\mem0[54][5] ), .QN(n25163) );
  SDFFX1 \mem0_reg[54][4]  ( .D(n16992), .SI(\mem0[54][3] ), .SE(test_se), 
        .CLK(n1715), .Q(\mem0[54][4] ), .QN(n25164) );
  SDFFX1 \mem0_reg[54][3]  ( .D(n16991), .SI(\mem0[54][2] ), .SE(test_se), 
        .CLK(n1715), .Q(\mem0[54][3] ), .QN(n25165) );
  SDFFX1 \mem0_reg[54][2]  ( .D(n16990), .SI(\mem0[54][1] ), .SE(test_se), 
        .CLK(n1715), .Q(\mem0[54][2] ), .QN(n25166) );
  SDFFX1 \mem0_reg[54][1]  ( .D(n16989), .SI(\mem0[54][0] ), .SE(test_se), 
        .CLK(n1715), .Q(\mem0[54][1] ), .QN(n25167) );
  SDFFX1 \mem0_reg[54][0]  ( .D(n16988), .SI(\mem0[53][7] ), .SE(test_se), 
        .CLK(n1715), .Q(\mem0[54][0] ), .QN(n25168) );
  SDFFX1 \mem0_reg[53][7]  ( .D(n16987), .SI(\mem0[53][6] ), .SE(test_se), 
        .CLK(n1715), .Q(\mem0[53][7] ), .QN(n25169) );
  SDFFX1 \mem0_reg[53][6]  ( .D(n16986), .SI(\mem0[53][5] ), .SE(test_se), 
        .CLK(n1715), .Q(\mem0[53][6] ), .QN(n25170) );
  SDFFX1 \mem0_reg[53][5]  ( .D(n16985), .SI(\mem0[53][4] ), .SE(test_se), 
        .CLK(n1716), .Q(\mem0[53][5] ), .QN(n25171) );
  SDFFX1 \mem0_reg[53][4]  ( .D(n16984), .SI(\mem0[53][3] ), .SE(test_se), 
        .CLK(n1716), .Q(\mem0[53][4] ), .QN(n25172) );
  SDFFX1 \mem0_reg[53][3]  ( .D(n16983), .SI(\mem0[53][2] ), .SE(test_se), 
        .CLK(n1716), .Q(\mem0[53][3] ), .QN(n25173) );
  SDFFX1 \mem0_reg[53][2]  ( .D(n16982), .SI(\mem0[53][1] ), .SE(test_se), 
        .CLK(n1716), .Q(\mem0[53][2] ), .QN(n25174) );
  SDFFX1 \mem0_reg[53][1]  ( .D(n16981), .SI(\mem0[53][0] ), .SE(test_se), 
        .CLK(n1716), .Q(\mem0[53][1] ), .QN(n25175) );
  SDFFX1 \mem0_reg[53][0]  ( .D(n16980), .SI(\mem0[52][7] ), .SE(test_se), 
        .CLK(n1716), .Q(\mem0[53][0] ), .QN(n25176) );
  SDFFX1 \mem0_reg[52][7]  ( .D(n16979), .SI(\mem0[52][6] ), .SE(test_se), 
        .CLK(n1716), .Q(\mem0[52][7] ), .QN(n25177) );
  SDFFX1 \mem0_reg[52][6]  ( .D(n16978), .SI(\mem0[52][5] ), .SE(test_se), 
        .CLK(n1716), .Q(\mem0[52][6] ), .QN(n25178) );
  SDFFX1 \mem0_reg[52][5]  ( .D(n16977), .SI(\mem0[52][4] ), .SE(test_se), 
        .CLK(n1716), .Q(\mem0[52][5] ), .QN(n25179) );
  SDFFX1 \mem0_reg[52][4]  ( .D(n16976), .SI(\mem0[52][3] ), .SE(test_se), 
        .CLK(n1716), .Q(\mem0[52][4] ), .QN(n25180) );
  SDFFX1 \mem0_reg[52][3]  ( .D(n16975), .SI(\mem0[52][2] ), .SE(test_se), 
        .CLK(n1716), .Q(\mem0[52][3] ), .QN(n25181) );
  SDFFX1 \mem0_reg[52][2]  ( .D(n16974), .SI(\mem0[52][1] ), .SE(test_se), 
        .CLK(n1716), .Q(\mem0[52][2] ), .QN(n25182) );
  SDFFX1 \mem0_reg[52][1]  ( .D(n16973), .SI(\mem0[52][0] ), .SE(test_se), 
        .CLK(n1717), .Q(\mem0[52][1] ), .QN(n25183) );
  SDFFX1 \mem0_reg[52][0]  ( .D(n16972), .SI(\mem0[51][7] ), .SE(test_se), 
        .CLK(n1717), .Q(\mem0[52][0] ), .QN(n25184) );
  SDFFX1 \mem0_reg[51][7]  ( .D(n16971), .SI(\mem0[51][6] ), .SE(test_se), 
        .CLK(n1717), .Q(\mem0[51][7] ), .QN(n25185) );
  SDFFX1 \mem0_reg[51][6]  ( .D(n16970), .SI(\mem0[51][5] ), .SE(test_se), 
        .CLK(n1717), .Q(\mem0[51][6] ), .QN(n25186) );
  SDFFX1 \mem0_reg[51][5]  ( .D(n16969), .SI(\mem0[51][4] ), .SE(test_se), 
        .CLK(n1717), .Q(\mem0[51][5] ), .QN(n25187) );
  SDFFX1 \mem0_reg[51][4]  ( .D(n16968), .SI(\mem0[51][3] ), .SE(test_se), 
        .CLK(n1717), .Q(\mem0[51][4] ), .QN(n25188) );
  SDFFX1 \mem0_reg[51][3]  ( .D(n16967), .SI(\mem0[51][2] ), .SE(test_se), 
        .CLK(n1717), .Q(\mem0[51][3] ), .QN(n25189) );
  SDFFX1 \mem0_reg[51][2]  ( .D(n16966), .SI(\mem0[51][1] ), .SE(test_se), 
        .CLK(n1717), .Q(\mem0[51][2] ), .QN(n25190) );
  SDFFX1 \mem0_reg[51][1]  ( .D(n16965), .SI(\mem0[51][0] ), .SE(test_se), 
        .CLK(n1717), .Q(\mem0[51][1] ), .QN(n25191) );
  SDFFX1 \mem0_reg[51][0]  ( .D(n16964), .SI(\mem0[50][7] ), .SE(test_se), 
        .CLK(n1717), .Q(\mem0[51][0] ), .QN(n25192) );
  SDFFX1 \mem0_reg[50][7]  ( .D(n16963), .SI(\mem0[50][6] ), .SE(test_se), 
        .CLK(n1717), .Q(\mem0[50][7] ), .QN(n25193) );
  SDFFX1 \mem0_reg[50][6]  ( .D(n16962), .SI(\mem0[50][5] ), .SE(test_se), 
        .CLK(n1717), .Q(\mem0[50][6] ), .QN(n25194) );
  SDFFX1 \mem0_reg[50][5]  ( .D(n16961), .SI(\mem0[50][4] ), .SE(test_se), 
        .CLK(n1718), .Q(\mem0[50][5] ), .QN(n25195) );
  SDFFX1 \mem0_reg[50][4]  ( .D(n16960), .SI(\mem0[50][3] ), .SE(test_se), 
        .CLK(n1718), .Q(\mem0[50][4] ), .QN(n25196) );
  SDFFX1 \mem0_reg[50][3]  ( .D(n16959), .SI(\mem0[50][2] ), .SE(test_se), 
        .CLK(n1718), .Q(\mem0[50][3] ), .QN(n25197) );
  SDFFX1 \mem0_reg[50][2]  ( .D(n16958), .SI(\mem0[50][1] ), .SE(test_se), 
        .CLK(n1718), .Q(\mem0[50][2] ), .QN(n25198) );
  SDFFX1 \mem0_reg[50][1]  ( .D(n16957), .SI(\mem0[50][0] ), .SE(test_se), 
        .CLK(n1718), .Q(\mem0[50][1] ), .QN(n25199) );
  SDFFX1 \mem0_reg[50][0]  ( .D(n16956), .SI(\mem0[49][7] ), .SE(test_se), 
        .CLK(n1718), .Q(\mem0[50][0] ), .QN(n25200) );
  SDFFX1 \mem0_reg[49][7]  ( .D(n16955), .SI(\mem0[49][6] ), .SE(test_se), 
        .CLK(n1718), .Q(\mem0[49][7] ), .QN(n25201) );
  SDFFX1 \mem0_reg[49][6]  ( .D(n16954), .SI(\mem0[49][5] ), .SE(test_se), 
        .CLK(n1718), .Q(\mem0[49][6] ), .QN(n25202) );
  SDFFX1 \mem0_reg[49][5]  ( .D(n16953), .SI(\mem0[49][4] ), .SE(test_se), 
        .CLK(n1718), .Q(\mem0[49][5] ), .QN(n25203) );
  SDFFX1 \mem0_reg[49][4]  ( .D(n16952), .SI(\mem0[49][3] ), .SE(test_se), 
        .CLK(n1718), .Q(\mem0[49][4] ), .QN(n25204) );
  SDFFX1 \mem0_reg[49][3]  ( .D(n16951), .SI(\mem0[49][2] ), .SE(test_se), 
        .CLK(n1718), .Q(\mem0[49][3] ), .QN(n25205) );
  SDFFX1 \mem0_reg[49][2]  ( .D(n16950), .SI(\mem0[49][1] ), .SE(test_se), 
        .CLK(n1718), .Q(\mem0[49][2] ), .QN(n25206) );
  SDFFX1 \mem0_reg[49][1]  ( .D(n16949), .SI(\mem0[49][0] ), .SE(test_se), 
        .CLK(n1719), .Q(\mem0[49][1] ), .QN(n25207) );
  SDFFX1 \mem0_reg[49][0]  ( .D(n16948), .SI(\mem0[48][7] ), .SE(test_se), 
        .CLK(n1719), .Q(\mem0[49][0] ), .QN(n25208) );
  SDFFX1 \mem0_reg[48][7]  ( .D(n16947), .SI(\mem0[48][6] ), .SE(test_se), 
        .CLK(n1719), .Q(\mem0[48][7] ), .QN(n25209) );
  SDFFX1 \mem0_reg[48][6]  ( .D(n16946), .SI(\mem0[48][5] ), .SE(test_se), 
        .CLK(n1719), .Q(\mem0[48][6] ), .QN(n25210) );
  SDFFX1 \mem0_reg[48][5]  ( .D(n16945), .SI(\mem0[48][4] ), .SE(test_se), 
        .CLK(n1719), .Q(\mem0[48][5] ), .QN(n25211) );
  SDFFX1 \mem0_reg[48][4]  ( .D(n16944), .SI(\mem0[48][3] ), .SE(test_se), 
        .CLK(n1719), .Q(\mem0[48][4] ), .QN(n25212) );
  SDFFX1 \mem0_reg[48][3]  ( .D(n16943), .SI(\mem0[48][2] ), .SE(test_se), 
        .CLK(n1719), .Q(\mem0[48][3] ), .QN(n25213) );
  SDFFX1 \mem0_reg[48][2]  ( .D(n16942), .SI(\mem0[48][1] ), .SE(test_se), 
        .CLK(n1719), .Q(\mem0[48][2] ), .QN(n25214) );
  SDFFX1 \mem0_reg[48][1]  ( .D(n16941), .SI(\mem0[48][0] ), .SE(test_se), 
        .CLK(n1719), .Q(\mem0[48][1] ), .QN(n25215) );
  SDFFX1 \mem0_reg[48][0]  ( .D(n16940), .SI(\mem0[47][7] ), .SE(test_se), 
        .CLK(n1719), .Q(\mem0[48][0] ), .QN(n25216) );
  SDFFX1 \mem0_reg[47][7]  ( .D(n16939), .SI(\mem0[47][6] ), .SE(test_se), 
        .CLK(n1719), .Q(\mem0[47][7] ), .QN(n25217) );
  SDFFX1 \mem0_reg[47][6]  ( .D(n16938), .SI(\mem0[47][5] ), .SE(test_se), 
        .CLK(n1719), .Q(\mem0[47][6] ), .QN(n25218) );
  SDFFX1 \mem0_reg[47][5]  ( .D(n16937), .SI(\mem0[47][4] ), .SE(test_se), 
        .CLK(n1720), .Q(\mem0[47][5] ), .QN(n25219) );
  SDFFX1 \mem0_reg[47][4]  ( .D(n16936), .SI(\mem0[47][3] ), .SE(test_se), 
        .CLK(n1720), .Q(\mem0[47][4] ), .QN(n25220) );
  SDFFX1 \mem0_reg[47][3]  ( .D(n16935), .SI(\mem0[47][2] ), .SE(test_se), 
        .CLK(n1720), .Q(\mem0[47][3] ), .QN(n25221) );
  SDFFX1 \mem0_reg[47][2]  ( .D(n16934), .SI(\mem0[47][1] ), .SE(test_se), 
        .CLK(n1720), .Q(\mem0[47][2] ), .QN(n25222) );
  SDFFX1 \mem0_reg[47][1]  ( .D(n16933), .SI(\mem0[47][0] ), .SE(test_se), 
        .CLK(n1720), .Q(\mem0[47][1] ), .QN(n25223) );
  SDFFX1 \mem0_reg[47][0]  ( .D(n16932), .SI(\mem0[46][7] ), .SE(test_se), 
        .CLK(n1720), .Q(\mem0[47][0] ), .QN(n25224) );
  SDFFX1 \mem0_reg[46][7]  ( .D(n16931), .SI(\mem0[46][6] ), .SE(test_se), 
        .CLK(n1720), .Q(\mem0[46][7] ), .QN(n25225) );
  SDFFX1 \mem0_reg[46][6]  ( .D(n16930), .SI(\mem0[46][5] ), .SE(test_se), 
        .CLK(n1720), .Q(\mem0[46][6] ), .QN(n25226) );
  SDFFX1 \mem0_reg[46][5]  ( .D(n16929), .SI(\mem0[46][4] ), .SE(test_se), 
        .CLK(n1720), .Q(\mem0[46][5] ), .QN(n25227) );
  SDFFX1 \mem0_reg[46][4]  ( .D(n16928), .SI(\mem0[46][3] ), .SE(test_se), 
        .CLK(n1720), .Q(\mem0[46][4] ), .QN(n25228) );
  SDFFX1 \mem0_reg[46][3]  ( .D(n16927), .SI(\mem0[46][2] ), .SE(test_se), 
        .CLK(n1720), .Q(\mem0[46][3] ), .QN(n25229) );
  SDFFX1 \mem0_reg[46][2]  ( .D(n16926), .SI(\mem0[46][1] ), .SE(test_se), 
        .CLK(n1720), .Q(\mem0[46][2] ), .QN(n25230) );
  SDFFX1 \mem0_reg[46][1]  ( .D(n16925), .SI(\mem0[46][0] ), .SE(test_se), 
        .CLK(n1721), .Q(\mem0[46][1] ), .QN(n25231) );
  SDFFX1 \mem0_reg[46][0]  ( .D(n16924), .SI(\mem0[45][7] ), .SE(test_se), 
        .CLK(n1721), .Q(\mem0[46][0] ), .QN(n25232) );
  SDFFX1 \mem0_reg[45][7]  ( .D(n16923), .SI(\mem0[45][6] ), .SE(test_se), 
        .CLK(n1721), .Q(\mem0[45][7] ), .QN(n25233) );
  SDFFX1 \mem0_reg[45][6]  ( .D(n16922), .SI(\mem0[45][5] ), .SE(test_se), 
        .CLK(n1721), .Q(\mem0[45][6] ), .QN(n25234) );
  SDFFX1 \mem0_reg[45][5]  ( .D(n16921), .SI(\mem0[45][4] ), .SE(test_se), 
        .CLK(n1721), .Q(\mem0[45][5] ), .QN(n25235) );
  SDFFX1 \mem0_reg[45][4]  ( .D(n16920), .SI(\mem0[45][3] ), .SE(test_se), 
        .CLK(n1721), .Q(\mem0[45][4] ), .QN(n25236) );
  SDFFX1 \mem0_reg[45][3]  ( .D(n16919), .SI(\mem0[45][2] ), .SE(test_se), 
        .CLK(n1721), .Q(\mem0[45][3] ), .QN(n25237) );
  SDFFX1 \mem0_reg[45][2]  ( .D(n16918), .SI(\mem0[45][1] ), .SE(test_se), 
        .CLK(n1721), .Q(\mem0[45][2] ), .QN(n25238) );
  SDFFX1 \mem0_reg[45][1]  ( .D(n16917), .SI(\mem0[45][0] ), .SE(test_se), 
        .CLK(n1721), .Q(\mem0[45][1] ), .QN(n25239) );
  SDFFX1 \mem0_reg[45][0]  ( .D(n16916), .SI(\mem0[44][7] ), .SE(test_se), 
        .CLK(n1721), .Q(\mem0[45][0] ), .QN(n25240) );
  SDFFX1 \mem0_reg[44][7]  ( .D(n16915), .SI(\mem0[44][6] ), .SE(test_se), 
        .CLK(n1721), .Q(\mem0[44][7] ), .QN(n25241) );
  SDFFX1 \mem0_reg[44][6]  ( .D(n16914), .SI(\mem0[44][5] ), .SE(test_se), 
        .CLK(n1721), .Q(\mem0[44][6] ), .QN(n25242) );
  SDFFX1 \mem0_reg[44][5]  ( .D(n16913), .SI(\mem0[44][4] ), .SE(test_se), 
        .CLK(n1722), .Q(\mem0[44][5] ), .QN(n25243) );
  SDFFX1 \mem0_reg[44][4]  ( .D(n16912), .SI(\mem0[44][3] ), .SE(test_se), 
        .CLK(n1722), .Q(\mem0[44][4] ), .QN(n25244) );
  SDFFX1 \mem0_reg[44][3]  ( .D(n16911), .SI(\mem0[44][2] ), .SE(test_se), 
        .CLK(n1722), .Q(\mem0[44][3] ), .QN(n25245) );
  SDFFX1 \mem0_reg[44][2]  ( .D(n16910), .SI(\mem0[44][1] ), .SE(test_se), 
        .CLK(n1722), .Q(\mem0[44][2] ), .QN(n25246) );
  SDFFX1 \mem0_reg[44][1]  ( .D(n16909), .SI(\mem0[44][0] ), .SE(test_se), 
        .CLK(n1722), .Q(\mem0[44][1] ), .QN(n25247) );
  SDFFX1 \mem0_reg[44][0]  ( .D(n16908), .SI(\mem0[43][7] ), .SE(test_se), 
        .CLK(n1722), .Q(\mem0[44][0] ), .QN(n25248) );
  SDFFX1 \mem0_reg[43][7]  ( .D(n16907), .SI(\mem0[43][6] ), .SE(test_se), 
        .CLK(n1722), .Q(\mem0[43][7] ), .QN(n25249) );
  SDFFX1 \mem0_reg[43][6]  ( .D(n16906), .SI(\mem0[43][5] ), .SE(test_se), 
        .CLK(n1722), .Q(\mem0[43][6] ), .QN(n25250) );
  SDFFX1 \mem0_reg[43][5]  ( .D(n16905), .SI(\mem0[43][4] ), .SE(test_se), 
        .CLK(n1722), .Q(\mem0[43][5] ), .QN(n25251) );
  SDFFX1 \mem0_reg[43][4]  ( .D(n16904), .SI(\mem0[43][3] ), .SE(test_se), 
        .CLK(n1722), .Q(\mem0[43][4] ), .QN(n25252) );
  SDFFX1 \mem0_reg[43][3]  ( .D(n16903), .SI(\mem0[43][2] ), .SE(test_se), 
        .CLK(n1722), .Q(\mem0[43][3] ), .QN(n25253) );
  SDFFX1 \mem0_reg[43][2]  ( .D(n16902), .SI(\mem0[43][1] ), .SE(test_se), 
        .CLK(n1722), .Q(\mem0[43][2] ), .QN(n25254) );
  SDFFX1 \mem0_reg[43][1]  ( .D(n16901), .SI(\mem0[43][0] ), .SE(test_se), 
        .CLK(n1723), .Q(\mem0[43][1] ), .QN(n25255) );
  SDFFX1 \mem0_reg[43][0]  ( .D(n16900), .SI(\mem0[42][7] ), .SE(test_se), 
        .CLK(n1723), .Q(\mem0[43][0] ), .QN(n25256) );
  SDFFX1 \mem0_reg[42][7]  ( .D(n16899), .SI(\mem0[42][6] ), .SE(test_se), 
        .CLK(n1723), .Q(\mem0[42][7] ), .QN(n25257) );
  SDFFX1 \mem0_reg[42][6]  ( .D(n16898), .SI(\mem0[42][5] ), .SE(test_se), 
        .CLK(n1723), .Q(\mem0[42][6] ), .QN(n25258) );
  SDFFX1 \mem0_reg[42][5]  ( .D(n16897), .SI(\mem0[42][4] ), .SE(test_se), 
        .CLK(n1723), .Q(\mem0[42][5] ), .QN(n25259) );
  SDFFX1 \mem0_reg[42][4]  ( .D(n16896), .SI(\mem0[42][3] ), .SE(test_se), 
        .CLK(n1723), .Q(\mem0[42][4] ), .QN(n25260) );
  SDFFX1 \mem0_reg[42][3]  ( .D(n16895), .SI(\mem0[42][2] ), .SE(test_se), 
        .CLK(n1723), .Q(\mem0[42][3] ), .QN(n25261) );
  SDFFX1 \mem0_reg[42][2]  ( .D(n16894), .SI(\mem0[42][1] ), .SE(test_se), 
        .CLK(n1723), .Q(\mem0[42][2] ), .QN(n25262) );
  SDFFX1 \mem0_reg[42][1]  ( .D(n16893), .SI(\mem0[42][0] ), .SE(test_se), 
        .CLK(n1723), .Q(\mem0[42][1] ), .QN(n25263) );
  SDFFX1 \mem0_reg[42][0]  ( .D(n16892), .SI(\mem0[41][7] ), .SE(test_se), 
        .CLK(n1723), .Q(\mem0[42][0] ), .QN(n25264) );
  SDFFX1 \mem0_reg[41][7]  ( .D(n16891), .SI(\mem0[41][6] ), .SE(test_se), 
        .CLK(n1723), .Q(\mem0[41][7] ), .QN(n25265) );
  SDFFX1 \mem0_reg[41][6]  ( .D(n16890), .SI(\mem0[41][5] ), .SE(test_se), 
        .CLK(n1723), .Q(\mem0[41][6] ), .QN(n25266) );
  SDFFX1 \mem0_reg[41][5]  ( .D(n16889), .SI(\mem0[41][4] ), .SE(test_se), 
        .CLK(n1724), .Q(\mem0[41][5] ), .QN(n25267) );
  SDFFX1 \mem0_reg[41][4]  ( .D(n16888), .SI(\mem0[41][3] ), .SE(test_se), 
        .CLK(n1724), .Q(\mem0[41][4] ), .QN(n25268) );
  SDFFX1 \mem0_reg[41][3]  ( .D(n16887), .SI(\mem0[41][2] ), .SE(test_se), 
        .CLK(n1724), .Q(\mem0[41][3] ), .QN(n25269) );
  SDFFX1 \mem0_reg[41][2]  ( .D(n16886), .SI(\mem0[41][1] ), .SE(test_se), 
        .CLK(n1724), .Q(\mem0[41][2] ), .QN(n25270) );
  SDFFX1 \mem0_reg[41][1]  ( .D(n16885), .SI(\mem0[41][0] ), .SE(test_se), 
        .CLK(n1724), .Q(\mem0[41][1] ), .QN(n25271) );
  SDFFX1 \mem0_reg[41][0]  ( .D(n16884), .SI(\mem0[40][7] ), .SE(test_se), 
        .CLK(n1724), .Q(\mem0[41][0] ), .QN(n25272) );
  SDFFX1 \mem0_reg[40][7]  ( .D(n16883), .SI(\mem0[40][6] ), .SE(test_se), 
        .CLK(n1724), .Q(\mem0[40][7] ), .QN(n25273) );
  SDFFX1 \mem0_reg[40][6]  ( .D(n16882), .SI(\mem0[40][5] ), .SE(test_se), 
        .CLK(n1724), .Q(\mem0[40][6] ), .QN(n25274) );
  SDFFX1 \mem0_reg[40][5]  ( .D(n16881), .SI(\mem0[40][4] ), .SE(test_se), 
        .CLK(n1724), .Q(\mem0[40][5] ), .QN(n25275) );
  SDFFX1 \mem0_reg[40][4]  ( .D(n16880), .SI(\mem0[40][3] ), .SE(test_se), 
        .CLK(n1724), .Q(\mem0[40][4] ), .QN(n25276) );
  SDFFX1 \mem0_reg[40][3]  ( .D(n16879), .SI(\mem0[40][2] ), .SE(test_se), 
        .CLK(n1724), .Q(\mem0[40][3] ), .QN(n25277) );
  SDFFX1 \mem0_reg[40][2]  ( .D(n16878), .SI(\mem0[40][1] ), .SE(test_se), 
        .CLK(n1724), .Q(\mem0[40][2] ), .QN(n25278) );
  SDFFX1 \mem0_reg[40][1]  ( .D(n16877), .SI(\mem0[40][0] ), .SE(test_se), 
        .CLK(n1725), .Q(\mem0[40][1] ), .QN(n25279) );
  SDFFX1 \mem0_reg[40][0]  ( .D(n16876), .SI(\mem0[39][7] ), .SE(test_se), 
        .CLK(n1725), .Q(\mem0[40][0] ), .QN(n25280) );
  SDFFX1 \mem0_reg[39][7]  ( .D(n16875), .SI(\mem0[39][6] ), .SE(test_se), 
        .CLK(n1725), .Q(\mem0[39][7] ), .QN(n25281) );
  SDFFX1 \mem0_reg[39][6]  ( .D(n16874), .SI(\mem0[39][5] ), .SE(test_se), 
        .CLK(n1725), .Q(\mem0[39][6] ), .QN(n25282) );
  SDFFX1 \mem0_reg[39][5]  ( .D(n16873), .SI(\mem0[39][4] ), .SE(test_se), 
        .CLK(n1725), .Q(\mem0[39][5] ), .QN(n25283) );
  SDFFX1 \mem0_reg[39][4]  ( .D(n16872), .SI(\mem0[39][3] ), .SE(test_se), 
        .CLK(n1725), .Q(\mem0[39][4] ), .QN(n25284) );
  SDFFX1 \mem0_reg[39][3]  ( .D(n16871), .SI(\mem0[39][2] ), .SE(test_se), 
        .CLK(n1725), .Q(\mem0[39][3] ), .QN(n25285) );
  SDFFX1 \mem0_reg[39][2]  ( .D(n16870), .SI(\mem0[39][1] ), .SE(test_se), 
        .CLK(n1725), .Q(\mem0[39][2] ), .QN(n25286) );
  SDFFX1 \mem0_reg[39][1]  ( .D(n16869), .SI(\mem0[39][0] ), .SE(test_se), 
        .CLK(n1725), .Q(\mem0[39][1] ), .QN(n25287) );
  SDFFX1 \mem0_reg[39][0]  ( .D(n16868), .SI(\mem0[38][7] ), .SE(test_se), 
        .CLK(n1725), .Q(\mem0[39][0] ), .QN(n25288) );
  SDFFX1 \mem0_reg[38][7]  ( .D(n16867), .SI(\mem0[38][6] ), .SE(test_se), 
        .CLK(n1725), .Q(\mem0[38][7] ), .QN(n25289) );
  SDFFX1 \mem0_reg[38][6]  ( .D(n16866), .SI(\mem0[38][5] ), .SE(test_se), 
        .CLK(n1725), .Q(\mem0[38][6] ), .QN(n25290) );
  SDFFX1 \mem0_reg[38][5]  ( .D(n16865), .SI(\mem0[38][4] ), .SE(test_se), 
        .CLK(n1726), .Q(\mem0[38][5] ), .QN(n25291) );
  SDFFX1 \mem0_reg[38][4]  ( .D(n16864), .SI(\mem0[38][3] ), .SE(test_se), 
        .CLK(n1726), .Q(\mem0[38][4] ), .QN(n25292) );
  SDFFX1 \mem0_reg[38][3]  ( .D(n16863), .SI(\mem0[38][2] ), .SE(test_se), 
        .CLK(n1726), .Q(\mem0[38][3] ), .QN(n25293) );
  SDFFX1 \mem0_reg[38][2]  ( .D(n16862), .SI(\mem0[38][1] ), .SE(test_se), 
        .CLK(n1726), .Q(\mem0[38][2] ), .QN(n25294) );
  SDFFX1 \mem0_reg[38][1]  ( .D(n16861), .SI(\mem0[38][0] ), .SE(test_se), 
        .CLK(n1726), .Q(\mem0[38][1] ), .QN(n25295) );
  SDFFX1 \mem0_reg[38][0]  ( .D(n16860), .SI(\mem0[37][7] ), .SE(test_se), 
        .CLK(n1726), .Q(\mem0[38][0] ), .QN(n25296) );
  SDFFX1 \mem0_reg[37][7]  ( .D(n16859), .SI(\mem0[37][6] ), .SE(test_se), 
        .CLK(n1726), .Q(\mem0[37][7] ), .QN(n25297) );
  SDFFX1 \mem0_reg[37][6]  ( .D(n16858), .SI(\mem0[37][5] ), .SE(test_se), 
        .CLK(n1726), .Q(\mem0[37][6] ), .QN(n25298) );
  SDFFX1 \mem0_reg[37][5]  ( .D(n16857), .SI(\mem0[37][4] ), .SE(test_se), 
        .CLK(n1726), .Q(\mem0[37][5] ), .QN(n25299) );
  SDFFX1 \mem0_reg[37][4]  ( .D(n16856), .SI(\mem0[37][3] ), .SE(test_se), 
        .CLK(n1726), .Q(\mem0[37][4] ), .QN(n25300) );
  SDFFX1 \mem0_reg[37][3]  ( .D(n16855), .SI(\mem0[37][2] ), .SE(test_se), 
        .CLK(n1726), .Q(\mem0[37][3] ), .QN(n25301) );
  SDFFX1 \mem0_reg[37][2]  ( .D(n16854), .SI(\mem0[37][1] ), .SE(test_se), 
        .CLK(n1726), .Q(\mem0[37][2] ), .QN(n25302) );
  SDFFX1 \mem0_reg[37][1]  ( .D(n16853), .SI(\mem0[37][0] ), .SE(test_se), 
        .CLK(n1727), .Q(\mem0[37][1] ), .QN(n25303) );
  SDFFX1 \mem0_reg[37][0]  ( .D(n16852), .SI(\mem0[36][7] ), .SE(test_se), 
        .CLK(n1727), .Q(\mem0[37][0] ), .QN(n25304) );
  SDFFX1 \mem0_reg[36][7]  ( .D(n16851), .SI(\mem0[36][6] ), .SE(test_se), 
        .CLK(n1727), .Q(\mem0[36][7] ), .QN(n25305) );
  SDFFX1 \mem0_reg[36][6]  ( .D(n16850), .SI(\mem0[36][5] ), .SE(test_se), 
        .CLK(n1727), .Q(\mem0[36][6] ), .QN(n25306) );
  SDFFX1 \mem0_reg[36][5]  ( .D(n16849), .SI(\mem0[36][4] ), .SE(test_se), 
        .CLK(n1727), .Q(\mem0[36][5] ), .QN(n25307) );
  SDFFX1 \mem0_reg[36][4]  ( .D(n16848), .SI(\mem0[36][3] ), .SE(test_se), 
        .CLK(n1727), .Q(\mem0[36][4] ), .QN(n25308) );
  SDFFX1 \mem0_reg[36][3]  ( .D(n16847), .SI(\mem0[36][2] ), .SE(test_se), 
        .CLK(n1727), .Q(\mem0[36][3] ), .QN(n25309) );
  SDFFX1 \mem0_reg[36][2]  ( .D(n16846), .SI(\mem0[36][1] ), .SE(test_se), 
        .CLK(n1727), .Q(\mem0[36][2] ), .QN(n25310) );
  SDFFX1 \mem0_reg[36][1]  ( .D(n16845), .SI(\mem0[36][0] ), .SE(test_se), 
        .CLK(n1727), .Q(\mem0[36][1] ), .QN(n25311) );
  SDFFX1 \mem0_reg[36][0]  ( .D(n16844), .SI(\mem0[35][7] ), .SE(test_se), 
        .CLK(n1727), .Q(\mem0[36][0] ), .QN(n25312) );
  SDFFX1 \mem0_reg[35][7]  ( .D(n16843), .SI(\mem0[35][6] ), .SE(test_se), 
        .CLK(n1727), .Q(\mem0[35][7] ), .QN(n25313) );
  SDFFX1 \mem0_reg[35][6]  ( .D(n16842), .SI(\mem0[35][5] ), .SE(test_se), 
        .CLK(n1727), .Q(\mem0[35][6] ), .QN(n25314) );
  SDFFX1 \mem0_reg[35][5]  ( .D(n16841), .SI(\mem0[35][4] ), .SE(test_se), 
        .CLK(n1728), .Q(\mem0[35][5] ), .QN(n25315) );
  SDFFX1 \mem0_reg[35][4]  ( .D(n16840), .SI(\mem0[35][3] ), .SE(test_se), 
        .CLK(n1728), .Q(\mem0[35][4] ), .QN(n25316) );
  SDFFX1 \mem0_reg[35][3]  ( .D(n16839), .SI(\mem0[35][2] ), .SE(test_se), 
        .CLK(n1728), .Q(\mem0[35][3] ), .QN(n25317) );
  SDFFX1 \mem0_reg[35][2]  ( .D(n16838), .SI(\mem0[35][1] ), .SE(test_se), 
        .CLK(n1728), .Q(\mem0[35][2] ), .QN(n25318) );
  SDFFX1 \mem0_reg[35][1]  ( .D(n16837), .SI(\mem0[35][0] ), .SE(test_se), 
        .CLK(n1728), .Q(\mem0[35][1] ), .QN(n25319) );
  SDFFX1 \mem0_reg[35][0]  ( .D(n16836), .SI(\mem0[34][7] ), .SE(test_se), 
        .CLK(n1728), .Q(\mem0[35][0] ), .QN(n25320) );
  SDFFX1 \mem0_reg[34][7]  ( .D(n16835), .SI(\mem0[34][6] ), .SE(test_se), 
        .CLK(n1728), .Q(\mem0[34][7] ), .QN(n25321) );
  SDFFX1 \mem0_reg[34][6]  ( .D(n16834), .SI(\mem0[34][5] ), .SE(test_se), 
        .CLK(n1728), .Q(\mem0[34][6] ), .QN(n25322) );
  SDFFX1 \mem0_reg[34][5]  ( .D(n16833), .SI(\mem0[34][4] ), .SE(test_se), 
        .CLK(n1728), .Q(\mem0[34][5] ), .QN(n25323) );
  SDFFX1 \mem0_reg[34][4]  ( .D(n16832), .SI(\mem0[34][3] ), .SE(test_se), 
        .CLK(n1728), .Q(\mem0[34][4] ), .QN(n25324) );
  SDFFX1 \mem0_reg[34][3]  ( .D(n16831), .SI(\mem0[34][2] ), .SE(test_se), 
        .CLK(n1728), .Q(\mem0[34][3] ), .QN(n25325) );
  SDFFX1 \mem0_reg[34][2]  ( .D(n16830), .SI(\mem0[34][1] ), .SE(test_se), 
        .CLK(n1728), .Q(\mem0[34][2] ), .QN(n25326) );
  SDFFX1 \mem0_reg[34][1]  ( .D(n16829), .SI(\mem0[34][0] ), .SE(test_se), 
        .CLK(n1729), .Q(\mem0[34][1] ), .QN(n25327) );
  SDFFX1 \mem0_reg[34][0]  ( .D(n16828), .SI(\mem0[33][7] ), .SE(test_se), 
        .CLK(n1729), .Q(\mem0[34][0] ), .QN(n25328) );
  SDFFX1 \mem0_reg[33][7]  ( .D(n16827), .SI(\mem0[33][6] ), .SE(test_se), 
        .CLK(n1729), .Q(\mem0[33][7] ), .QN(n25329) );
  SDFFX1 \mem0_reg[33][6]  ( .D(n16826), .SI(\mem0[33][5] ), .SE(test_se), 
        .CLK(n1729), .Q(\mem0[33][6] ), .QN(n25330) );
  SDFFX1 \mem0_reg[33][5]  ( .D(n16825), .SI(\mem0[33][4] ), .SE(test_se), 
        .CLK(n1729), .Q(\mem0[33][5] ), .QN(n25331) );
  SDFFX1 \mem0_reg[33][4]  ( .D(n16824), .SI(\mem0[33][3] ), .SE(test_se), 
        .CLK(n1729), .Q(\mem0[33][4] ), .QN(n25332) );
  SDFFX1 \mem0_reg[33][3]  ( .D(n16823), .SI(\mem0[33][2] ), .SE(test_se), 
        .CLK(n1729), .Q(\mem0[33][3] ), .QN(n25333) );
  SDFFX1 \mem0_reg[33][2]  ( .D(n16822), .SI(\mem0[33][1] ), .SE(test_se), 
        .CLK(n1729), .Q(\mem0[33][2] ), .QN(n25334) );
  SDFFX1 \mem0_reg[33][1]  ( .D(n16821), .SI(\mem0[33][0] ), .SE(test_se), 
        .CLK(n1729), .Q(\mem0[33][1] ), .QN(n25335) );
  SDFFX1 \mem0_reg[33][0]  ( .D(n16820), .SI(\mem0[32][7] ), .SE(test_se), 
        .CLK(n1729), .Q(\mem0[33][0] ), .QN(n25336) );
  SDFFX1 \mem0_reg[32][7]  ( .D(n16819), .SI(\mem0[32][6] ), .SE(test_se), 
        .CLK(n1729), .Q(\mem0[32][7] ), .QN(n25337) );
  SDFFX1 \mem0_reg[32][6]  ( .D(n16818), .SI(\mem0[32][5] ), .SE(test_se), 
        .CLK(n1729), .Q(\mem0[32][6] ), .QN(n25338) );
  SDFFX1 \mem0_reg[32][5]  ( .D(n16817), .SI(\mem0[32][4] ), .SE(test_se), 
        .CLK(n1730), .Q(\mem0[32][5] ), .QN(n25339) );
  SDFFX1 \mem0_reg[32][4]  ( .D(n16816), .SI(\mem0[32][3] ), .SE(test_se), 
        .CLK(n1730), .Q(\mem0[32][4] ), .QN(n25340) );
  SDFFX1 \mem0_reg[32][3]  ( .D(n16815), .SI(\mem0[32][2] ), .SE(test_se), 
        .CLK(n1730), .Q(\mem0[32][3] ), .QN(n25341) );
  SDFFX1 \mem0_reg[32][2]  ( .D(n16814), .SI(\mem0[32][1] ), .SE(test_se), 
        .CLK(n1730), .Q(\mem0[32][2] ), .QN(n25342) );
  SDFFX1 \mem0_reg[32][1]  ( .D(n16813), .SI(\mem0[32][0] ), .SE(test_se), 
        .CLK(n1730), .Q(\mem0[32][1] ), .QN(n25343) );
  SDFFX1 \mem0_reg[32][0]  ( .D(n16812), .SI(\mem0[31][7] ), .SE(test_se), 
        .CLK(n1730), .Q(\mem0[32][0] ), .QN(n25344) );
  SDFFX1 \mem0_reg[31][7]  ( .D(n16811), .SI(\mem0[31][6] ), .SE(test_se), 
        .CLK(n1730), .Q(\mem0[31][7] ), .QN(n25345) );
  SDFFX1 \mem0_reg[31][6]  ( .D(n16810), .SI(\mem0[31][5] ), .SE(test_se), 
        .CLK(n1730), .Q(\mem0[31][6] ), .QN(n25346) );
  SDFFX1 \mem0_reg[31][5]  ( .D(n16809), .SI(\mem0[31][4] ), .SE(test_se), 
        .CLK(n1730), .Q(\mem0[31][5] ), .QN(n25347) );
  SDFFX1 \mem0_reg[31][4]  ( .D(n16808), .SI(\mem0[31][3] ), .SE(test_se), 
        .CLK(n1730), .Q(\mem0[31][4] ), .QN(n25348) );
  SDFFX1 \mem0_reg[31][3]  ( .D(n16807), .SI(\mem0[31][2] ), .SE(test_se), 
        .CLK(n1730), .Q(\mem0[31][3] ), .QN(n25349) );
  SDFFX1 \mem0_reg[31][2]  ( .D(n16806), .SI(\mem0[31][1] ), .SE(test_se), 
        .CLK(n1730), .Q(\mem0[31][2] ), .QN(n25350) );
  SDFFX1 \mem0_reg[31][1]  ( .D(n16805), .SI(\mem0[31][0] ), .SE(test_se), 
        .CLK(n1731), .Q(\mem0[31][1] ), .QN(n25351) );
  SDFFX1 \mem0_reg[31][0]  ( .D(n16804), .SI(\mem0[30][7] ), .SE(test_se), 
        .CLK(n1731), .Q(\mem0[31][0] ), .QN(n25352) );
  SDFFX1 \mem0_reg[30][7]  ( .D(n16803), .SI(\mem0[30][6] ), .SE(test_se), 
        .CLK(n1731), .Q(\mem0[30][7] ), .QN(n25353) );
  SDFFX1 \mem0_reg[30][6]  ( .D(n16802), .SI(\mem0[30][5] ), .SE(test_se), 
        .CLK(n1731), .Q(\mem0[30][6] ), .QN(n25354) );
  SDFFX1 \mem0_reg[30][5]  ( .D(n16801), .SI(\mem0[30][4] ), .SE(test_se), 
        .CLK(n1731), .Q(\mem0[30][5] ), .QN(n25355) );
  SDFFX1 \mem0_reg[30][4]  ( .D(n16800), .SI(\mem0[30][3] ), .SE(test_se), 
        .CLK(n1731), .Q(\mem0[30][4] ), .QN(n25356) );
  SDFFX1 \mem0_reg[30][3]  ( .D(n16799), .SI(\mem0[30][2] ), .SE(test_se), 
        .CLK(n1731), .Q(\mem0[30][3] ), .QN(n25357) );
  SDFFX1 \mem0_reg[30][2]  ( .D(n16798), .SI(\mem0[30][1] ), .SE(test_se), 
        .CLK(n1731), .Q(\mem0[30][2] ), .QN(n25358) );
  SDFFX1 \mem0_reg[30][1]  ( .D(n16797), .SI(\mem0[30][0] ), .SE(test_se), 
        .CLK(n1731), .Q(\mem0[30][1] ), .QN(n25359) );
  SDFFX1 \mem0_reg[30][0]  ( .D(n16796), .SI(\mem0[29][7] ), .SE(test_se), 
        .CLK(n1731), .Q(\mem0[30][0] ), .QN(n25360) );
  SDFFX1 \mem0_reg[29][7]  ( .D(n16795), .SI(\mem0[29][6] ), .SE(test_se), 
        .CLK(n1731), .Q(\mem0[29][7] ), .QN(n25361) );
  SDFFX1 \mem0_reg[29][6]  ( .D(n16794), .SI(\mem0[29][5] ), .SE(test_se), 
        .CLK(n1731), .Q(\mem0[29][6] ), .QN(n25362) );
  SDFFX1 \mem0_reg[29][5]  ( .D(n16793), .SI(\mem0[29][4] ), .SE(test_se), 
        .CLK(n1732), .Q(\mem0[29][5] ), .QN(n25363) );
  SDFFX1 \mem0_reg[29][4]  ( .D(n16792), .SI(\mem0[29][3] ), .SE(test_se), 
        .CLK(n1732), .Q(\mem0[29][4] ), .QN(n25364) );
  SDFFX1 \mem0_reg[29][3]  ( .D(n16791), .SI(\mem0[29][2] ), .SE(test_se), 
        .CLK(n1732), .Q(\mem0[29][3] ), .QN(n25365) );
  SDFFX1 \mem0_reg[29][2]  ( .D(n16790), .SI(\mem0[29][1] ), .SE(test_se), 
        .CLK(n1732), .Q(\mem0[29][2] ), .QN(n25366) );
  SDFFX1 \mem0_reg[29][1]  ( .D(n16789), .SI(\mem0[29][0] ), .SE(test_se), 
        .CLK(n1732), .Q(\mem0[29][1] ), .QN(n25367) );
  SDFFX1 \mem0_reg[29][0]  ( .D(n16788), .SI(\mem0[28][7] ), .SE(test_se), 
        .CLK(n1732), .Q(\mem0[29][0] ), .QN(n25368) );
  SDFFX1 \mem0_reg[28][7]  ( .D(n16787), .SI(\mem0[28][6] ), .SE(test_se), 
        .CLK(n1732), .Q(\mem0[28][7] ), .QN(n25369) );
  SDFFX1 \mem0_reg[28][6]  ( .D(n16786), .SI(\mem0[28][5] ), .SE(test_se), 
        .CLK(n1732), .Q(\mem0[28][6] ), .QN(n25370) );
  SDFFX1 \mem0_reg[28][5]  ( .D(n16785), .SI(\mem0[28][4] ), .SE(test_se), 
        .CLK(n1732), .Q(\mem0[28][5] ), .QN(n25371) );
  SDFFX1 \mem0_reg[28][4]  ( .D(n16784), .SI(\mem0[28][3] ), .SE(test_se), 
        .CLK(n1732), .Q(\mem0[28][4] ), .QN(n25372) );
  SDFFX1 \mem0_reg[28][3]  ( .D(n16783), .SI(\mem0[28][2] ), .SE(test_se), 
        .CLK(n1732), .Q(\mem0[28][3] ), .QN(n25373) );
  SDFFX1 \mem0_reg[28][2]  ( .D(n16782), .SI(\mem0[28][1] ), .SE(test_se), 
        .CLK(n1732), .Q(\mem0[28][2] ), .QN(n25374) );
  SDFFX1 \mem0_reg[28][1]  ( .D(n16781), .SI(\mem0[28][0] ), .SE(test_se), 
        .CLK(n1733), .Q(\mem0[28][1] ), .QN(n25375) );
  SDFFX1 \mem0_reg[28][0]  ( .D(n16780), .SI(\mem0[27][7] ), .SE(test_se), 
        .CLK(n1733), .Q(\mem0[28][0] ), .QN(n25376) );
  SDFFX1 \mem0_reg[27][7]  ( .D(n16779), .SI(\mem0[27][6] ), .SE(test_se), 
        .CLK(n1733), .Q(\mem0[27][7] ), .QN(n25377) );
  SDFFX1 \mem0_reg[27][6]  ( .D(n16778), .SI(\mem0[27][5] ), .SE(test_se), 
        .CLK(n1733), .Q(\mem0[27][6] ), .QN(n25378) );
  SDFFX1 \mem0_reg[27][5]  ( .D(n16777), .SI(\mem0[27][4] ), .SE(test_se), 
        .CLK(n1733), .Q(\mem0[27][5] ), .QN(n25379) );
  SDFFX1 \mem0_reg[27][4]  ( .D(n16776), .SI(\mem0[27][3] ), .SE(test_se), 
        .CLK(n1733), .Q(\mem0[27][4] ), .QN(n25380) );
  SDFFX1 \mem0_reg[27][3]  ( .D(n16775), .SI(\mem0[27][2] ), .SE(test_se), 
        .CLK(n1733), .Q(\mem0[27][3] ), .QN(n25381) );
  SDFFX1 \mem0_reg[27][2]  ( .D(n16774), .SI(\mem0[27][1] ), .SE(test_se), 
        .CLK(n1733), .Q(\mem0[27][2] ), .QN(n25382) );
  SDFFX1 \mem0_reg[27][1]  ( .D(n16773), .SI(\mem0[27][0] ), .SE(test_se), 
        .CLK(n1733), .Q(\mem0[27][1] ), .QN(n25383) );
  SDFFX1 \mem0_reg[27][0]  ( .D(n16772), .SI(\mem0[26][7] ), .SE(test_se), 
        .CLK(n1733), .Q(\mem0[27][0] ), .QN(n25384) );
  SDFFX1 \mem0_reg[26][7]  ( .D(n16771), .SI(\mem0[26][6] ), .SE(test_se), 
        .CLK(n1733), .Q(\mem0[26][7] ), .QN(n25385) );
  SDFFX1 \mem0_reg[26][6]  ( .D(n16770), .SI(\mem0[26][5] ), .SE(test_se), 
        .CLK(n1733), .Q(\mem0[26][6] ), .QN(n25386) );
  SDFFX1 \mem0_reg[26][5]  ( .D(n16769), .SI(\mem0[26][4] ), .SE(test_se), 
        .CLK(n1734), .Q(\mem0[26][5] ), .QN(n25387) );
  SDFFX1 \mem0_reg[26][4]  ( .D(n16768), .SI(\mem0[26][3] ), .SE(test_se), 
        .CLK(n1734), .Q(\mem0[26][4] ), .QN(n25388) );
  SDFFX1 \mem0_reg[26][3]  ( .D(n16767), .SI(\mem0[26][2] ), .SE(test_se), 
        .CLK(n1734), .Q(\mem0[26][3] ), .QN(n25389) );
  SDFFX1 \mem0_reg[26][2]  ( .D(n16766), .SI(\mem0[26][1] ), .SE(test_se), 
        .CLK(n1734), .Q(\mem0[26][2] ), .QN(n25390) );
  SDFFX1 \mem0_reg[26][1]  ( .D(n16765), .SI(\mem0[26][0] ), .SE(test_se), 
        .CLK(n1734), .Q(\mem0[26][1] ), .QN(n25391) );
  SDFFX1 \mem0_reg[26][0]  ( .D(n16764), .SI(\mem0[25][7] ), .SE(test_se), 
        .CLK(n1734), .Q(\mem0[26][0] ), .QN(n25392) );
  SDFFX1 \mem0_reg[25][7]  ( .D(n16763), .SI(\mem0[25][6] ), .SE(test_se), 
        .CLK(n1734), .Q(\mem0[25][7] ), .QN(n25393) );
  SDFFX1 \mem0_reg[25][6]  ( .D(n16762), .SI(\mem0[25][5] ), .SE(test_se), 
        .CLK(n1734), .Q(\mem0[25][6] ), .QN(n25394) );
  SDFFX1 \mem0_reg[25][5]  ( .D(n16761), .SI(\mem0[25][4] ), .SE(test_se), 
        .CLK(n1734), .Q(\mem0[25][5] ), .QN(n25395) );
  SDFFX1 \mem0_reg[25][4]  ( .D(n16760), .SI(\mem0[25][3] ), .SE(test_se), 
        .CLK(n1734), .Q(\mem0[25][4] ), .QN(n25396) );
  SDFFX1 \mem0_reg[25][3]  ( .D(n16759), .SI(\mem0[25][2] ), .SE(test_se), 
        .CLK(n1734), .Q(\mem0[25][3] ), .QN(n25397) );
  SDFFX1 \mem0_reg[25][2]  ( .D(n16758), .SI(\mem0[25][1] ), .SE(test_se), 
        .CLK(n1734), .Q(\mem0[25][2] ), .QN(n25398) );
  SDFFX1 \mem0_reg[25][1]  ( .D(n16757), .SI(\mem0[25][0] ), .SE(test_se), 
        .CLK(n1735), .Q(\mem0[25][1] ), .QN(n25399) );
  SDFFX1 \mem0_reg[25][0]  ( .D(n16756), .SI(\mem0[24][7] ), .SE(test_se), 
        .CLK(n1735), .Q(\mem0[25][0] ), .QN(n25400) );
  SDFFX1 \mem0_reg[24][7]  ( .D(n16755), .SI(\mem0[24][6] ), .SE(test_se), 
        .CLK(n1735), .Q(\mem0[24][7] ), .QN(n25401) );
  SDFFX1 \mem0_reg[24][6]  ( .D(n16754), .SI(\mem0[24][5] ), .SE(test_se), 
        .CLK(n1735), .Q(\mem0[24][6] ), .QN(n25402) );
  SDFFX1 \mem0_reg[24][5]  ( .D(n16753), .SI(\mem0[24][4] ), .SE(test_se), 
        .CLK(n1735), .Q(\mem0[24][5] ), .QN(n25403) );
  SDFFX1 \mem0_reg[24][4]  ( .D(n16752), .SI(\mem0[24][3] ), .SE(test_se), 
        .CLK(n1735), .Q(\mem0[24][4] ), .QN(n25404) );
  SDFFX1 \mem0_reg[24][3]  ( .D(n16751), .SI(\mem0[24][2] ), .SE(test_se), 
        .CLK(n1735), .Q(\mem0[24][3] ), .QN(n25405) );
  SDFFX1 \mem0_reg[24][2]  ( .D(n16750), .SI(\mem0[24][1] ), .SE(test_se), 
        .CLK(n1735), .Q(\mem0[24][2] ), .QN(n25406) );
  SDFFX1 \mem0_reg[24][1]  ( .D(n16749), .SI(\mem0[24][0] ), .SE(test_se), 
        .CLK(n1735), .Q(\mem0[24][1] ), .QN(n25407) );
  SDFFX1 \mem0_reg[24][0]  ( .D(n16748), .SI(\mem0[23][7] ), .SE(test_se), 
        .CLK(n1735), .Q(\mem0[24][0] ), .QN(n25408) );
  SDFFX1 \mem0_reg[23][7]  ( .D(n16747), .SI(\mem0[23][6] ), .SE(test_se), 
        .CLK(n1735), .Q(\mem0[23][7] ), .QN(n25409) );
  SDFFX1 \mem0_reg[23][6]  ( .D(n16746), .SI(\mem0[23][5] ), .SE(test_se), 
        .CLK(n1735), .Q(\mem0[23][6] ), .QN(n25410) );
  SDFFX1 \mem0_reg[23][5]  ( .D(n16745), .SI(\mem0[23][4] ), .SE(test_se), 
        .CLK(n1736), .Q(\mem0[23][5] ), .QN(n25411) );
  SDFFX1 \mem0_reg[23][4]  ( .D(n16744), .SI(\mem0[23][3] ), .SE(test_se), 
        .CLK(n1736), .Q(\mem0[23][4] ), .QN(n25412) );
  SDFFX1 \mem0_reg[23][3]  ( .D(n16743), .SI(\mem0[23][2] ), .SE(test_se), 
        .CLK(n1736), .Q(\mem0[23][3] ), .QN(n25413) );
  SDFFX1 \mem0_reg[23][2]  ( .D(n16742), .SI(\mem0[23][1] ), .SE(test_se), 
        .CLK(n1736), .Q(\mem0[23][2] ), .QN(n25414) );
  SDFFX1 \mem0_reg[23][1]  ( .D(n16741), .SI(\mem0[23][0] ), .SE(test_se), 
        .CLK(n1736), .Q(\mem0[23][1] ), .QN(n25415) );
  SDFFX1 \mem0_reg[23][0]  ( .D(n16740), .SI(\mem0[22][7] ), .SE(test_se), 
        .CLK(n1736), .Q(\mem0[23][0] ), .QN(n25416) );
  SDFFX1 \mem0_reg[22][7]  ( .D(n16739), .SI(\mem0[22][6] ), .SE(test_se), 
        .CLK(n1736), .Q(\mem0[22][7] ), .QN(n25417) );
  SDFFX1 \mem0_reg[22][6]  ( .D(n16738), .SI(\mem0[22][5] ), .SE(test_se), 
        .CLK(n1736), .Q(\mem0[22][6] ), .QN(n25418) );
  SDFFX1 \mem0_reg[22][5]  ( .D(n16737), .SI(\mem0[22][4] ), .SE(test_se), 
        .CLK(n1736), .Q(\mem0[22][5] ), .QN(n25419) );
  SDFFX1 \mem0_reg[22][4]  ( .D(n16736), .SI(\mem0[22][3] ), .SE(test_se), 
        .CLK(n1736), .Q(\mem0[22][4] ), .QN(n25420) );
  SDFFX1 \mem0_reg[22][3]  ( .D(n16735), .SI(\mem0[22][2] ), .SE(test_se), 
        .CLK(n1736), .Q(\mem0[22][3] ), .QN(n25421) );
  SDFFX1 \mem0_reg[22][2]  ( .D(n16734), .SI(\mem0[22][1] ), .SE(test_se), 
        .CLK(n1736), .Q(\mem0[22][2] ), .QN(n25422) );
  SDFFX1 \mem0_reg[22][1]  ( .D(n16733), .SI(\mem0[22][0] ), .SE(test_se), 
        .CLK(n1737), .Q(\mem0[22][1] ), .QN(n25423) );
  SDFFX1 \mem0_reg[22][0]  ( .D(n16732), .SI(test_si2), .SE(test_se), .CLK(
        n1737), .Q(\mem0[22][0] ), .QN(n25424) );
  SDFFX1 \mem0_reg[21][7]  ( .D(n16731), .SI(\mem0[21][6] ), .SE(test_se), 
        .CLK(n1393), .Q(\mem0[21][7] ), .QN(n25425) );
  SDFFX1 \mem0_reg[21][6]  ( .D(n16730), .SI(\mem0[21][5] ), .SE(test_se), 
        .CLK(n1393), .Q(\mem0[21][6] ), .QN(n25426) );
  SDFFX1 \mem0_reg[21][5]  ( .D(n16729), .SI(\mem0[21][4] ), .SE(test_se), 
        .CLK(n1393), .Q(\mem0[21][5] ), .QN(n25427) );
  SDFFX1 \mem0_reg[21][4]  ( .D(n16728), .SI(\mem0[21][3] ), .SE(test_se), 
        .CLK(n1393), .Q(\mem0[21][4] ), .QN(n25428) );
  SDFFX1 \mem0_reg[21][3]  ( .D(n16727), .SI(\mem0[21][2] ), .SE(test_se), 
        .CLK(n1393), .Q(\mem0[21][3] ), .QN(n25429) );
  SDFFX1 \mem0_reg[21][2]  ( .D(n16726), .SI(\mem0[21][1] ), .SE(test_se), 
        .CLK(n1393), .Q(\mem0[21][2] ), .QN(n25430) );
  SDFFX1 \mem0_reg[21][1]  ( .D(n16725), .SI(\mem0[21][0] ), .SE(test_se), 
        .CLK(n1393), .Q(\mem0[21][1] ), .QN(n25431) );
  SDFFX1 \mem0_reg[21][0]  ( .D(n16724), .SI(\mem0[20][7] ), .SE(test_se), 
        .CLK(n1393), .Q(\mem0[21][0] ), .QN(n25432) );
  SDFFX1 \mem0_reg[20][7]  ( .D(n16723), .SI(\mem0[20][6] ), .SE(test_se), 
        .CLK(n1393), .Q(\mem0[20][7] ), .QN(n25433) );
  SDFFX1 \mem0_reg[20][6]  ( .D(n16722), .SI(\mem0[20][5] ), .SE(test_se), 
        .CLK(n1393), .Q(\mem0[20][6] ), .QN(n25434) );
  SDFFX1 \mem0_reg[20][5]  ( .D(n16721), .SI(\mem0[20][4] ), .SE(test_se), 
        .CLK(n1393), .Q(\mem0[20][5] ), .QN(n25435) );
  SDFFX1 \mem0_reg[20][4]  ( .D(n16720), .SI(\mem0[20][3] ), .SE(test_se), 
        .CLK(n1393), .Q(\mem0[20][4] ), .QN(n25436) );
  SDFFX1 \mem0_reg[20][3]  ( .D(n16719), .SI(\mem0[20][2] ), .SE(test_se), 
        .CLK(n1394), .Q(\mem0[20][3] ), .QN(n25437) );
  SDFFX1 \mem0_reg[20][2]  ( .D(n16718), .SI(\mem0[20][1] ), .SE(test_se), 
        .CLK(n1394), .Q(\mem0[20][2] ), .QN(n25438) );
  SDFFX1 \mem0_reg[20][1]  ( .D(n16717), .SI(\mem0[20][0] ), .SE(test_se), 
        .CLK(n1394), .Q(\mem0[20][1] ), .QN(n25439) );
  SDFFX1 \mem0_reg[20][0]  ( .D(n16716), .SI(\mem0[19][7] ), .SE(test_se), 
        .CLK(n1394), .Q(\mem0[20][0] ), .QN(n25440) );
  SDFFX1 \mem0_reg[19][7]  ( .D(n16715), .SI(\mem0[19][6] ), .SE(test_se), 
        .CLK(n1394), .Q(\mem0[19][7] ), .QN(n25441) );
  SDFFX1 \mem0_reg[19][6]  ( .D(n16714), .SI(\mem0[19][5] ), .SE(test_se), 
        .CLK(n1394), .Q(\mem0[19][6] ), .QN(n25442) );
  SDFFX1 \mem0_reg[19][5]  ( .D(n16713), .SI(\mem0[19][4] ), .SE(test_se), 
        .CLK(n1394), .Q(\mem0[19][5] ), .QN(n25443) );
  SDFFX1 \mem0_reg[19][4]  ( .D(n16712), .SI(\mem0[19][3] ), .SE(test_se), 
        .CLK(n1394), .Q(\mem0[19][4] ), .QN(n25444) );
  SDFFX1 \mem0_reg[19][3]  ( .D(n16711), .SI(\mem0[19][2] ), .SE(test_se), 
        .CLK(n1394), .Q(\mem0[19][3] ), .QN(n25445) );
  SDFFX1 \mem0_reg[19][2]  ( .D(n16710), .SI(\mem0[19][1] ), .SE(test_se), 
        .CLK(n1394), .Q(\mem0[19][2] ), .QN(n25446) );
  SDFFX1 \mem0_reg[19][1]  ( .D(n16709), .SI(\mem0[19][0] ), .SE(test_se), 
        .CLK(n1394), .Q(\mem0[19][1] ), .QN(n25447) );
  SDFFX1 \mem0_reg[19][0]  ( .D(n16708), .SI(\mem0[18][7] ), .SE(test_se), 
        .CLK(n1394), .Q(\mem0[19][0] ), .QN(n25448) );
  SDFFX1 \mem0_reg[18][7]  ( .D(n16707), .SI(\mem0[18][6] ), .SE(test_se), 
        .CLK(n1395), .Q(\mem0[18][7] ), .QN(n25449) );
  SDFFX1 \mem0_reg[18][6]  ( .D(n16706), .SI(\mem0[18][5] ), .SE(test_se), 
        .CLK(n1395), .Q(\mem0[18][6] ), .QN(n25450) );
  SDFFX1 \mem0_reg[18][5]  ( .D(n16705), .SI(\mem0[18][4] ), .SE(test_se), 
        .CLK(n1395), .Q(\mem0[18][5] ), .QN(n25451) );
  SDFFX1 \mem0_reg[18][4]  ( .D(n16704), .SI(\mem0[18][3] ), .SE(test_se), 
        .CLK(n1395), .Q(\mem0[18][4] ), .QN(n25452) );
  SDFFX1 \mem0_reg[18][3]  ( .D(n16703), .SI(\mem0[18][2] ), .SE(test_se), 
        .CLK(n1395), .Q(\mem0[18][3] ), .QN(n25453) );
  SDFFX1 \mem0_reg[18][2]  ( .D(n16702), .SI(\mem0[18][1] ), .SE(test_se), 
        .CLK(n1395), .Q(\mem0[18][2] ), .QN(n25454) );
  SDFFX1 \mem0_reg[18][1]  ( .D(n16701), .SI(\mem0[18][0] ), .SE(test_se), 
        .CLK(n1395), .Q(\mem0[18][1] ), .QN(n25455) );
  SDFFX1 \mem0_reg[18][0]  ( .D(n16700), .SI(\mem0[17][7] ), .SE(test_se), 
        .CLK(n1395), .Q(\mem0[18][0] ), .QN(n25456) );
  SDFFX1 \mem0_reg[17][7]  ( .D(n16699), .SI(\mem0[17][6] ), .SE(test_se), 
        .CLK(n1395), .Q(\mem0[17][7] ), .QN(n25457) );
  SDFFX1 \mem0_reg[17][6]  ( .D(n16698), .SI(\mem0[17][5] ), .SE(test_se), 
        .CLK(n1395), .Q(\mem0[17][6] ), .QN(n25458) );
  SDFFX1 \mem0_reg[17][5]  ( .D(n16697), .SI(\mem0[17][4] ), .SE(test_se), 
        .CLK(n1395), .Q(\mem0[17][5] ), .QN(n25459) );
  SDFFX1 \mem0_reg[17][4]  ( .D(n16696), .SI(\mem0[17][3] ), .SE(test_se), 
        .CLK(n1395), .Q(\mem0[17][4] ), .QN(n25460) );
  SDFFX1 \mem0_reg[17][3]  ( .D(n16695), .SI(\mem0[17][2] ), .SE(test_se), 
        .CLK(n1396), .Q(\mem0[17][3] ), .QN(n25461) );
  SDFFX1 \mem0_reg[17][2]  ( .D(n16694), .SI(\mem0[17][1] ), .SE(test_se), 
        .CLK(n1396), .Q(\mem0[17][2] ), .QN(n25462) );
  SDFFX1 \mem0_reg[17][1]  ( .D(n16693), .SI(\mem0[17][0] ), .SE(test_se), 
        .CLK(n1396), .Q(\mem0[17][1] ), .QN(n25463) );
  SDFFX1 \mem0_reg[17][0]  ( .D(n16692), .SI(\mem0[16][7] ), .SE(test_se), 
        .CLK(n1396), .Q(\mem0[17][0] ), .QN(n25464) );
  SDFFX1 \mem0_reg[16][7]  ( .D(n16691), .SI(\mem0[16][6] ), .SE(test_se), 
        .CLK(n1396), .Q(\mem0[16][7] ), .QN(n25465) );
  SDFFX1 \mem0_reg[16][6]  ( .D(n16690), .SI(\mem0[16][5] ), .SE(test_se), 
        .CLK(n1396), .Q(\mem0[16][6] ), .QN(n25466) );
  SDFFX1 \mem0_reg[16][5]  ( .D(n16689), .SI(\mem0[16][4] ), .SE(test_se), 
        .CLK(n1396), .Q(\mem0[16][5] ), .QN(n25467) );
  SDFFX1 \mem0_reg[16][4]  ( .D(n16688), .SI(\mem0[16][3] ), .SE(test_se), 
        .CLK(n1396), .Q(\mem0[16][4] ), .QN(n25468) );
  SDFFX1 \mem0_reg[16][3]  ( .D(n16687), .SI(\mem0[16][2] ), .SE(test_se), 
        .CLK(n1396), .Q(\mem0[16][3] ), .QN(n25469) );
  SDFFX1 \mem0_reg[16][2]  ( .D(n16686), .SI(\mem0[16][1] ), .SE(test_se), 
        .CLK(n1396), .Q(\mem0[16][2] ), .QN(n25470) );
  SDFFX1 \mem0_reg[16][1]  ( .D(n16685), .SI(\mem0[16][0] ), .SE(test_se), 
        .CLK(n1396), .Q(\mem0[16][1] ), .QN(n25471) );
  SDFFX1 \mem0_reg[16][0]  ( .D(n16684), .SI(\mem0[15][7] ), .SE(test_se), 
        .CLK(n1396), .Q(\mem0[16][0] ), .QN(n25472) );
  SDFFX1 \mem0_reg[15][7]  ( .D(n16683), .SI(\mem0[15][6] ), .SE(test_se), 
        .CLK(n1397), .Q(\mem0[15][7] ), .QN(n25473) );
  SDFFX1 \mem0_reg[15][6]  ( .D(n16682), .SI(\mem0[15][5] ), .SE(test_se), 
        .CLK(n1397), .Q(\mem0[15][6] ), .QN(n25474) );
  SDFFX1 \mem0_reg[15][5]  ( .D(n16681), .SI(\mem0[15][4] ), .SE(test_se), 
        .CLK(n1397), .Q(\mem0[15][5] ), .QN(n25475) );
  SDFFX1 \mem0_reg[15][4]  ( .D(n16680), .SI(\mem0[15][3] ), .SE(test_se), 
        .CLK(n1397), .Q(\mem0[15][4] ), .QN(n25476) );
  SDFFX1 \mem0_reg[15][3]  ( .D(n16679), .SI(\mem0[15][2] ), .SE(test_se), 
        .CLK(n1397), .Q(\mem0[15][3] ), .QN(n25477) );
  SDFFX1 \mem0_reg[15][2]  ( .D(n16678), .SI(\mem0[15][1] ), .SE(test_se), 
        .CLK(n1397), .Q(\mem0[15][2] ), .QN(n25478) );
  SDFFX1 \mem0_reg[15][1]  ( .D(n16677), .SI(\mem0[15][0] ), .SE(test_se), 
        .CLK(n1397), .Q(\mem0[15][1] ), .QN(n25479) );
  SDFFX1 \mem0_reg[15][0]  ( .D(n16676), .SI(\mem0[14][7] ), .SE(test_se), 
        .CLK(n1397), .Q(\mem0[15][0] ), .QN(n25480) );
  SDFFX1 \mem0_reg[14][7]  ( .D(n16675), .SI(\mem0[14][6] ), .SE(test_se), 
        .CLK(n1397), .Q(\mem0[14][7] ), .QN(n25481) );
  SDFFX1 \mem0_reg[14][6]  ( .D(n16674), .SI(\mem0[14][5] ), .SE(test_se), 
        .CLK(n1397), .Q(\mem0[14][6] ), .QN(n25482) );
  SDFFX1 \mem0_reg[14][5]  ( .D(n16673), .SI(\mem0[14][4] ), .SE(test_se), 
        .CLK(n1397), .Q(\mem0[14][5] ), .QN(n25483) );
  SDFFX1 \mem0_reg[14][4]  ( .D(n16672), .SI(\mem0[14][3] ), .SE(test_se), 
        .CLK(n1397), .Q(\mem0[14][4] ), .QN(n25484) );
  SDFFX1 \mem0_reg[14][3]  ( .D(n16671), .SI(\mem0[14][2] ), .SE(test_se), 
        .CLK(n1398), .Q(\mem0[14][3] ), .QN(n25485) );
  SDFFX1 \mem0_reg[14][2]  ( .D(n16670), .SI(\mem0[14][1] ), .SE(test_se), 
        .CLK(n1398), .Q(\mem0[14][2] ), .QN(n25486) );
  SDFFX1 \mem0_reg[14][1]  ( .D(n16669), .SI(\mem0[14][0] ), .SE(test_se), 
        .CLK(n1398), .Q(\mem0[14][1] ), .QN(n25487) );
  SDFFX1 \mem0_reg[14][0]  ( .D(n16668), .SI(\mem0[13][7] ), .SE(test_se), 
        .CLK(n1398), .Q(\mem0[14][0] ), .QN(n25488) );
  SDFFX1 \mem0_reg[13][7]  ( .D(n16667), .SI(\mem0[13][6] ), .SE(test_se), 
        .CLK(n1398), .Q(\mem0[13][7] ), .QN(n25489) );
  SDFFX1 \mem0_reg[13][6]  ( .D(n16666), .SI(\mem0[13][5] ), .SE(test_se), 
        .CLK(n1398), .Q(\mem0[13][6] ), .QN(n25490) );
  SDFFX1 \mem0_reg[13][5]  ( .D(n16665), .SI(\mem0[13][4] ), .SE(test_se), 
        .CLK(n1398), .Q(\mem0[13][5] ), .QN(n25491) );
  SDFFX1 \mem0_reg[13][4]  ( .D(n16664), .SI(\mem0[13][3] ), .SE(test_se), 
        .CLK(n1398), .Q(\mem0[13][4] ), .QN(n25492) );
  SDFFX1 \mem0_reg[13][3]  ( .D(n16663), .SI(\mem0[13][2] ), .SE(test_se), 
        .CLK(n1398), .Q(\mem0[13][3] ), .QN(n25493) );
  SDFFX1 \mem0_reg[13][2]  ( .D(n16662), .SI(\mem0[13][1] ), .SE(test_se), 
        .CLK(n1398), .Q(\mem0[13][2] ), .QN(n25494) );
  SDFFX1 \mem0_reg[13][1]  ( .D(n16661), .SI(\mem0[13][0] ), .SE(test_se), 
        .CLK(n1398), .Q(\mem0[13][1] ), .QN(n25495) );
  SDFFX1 \mem0_reg[13][0]  ( .D(n16660), .SI(\mem0[12][7] ), .SE(test_se), 
        .CLK(n1398), .Q(\mem0[13][0] ), .QN(n25496) );
  SDFFX1 \mem0_reg[12][7]  ( .D(n16659), .SI(\mem0[12][6] ), .SE(test_se), 
        .CLK(n1399), .Q(\mem0[12][7] ), .QN(n25497) );
  SDFFX1 \mem0_reg[12][6]  ( .D(n16658), .SI(\mem0[12][5] ), .SE(test_se), 
        .CLK(n1399), .Q(\mem0[12][6] ), .QN(n25498) );
  SDFFX1 \mem0_reg[12][5]  ( .D(n16657), .SI(\mem0[12][4] ), .SE(test_se), 
        .CLK(n1399), .Q(\mem0[12][5] ), .QN(n25499) );
  SDFFX1 \mem0_reg[12][4]  ( .D(n16656), .SI(\mem0[12][3] ), .SE(test_se), 
        .CLK(n1399), .Q(\mem0[12][4] ), .QN(n25500) );
  SDFFX1 \mem0_reg[12][3]  ( .D(n16655), .SI(\mem0[12][2] ), .SE(test_se), 
        .CLK(n1399), .Q(\mem0[12][3] ), .QN(n25501) );
  SDFFX1 \mem0_reg[12][2]  ( .D(n16654), .SI(\mem0[12][1] ), .SE(test_se), 
        .CLK(n1399), .Q(\mem0[12][2] ), .QN(n25502) );
  SDFFX1 \mem0_reg[12][1]  ( .D(n16653), .SI(\mem0[12][0] ), .SE(test_se), 
        .CLK(n1399), .Q(\mem0[12][1] ), .QN(n25503) );
  SDFFX1 \mem0_reg[12][0]  ( .D(n16652), .SI(\mem0[11][7] ), .SE(test_se), 
        .CLK(n1399), .Q(\mem0[12][0] ), .QN(n25504) );
  SDFFX1 \mem0_reg[11][7]  ( .D(n16651), .SI(\mem0[11][6] ), .SE(test_se), 
        .CLK(n1399), .Q(\mem0[11][7] ), .QN(n25505) );
  SDFFX1 \mem0_reg[11][6]  ( .D(n16650), .SI(\mem0[11][5] ), .SE(test_se), 
        .CLK(n1399), .Q(\mem0[11][6] ), .QN(n25506) );
  SDFFX1 \mem0_reg[11][5]  ( .D(n16649), .SI(\mem0[11][4] ), .SE(test_se), 
        .CLK(n1399), .Q(\mem0[11][5] ), .QN(n25507) );
  SDFFX1 \mem0_reg[11][4]  ( .D(n16648), .SI(\mem0[11][3] ), .SE(test_se), 
        .CLK(n1399), .Q(\mem0[11][4] ), .QN(n25508) );
  SDFFX1 \mem0_reg[11][3]  ( .D(n16647), .SI(\mem0[11][2] ), .SE(test_se), 
        .CLK(n1400), .Q(\mem0[11][3] ), .QN(n25509) );
  SDFFX1 \mem0_reg[11][2]  ( .D(n16646), .SI(\mem0[11][1] ), .SE(test_se), 
        .CLK(n1400), .Q(\mem0[11][2] ), .QN(n25510) );
  SDFFX1 \mem0_reg[11][1]  ( .D(n16645), .SI(\mem0[11][0] ), .SE(test_se), 
        .CLK(n1400), .Q(\mem0[11][1] ), .QN(n25511) );
  SDFFX1 \mem0_reg[11][0]  ( .D(n16644), .SI(\mem0[10][7] ), .SE(test_se), 
        .CLK(n1400), .Q(\mem0[11][0] ), .QN(n25512) );
  SDFFX1 \mem0_reg[10][7]  ( .D(n16643), .SI(\mem0[10][6] ), .SE(test_se), 
        .CLK(n1400), .Q(\mem0[10][7] ), .QN(n25513) );
  SDFFX1 \mem0_reg[10][6]  ( .D(n16642), .SI(\mem0[10][5] ), .SE(test_se), 
        .CLK(n1400), .Q(\mem0[10][6] ), .QN(n25514) );
  SDFFX1 \mem0_reg[10][5]  ( .D(n16641), .SI(\mem0[10][4] ), .SE(test_se), 
        .CLK(n1400), .Q(\mem0[10][5] ), .QN(n25515) );
  SDFFX1 \mem0_reg[10][4]  ( .D(n16640), .SI(\mem0[10][3] ), .SE(test_se), 
        .CLK(n1400), .Q(\mem0[10][4] ), .QN(n25516) );
  SDFFX1 \mem0_reg[10][3]  ( .D(n16639), .SI(\mem0[10][2] ), .SE(test_se), 
        .CLK(n1400), .Q(\mem0[10][3] ), .QN(n25517) );
  SDFFX1 \mem0_reg[10][2]  ( .D(n16638), .SI(\mem0[10][1] ), .SE(test_se), 
        .CLK(n1400), .Q(\mem0[10][2] ), .QN(n25518) );
  SDFFX1 \mem0_reg[10][1]  ( .D(n16637), .SI(\mem0[10][0] ), .SE(test_se), 
        .CLK(n1400), .Q(\mem0[10][1] ), .QN(n25519) );
  SDFFX1 \mem0_reg[10][0]  ( .D(n16636), .SI(\mem0[9][7] ), .SE(test_se), 
        .CLK(n1400), .Q(\mem0[10][0] ), .QN(n25520) );
  SDFFX1 \mem0_reg[9][7]  ( .D(n16635), .SI(\mem0[9][6] ), .SE(test_se), .CLK(
        n1401), .Q(\mem0[9][7] ), .QN(n25521) );
  SDFFX1 \mem0_reg[9][6]  ( .D(n16634), .SI(\mem0[9][5] ), .SE(test_se), .CLK(
        n1401), .Q(\mem0[9][6] ), .QN(n25522) );
  SDFFX1 \mem0_reg[9][5]  ( .D(n16633), .SI(\mem0[9][4] ), .SE(test_se), .CLK(
        n1401), .Q(\mem0[9][5] ), .QN(n25523) );
  SDFFX1 \mem0_reg[9][4]  ( .D(n16632), .SI(\mem0[9][3] ), .SE(test_se), .CLK(
        n1401), .Q(\mem0[9][4] ), .QN(n25524) );
  SDFFX1 \mem0_reg[9][3]  ( .D(n16631), .SI(\mem0[9][2] ), .SE(test_se), .CLK(
        n1401), .Q(\mem0[9][3] ), .QN(n25525) );
  SDFFX1 \mem0_reg[9][2]  ( .D(n16630), .SI(\mem0[9][1] ), .SE(test_se), .CLK(
        n1401), .Q(\mem0[9][2] ), .QN(n25526) );
  SDFFX1 \mem0_reg[9][1]  ( .D(n16629), .SI(\mem0[9][0] ), .SE(test_se), .CLK(
        n1401), .Q(\mem0[9][1] ), .QN(n25527) );
  SDFFX1 \mem0_reg[9][0]  ( .D(n16628), .SI(\mem0[8][7] ), .SE(test_se), .CLK(
        n1401), .Q(\mem0[9][0] ), .QN(n25528) );
  SDFFX1 \mem0_reg[8][7]  ( .D(n16627), .SI(\mem0[8][6] ), .SE(test_se), .CLK(
        n1401), .Q(\mem0[8][7] ), .QN(n25529) );
  SDFFX1 \mem0_reg[8][6]  ( .D(n16626), .SI(\mem0[8][5] ), .SE(test_se), .CLK(
        n1401), .Q(\mem0[8][6] ), .QN(n25530) );
  SDFFX1 \mem0_reg[8][5]  ( .D(n16625), .SI(\mem0[8][4] ), .SE(test_se), .CLK(
        n1401), .Q(\mem0[8][5] ), .QN(n25531) );
  SDFFX1 \mem0_reg[8][4]  ( .D(n16624), .SI(\mem0[8][3] ), .SE(test_se), .CLK(
        n1401), .Q(\mem0[8][4] ), .QN(n25532) );
  SDFFX1 \mem0_reg[8][3]  ( .D(n16623), .SI(\mem0[8][2] ), .SE(test_se), .CLK(
        n1402), .Q(\mem0[8][3] ), .QN(n25533) );
  SDFFX1 \mem0_reg[8][2]  ( .D(n16622), .SI(\mem0[8][1] ), .SE(test_se), .CLK(
        n1402), .Q(\mem0[8][2] ), .QN(n25534) );
  SDFFX1 \mem0_reg[8][1]  ( .D(n16621), .SI(\mem0[8][0] ), .SE(test_se), .CLK(
        n1402), .Q(\mem0[8][1] ), .QN(n25535) );
  SDFFX1 \mem0_reg[8][0]  ( .D(n16620), .SI(\mem0[7][7] ), .SE(test_se), .CLK(
        n1402), .Q(\mem0[8][0] ), .QN(n25536) );
  SDFFX1 \mem0_reg[7][7]  ( .D(n16619), .SI(\mem0[7][6] ), .SE(test_se), .CLK(
        n1402), .Q(\mem0[7][7] ), .QN(n25537) );
  SDFFX1 \mem0_reg[7][6]  ( .D(n16618), .SI(\mem0[7][5] ), .SE(test_se), .CLK(
        n1402), .Q(\mem0[7][6] ), .QN(n25538) );
  SDFFX1 \mem0_reg[7][5]  ( .D(n16617), .SI(\mem0[7][4] ), .SE(test_se), .CLK(
        n1402), .Q(\mem0[7][5] ), .QN(n25539) );
  SDFFX1 \mem0_reg[7][4]  ( .D(n16616), .SI(\mem0[7][3] ), .SE(test_se), .CLK(
        n1402), .Q(\mem0[7][4] ), .QN(n25540) );
  SDFFX1 \mem0_reg[7][3]  ( .D(n16615), .SI(\mem0[7][2] ), .SE(test_se), .CLK(
        n1402), .Q(\mem0[7][3] ), .QN(n25541) );
  SDFFX1 \mem0_reg[7][2]  ( .D(n16614), .SI(\mem0[7][1] ), .SE(test_se), .CLK(
        n1402), .Q(\mem0[7][2] ), .QN(n25542) );
  SDFFX1 \mem0_reg[7][1]  ( .D(n16613), .SI(\mem0[7][0] ), .SE(test_se), .CLK(
        n1402), .Q(\mem0[7][1] ), .QN(n25543) );
  SDFFX1 \mem0_reg[7][0]  ( .D(n16612), .SI(\mem0[6][7] ), .SE(test_se), .CLK(
        n1402), .Q(\mem0[7][0] ), .QN(n25544) );
  SDFFX1 \mem0_reg[6][7]  ( .D(n16611), .SI(\mem0[6][6] ), .SE(test_se), .CLK(
        n1403), .Q(\mem0[6][7] ), .QN(n25545) );
  SDFFX1 \mem0_reg[6][6]  ( .D(n16610), .SI(\mem0[6][5] ), .SE(test_se), .CLK(
        n1403), .Q(\mem0[6][6] ), .QN(n25546) );
  SDFFX1 \mem0_reg[6][5]  ( .D(n16609), .SI(\mem0[6][4] ), .SE(test_se), .CLK(
        n1403), .Q(\mem0[6][5] ), .QN(n25547) );
  SDFFX1 \mem0_reg[6][4]  ( .D(n16608), .SI(\mem0[6][3] ), .SE(test_se), .CLK(
        n1403), .Q(\mem0[6][4] ), .QN(n25548) );
  SDFFX1 \mem0_reg[6][3]  ( .D(n16607), .SI(\mem0[6][2] ), .SE(test_se), .CLK(
        n1403), .Q(\mem0[6][3] ), .QN(n25549) );
  SDFFX1 \mem0_reg[6][2]  ( .D(n16606), .SI(\mem0[6][1] ), .SE(test_se), .CLK(
        n1403), .Q(\mem0[6][2] ), .QN(n25550) );
  SDFFX1 \mem0_reg[6][1]  ( .D(n16605), .SI(\mem0[6][0] ), .SE(test_se), .CLK(
        n1403), .Q(\mem0[6][1] ), .QN(n25551) );
  SDFFX1 \mem0_reg[6][0]  ( .D(n16604), .SI(\mem0[5][7] ), .SE(test_se), .CLK(
        n1403), .Q(\mem0[6][0] ), .QN(n25552) );
  SDFFX1 \mem0_reg[5][7]  ( .D(n16603), .SI(\mem0[5][6] ), .SE(test_se), .CLK(
        n1403), .Q(\mem0[5][7] ), .QN(n25553) );
  SDFFX1 \mem0_reg[5][6]  ( .D(n16602), .SI(\mem0[5][5] ), .SE(test_se), .CLK(
        n1403), .Q(\mem0[5][6] ), .QN(n25554) );
  SDFFX1 \mem0_reg[5][5]  ( .D(n16601), .SI(\mem0[5][4] ), .SE(test_se), .CLK(
        n1403), .Q(\mem0[5][5] ), .QN(n25555) );
  SDFFX1 \mem0_reg[5][4]  ( .D(n16600), .SI(\mem0[5][3] ), .SE(test_se), .CLK(
        n1403), .Q(\mem0[5][4] ), .QN(n25556) );
  SDFFX1 \mem0_reg[5][3]  ( .D(n16599), .SI(\mem0[5][2] ), .SE(test_se), .CLK(
        n1404), .Q(\mem0[5][3] ), .QN(n25557) );
  SDFFX1 \mem0_reg[5][2]  ( .D(n16598), .SI(\mem0[5][1] ), .SE(test_se), .CLK(
        n1404), .Q(\mem0[5][2] ), .QN(n25558) );
  SDFFX1 \mem0_reg[5][1]  ( .D(n16597), .SI(\mem0[5][0] ), .SE(test_se), .CLK(
        n1404), .Q(\mem0[5][1] ), .QN(n25559) );
  SDFFX1 \mem0_reg[5][0]  ( .D(n16596), .SI(\mem0[4][7] ), .SE(test_se), .CLK(
        n1404), .Q(\mem0[5][0] ), .QN(n25560) );
  SDFFX1 \mem0_reg[4][7]  ( .D(n16595), .SI(\mem0[4][6] ), .SE(test_se), .CLK(
        n1404), .Q(\mem0[4][7] ), .QN(n25561) );
  SDFFX1 \mem0_reg[4][6]  ( .D(n16594), .SI(\mem0[4][5] ), .SE(test_se), .CLK(
        n1404), .Q(\mem0[4][6] ), .QN(n25562) );
  SDFFX1 \mem0_reg[4][5]  ( .D(n16593), .SI(\mem0[4][4] ), .SE(test_se), .CLK(
        n1404), .Q(\mem0[4][5] ), .QN(n25563) );
  SDFFX1 \mem0_reg[4][4]  ( .D(n16592), .SI(\mem0[4][3] ), .SE(test_se), .CLK(
        n1404), .Q(\mem0[4][4] ), .QN(n25564) );
  SDFFX1 \mem0_reg[4][3]  ( .D(n16591), .SI(\mem0[4][2] ), .SE(test_se), .CLK(
        n1404), .Q(\mem0[4][3] ), .QN(n25565) );
  SDFFX1 \mem0_reg[4][2]  ( .D(n16590), .SI(\mem0[4][1] ), .SE(test_se), .CLK(
        n1404), .Q(\mem0[4][2] ), .QN(n25566) );
  SDFFX1 \mem0_reg[4][1]  ( .D(n16589), .SI(\mem0[4][0] ), .SE(test_se), .CLK(
        n1404), .Q(\mem0[4][1] ), .QN(n25567) );
  SDFFX1 \mem0_reg[4][0]  ( .D(n16588), .SI(\mem0[3][7] ), .SE(test_se), .CLK(
        n1404), .Q(\mem0[4][0] ), .QN(n25568) );
  SDFFX1 \mem0_reg[3][7]  ( .D(n16587), .SI(\mem0[3][6] ), .SE(test_se), .CLK(
        n1405), .Q(\mem0[3][7] ), .QN(n25569) );
  SDFFX1 \mem0_reg[3][6]  ( .D(n16586), .SI(\mem0[3][5] ), .SE(test_se), .CLK(
        n1405), .Q(\mem0[3][6] ), .QN(n25570) );
  SDFFX1 \mem0_reg[3][5]  ( .D(n16585), .SI(\mem0[3][4] ), .SE(test_se), .CLK(
        n1405), .Q(\mem0[3][5] ), .QN(n25571) );
  SDFFX1 \mem0_reg[3][4]  ( .D(n16584), .SI(\mem0[3][3] ), .SE(test_se), .CLK(
        n1405), .Q(\mem0[3][4] ), .QN(n25572) );
  SDFFX1 \mem0_reg[3][3]  ( .D(n16583), .SI(\mem0[3][2] ), .SE(test_se), .CLK(
        n1405), .Q(\mem0[3][3] ), .QN(n25573) );
  SDFFX1 \mem0_reg[3][2]  ( .D(n16582), .SI(\mem0[3][1] ), .SE(test_se), .CLK(
        n1405), .Q(\mem0[3][2] ), .QN(n25574) );
  SDFFX1 \mem0_reg[3][1]  ( .D(n16581), .SI(\mem0[3][0] ), .SE(test_se), .CLK(
        n1405), .Q(\mem0[3][1] ), .QN(n25575) );
  SDFFX1 \mem0_reg[3][0]  ( .D(n16580), .SI(\mem0[2][7] ), .SE(test_se), .CLK(
        n1405), .Q(\mem0[3][0] ), .QN(n25576) );
  SDFFX1 \mem0_reg[2][7]  ( .D(n16579), .SI(\mem0[2][6] ), .SE(test_se), .CLK(
        n1405), .Q(\mem0[2][7] ), .QN(n25577) );
  SDFFX1 \mem0_reg[2][6]  ( .D(n16578), .SI(\mem0[2][5] ), .SE(test_se), .CLK(
        n1405), .Q(\mem0[2][6] ), .QN(n25578) );
  SDFFX1 \mem0_reg[2][5]  ( .D(n16577), .SI(\mem0[2][4] ), .SE(test_se), .CLK(
        n1405), .Q(\mem0[2][5] ), .QN(n25579) );
  SDFFX1 \mem0_reg[2][4]  ( .D(n16576), .SI(\mem0[2][3] ), .SE(test_se), .CLK(
        n1405), .Q(\mem0[2][4] ), .QN(n25580) );
  SDFFX1 \mem0_reg[2][3]  ( .D(n16575), .SI(\mem0[2][2] ), .SE(test_se), .CLK(
        n1406), .Q(\mem0[2][3] ), .QN(n25581) );
  SDFFX1 \mem0_reg[2][2]  ( .D(n16574), .SI(\mem0[2][1] ), .SE(test_se), .CLK(
        n1406), .Q(\mem0[2][2] ), .QN(n25582) );
  SDFFX1 \mem0_reg[2][1]  ( .D(n16573), .SI(\mem0[2][0] ), .SE(test_se), .CLK(
        n1406), .Q(\mem0[2][1] ), .QN(n25583) );
  SDFFX1 \mem0_reg[2][0]  ( .D(n16572), .SI(\mem0[1][7] ), .SE(test_se), .CLK(
        n1406), .Q(\mem0[2][0] ), .QN(n25584) );
  SDFFX1 \mem0_reg[1][7]  ( .D(n16571), .SI(\mem0[1][6] ), .SE(test_se), .CLK(
        n1406), .Q(\mem0[1][7] ), .QN(n25585) );
  SDFFX1 \mem0_reg[1][6]  ( .D(n16570), .SI(\mem0[1][5] ), .SE(test_se), .CLK(
        n1406), .Q(\mem0[1][6] ), .QN(n25586) );
  SDFFX1 \mem0_reg[1][5]  ( .D(n16569), .SI(\mem0[1][4] ), .SE(test_se), .CLK(
        n1406), .Q(\mem0[1][5] ), .QN(n25587) );
  SDFFX1 \mem0_reg[1][4]  ( .D(n16568), .SI(\mem0[1][3] ), .SE(test_se), .CLK(
        n1406), .Q(\mem0[1][4] ), .QN(n25588) );
  SDFFX1 \mem0_reg[1][3]  ( .D(n16567), .SI(\mem0[1][2] ), .SE(test_se), .CLK(
        n1406), .Q(\mem0[1][3] ), .QN(n25589) );
  SDFFX1 \mem0_reg[1][2]  ( .D(n16566), .SI(\mem0[1][1] ), .SE(test_se), .CLK(
        n1406), .Q(\mem0[1][2] ), .QN(n25590) );
  SDFFX1 \mem0_reg[1][1]  ( .D(n16565), .SI(\mem0[1][0] ), .SE(test_se), .CLK(
        n1406), .Q(\mem0[1][1] ), .QN(n25591) );
  SDFFX1 \mem0_reg[1][0]  ( .D(n16564), .SI(\mem0[0][7] ), .SE(test_se), .CLK(
        n1406), .Q(\mem0[1][0] ), .QN(n25592) );
  SDFFX1 \mem0_reg[0][7]  ( .D(n16563), .SI(\mem0[0][6] ), .SE(test_se), .CLK(
        n1407), .Q(\mem0[0][7] ), .QN(n25593) );
  SDFFX1 \mem0_reg[0][6]  ( .D(n16562), .SI(\mem0[0][5] ), .SE(test_se), .CLK(
        n1407), .Q(\mem0[0][6] ), .QN(n25594) );
  SDFFX1 \mem0_reg[0][5]  ( .D(n16561), .SI(\mem0[0][4] ), .SE(test_se), .CLK(
        n1407), .Q(\mem0[0][5] ), .QN(n25595) );
  SDFFX1 \mem0_reg[0][4]  ( .D(n16560), .SI(\mem0[0][3] ), .SE(test_se), .CLK(
        n1407), .Q(\mem0[0][4] ), .QN(n25596) );
  SDFFX1 \mem0_reg[0][3]  ( .D(n16559), .SI(\mem0[0][2] ), .SE(test_se), .CLK(
        n1407), .Q(\mem0[0][3] ), .QN(n25597) );
  SDFFX1 \mem0_reg[0][2]  ( .D(n16558), .SI(\mem0[0][1] ), .SE(test_se), .CLK(
        n1407), .Q(\mem0[0][2] ), .QN(n25598) );
  SDFFX1 \mem0_reg[0][1]  ( .D(n16557), .SI(\mem0[0][0] ), .SE(test_se), .CLK(
        n1407), .Q(\mem0[0][1] ), .QN(n25599) );
  SDFFX1 \mem0_reg[0][0]  ( .D(n16556), .SI(test_si1), .SE(test_se), .CLK(
        n1407), .Q(\mem0[0][0] ), .QN(n25600) );
  SDFFX1 \mem1_reg[255][15]  ( .D(n16555), .SI(\mem1[255][14] ), .SE(test_se), 
        .CLK(n1410), .Q(\mem1[255][15] ), .QN(n25601) );
  SDFFX1 \mem1_reg[255][14]  ( .D(n16554), .SI(\mem1[255][13] ), .SE(test_se), 
        .CLK(n1410), .Q(\mem1[255][14] ), .QN(n25602) );
  SDFFX1 \mem1_reg[255][13]  ( .D(n16553), .SI(\mem1[255][12] ), .SE(test_se), 
        .CLK(n1410), .Q(\mem1[255][13] ), .QN(n25603) );
  SDFFX1 \mem1_reg[255][12]  ( .D(n16552), .SI(\mem1[255][11] ), .SE(test_se), 
        .CLK(n1410), .Q(\mem1[255][12] ), .QN(n25604) );
  SDFFX1 \mem1_reg[255][11]  ( .D(n16551), .SI(\mem1[255][10] ), .SE(test_se), 
        .CLK(n1410), .Q(\mem1[255][11] ), .QN(n25605) );
  SDFFX1 \mem1_reg[255][10]  ( .D(n16550), .SI(\mem1[255][9] ), .SE(test_se), 
        .CLK(n1410), .Q(\mem1[255][10] ), .QN(n25606) );
  SDFFX1 \mem1_reg[255][9]  ( .D(n16549), .SI(\mem1[255][8] ), .SE(test_se), 
        .CLK(n1411), .Q(\mem1[255][9] ), .QN(n25607) );
  SDFFX1 \mem1_reg[255][8]  ( .D(n16548), .SI(\mem1[254][15] ), .SE(test_se), 
        .CLK(n1411), .Q(\mem1[255][8] ), .QN(n25608) );
  SDFFX1 \mem1_reg[254][15]  ( .D(n16547), .SI(\mem1[254][14] ), .SE(test_se), 
        .CLK(n1411), .Q(\mem1[254][15] ), .QN(n25609) );
  SDFFX1 \mem1_reg[254][14]  ( .D(n16546), .SI(\mem1[254][13] ), .SE(test_se), 
        .CLK(n1411), .Q(\mem1[254][14] ), .QN(n25610) );
  SDFFX1 \mem1_reg[254][13]  ( .D(n16545), .SI(\mem1[254][12] ), .SE(test_se), 
        .CLK(n1411), .Q(\mem1[254][13] ), .QN(n25611) );
  SDFFX1 \mem1_reg[254][12]  ( .D(n16544), .SI(\mem1[254][11] ), .SE(test_se), 
        .CLK(n1411), .Q(\mem1[254][12] ), .QN(n25612) );
  SDFFX1 \mem1_reg[254][11]  ( .D(n16543), .SI(\mem1[254][10] ), .SE(test_se), 
        .CLK(n1411), .Q(\mem1[254][11] ), .QN(n25613) );
  SDFFX1 \mem1_reg[254][10]  ( .D(n16542), .SI(\mem1[254][9] ), .SE(test_se), 
        .CLK(n1411), .Q(\mem1[254][10] ), .QN(n25614) );
  SDFFX1 \mem1_reg[254][9]  ( .D(n16541), .SI(\mem1[254][8] ), .SE(test_se), 
        .CLK(n1411), .Q(\mem1[254][9] ), .QN(n25615) );
  SDFFX1 \mem1_reg[254][8]  ( .D(n16540), .SI(\mem1[253][15] ), .SE(test_se), 
        .CLK(n1411), .Q(\mem1[254][8] ), .QN(n25616) );
  SDFFX1 \mem1_reg[253][15]  ( .D(n16539), .SI(\mem1[253][14] ), .SE(test_se), 
        .CLK(n1411), .Q(\mem1[253][15] ), .QN(n25617) );
  SDFFX1 \mem1_reg[253][14]  ( .D(n16538), .SI(\mem1[253][13] ), .SE(test_se), 
        .CLK(n1411), .Q(\mem1[253][14] ), .QN(n25618) );
  SDFFX1 \mem1_reg[253][13]  ( .D(n16537), .SI(\mem1[253][12] ), .SE(test_se), 
        .CLK(n1412), .Q(\mem1[253][13] ), .QN(n25619) );
  SDFFX1 \mem1_reg[253][12]  ( .D(n16536), .SI(\mem1[253][11] ), .SE(test_se), 
        .CLK(n1412), .Q(\mem1[253][12] ), .QN(n25620) );
  SDFFX1 \mem1_reg[253][11]  ( .D(n16535), .SI(\mem1[253][10] ), .SE(test_se), 
        .CLK(n1412), .Q(\mem1[253][11] ), .QN(n25621) );
  SDFFX1 \mem1_reg[253][10]  ( .D(n16534), .SI(\mem1[253][9] ), .SE(test_se), 
        .CLK(n1412), .Q(\mem1[253][10] ), .QN(n25622) );
  SDFFX1 \mem1_reg[253][9]  ( .D(n16533), .SI(\mem1[253][8] ), .SE(test_se), 
        .CLK(n1412), .Q(\mem1[253][9] ), .QN(n25623) );
  SDFFX1 \mem1_reg[253][8]  ( .D(n16532), .SI(\mem1[252][15] ), .SE(test_se), 
        .CLK(n1412), .Q(\mem1[253][8] ), .QN(n25624) );
  SDFFX1 \mem1_reg[252][15]  ( .D(n16531), .SI(\mem1[252][14] ), .SE(test_se), 
        .CLK(n1412), .Q(\mem1[252][15] ), .QN(n25625) );
  SDFFX1 \mem1_reg[252][14]  ( .D(n16530), .SI(\mem1[252][13] ), .SE(test_se), 
        .CLK(n1412), .Q(\mem1[252][14] ), .QN(n25626) );
  SDFFX1 \mem1_reg[252][13]  ( .D(n16529), .SI(\mem1[252][12] ), .SE(test_se), 
        .CLK(n1412), .Q(\mem1[252][13] ), .QN(n25627) );
  SDFFX1 \mem1_reg[252][12]  ( .D(n16528), .SI(\mem1[252][11] ), .SE(test_se), 
        .CLK(n1412), .Q(\mem1[252][12] ), .QN(n25628) );
  SDFFX1 \mem1_reg[252][11]  ( .D(n16527), .SI(\mem1[252][10] ), .SE(test_se), 
        .CLK(n1412), .Q(\mem1[252][11] ), .QN(n25629) );
  SDFFX1 \mem1_reg[252][10]  ( .D(n16526), .SI(\mem1[252][9] ), .SE(test_se), 
        .CLK(n1412), .Q(\mem1[252][10] ), .QN(n25630) );
  SDFFX1 \mem1_reg[252][9]  ( .D(n16525), .SI(\mem1[252][8] ), .SE(test_se), 
        .CLK(n1413), .Q(\mem1[252][9] ), .QN(n25631) );
  SDFFX1 \mem1_reg[252][8]  ( .D(n16524), .SI(\mem1[251][15] ), .SE(test_se), 
        .CLK(n1413), .Q(\mem1[252][8] ), .QN(n25632) );
  SDFFX1 \mem1_reg[251][15]  ( .D(n16523), .SI(\mem1[251][14] ), .SE(test_se), 
        .CLK(n1413), .Q(\mem1[251][15] ), .QN(n25633) );
  SDFFX1 \mem1_reg[251][14]  ( .D(n16522), .SI(\mem1[251][13] ), .SE(test_se), 
        .CLK(n1413), .Q(\mem1[251][14] ), .QN(n25634) );
  SDFFX1 \mem1_reg[251][13]  ( .D(n16521), .SI(\mem1[251][12] ), .SE(test_se), 
        .CLK(n1413), .Q(\mem1[251][13] ), .QN(n25635) );
  SDFFX1 \mem1_reg[251][12]  ( .D(n16520), .SI(\mem1[251][11] ), .SE(test_se), 
        .CLK(n1413), .Q(\mem1[251][12] ), .QN(n25636) );
  SDFFX1 \mem1_reg[251][11]  ( .D(n16519), .SI(\mem1[251][10] ), .SE(test_se), 
        .CLK(n1413), .Q(\mem1[251][11] ), .QN(n25637) );
  SDFFX1 \mem1_reg[251][10]  ( .D(n16518), .SI(\mem1[251][9] ), .SE(test_se), 
        .CLK(n1413), .Q(\mem1[251][10] ), .QN(n25638) );
  SDFFX1 \mem1_reg[251][9]  ( .D(n16517), .SI(\mem1[251][8] ), .SE(test_se), 
        .CLK(n1413), .Q(\mem1[251][9] ), .QN(n25639) );
  SDFFX1 \mem1_reg[251][8]  ( .D(n16516), .SI(\mem1[250][15] ), .SE(test_se), 
        .CLK(n1413), .Q(\mem1[251][8] ), .QN(n25640) );
  SDFFX1 \mem1_reg[250][15]  ( .D(n16515), .SI(\mem1[250][14] ), .SE(test_se), 
        .CLK(n1413), .Q(\mem1[250][15] ), .QN(n25641) );
  SDFFX1 \mem1_reg[250][14]  ( .D(n16514), .SI(\mem1[250][13] ), .SE(test_se), 
        .CLK(n1413), .Q(\mem1[250][14] ), .QN(n25642) );
  SDFFX1 \mem1_reg[250][13]  ( .D(n16513), .SI(\mem1[250][12] ), .SE(test_se), 
        .CLK(n1414), .Q(\mem1[250][13] ), .QN(n25643) );
  SDFFX1 \mem1_reg[250][12]  ( .D(n16512), .SI(\mem1[250][11] ), .SE(test_se), 
        .CLK(n1414), .Q(\mem1[250][12] ), .QN(n25644) );
  SDFFX1 \mem1_reg[250][11]  ( .D(n16511), .SI(\mem1[250][10] ), .SE(test_se), 
        .CLK(n1414), .Q(\mem1[250][11] ), .QN(n25645) );
  SDFFX1 \mem1_reg[250][10]  ( .D(n16510), .SI(\mem1[250][9] ), .SE(test_se), 
        .CLK(n1414), .Q(\mem1[250][10] ), .QN(n25646) );
  SDFFX1 \mem1_reg[250][9]  ( .D(n16509), .SI(\mem1[250][8] ), .SE(test_se), 
        .CLK(n1414), .Q(\mem1[250][9] ), .QN(n25647) );
  SDFFX1 \mem1_reg[250][8]  ( .D(n16508), .SI(\mem1[249][15] ), .SE(test_se), 
        .CLK(n1414), .Q(\mem1[250][8] ), .QN(n25648) );
  SDFFX1 \mem1_reg[249][15]  ( .D(n16507), .SI(\mem1[249][14] ), .SE(test_se), 
        .CLK(n1414), .Q(\mem1[249][15] ), .QN(n25649) );
  SDFFX1 \mem1_reg[249][14]  ( .D(n16506), .SI(\mem1[249][13] ), .SE(test_se), 
        .CLK(n1414), .Q(\mem1[249][14] ), .QN(n25650) );
  SDFFX1 \mem1_reg[249][13]  ( .D(n16505), .SI(\mem1[249][12] ), .SE(test_se), 
        .CLK(n1414), .Q(\mem1[249][13] ), .QN(n25651) );
  SDFFX1 \mem1_reg[249][12]  ( .D(n16504), .SI(\mem1[249][11] ), .SE(test_se), 
        .CLK(n1414), .Q(\mem1[249][12] ), .QN(n25652) );
  SDFFX1 \mem1_reg[249][11]  ( .D(n16503), .SI(\mem1[249][10] ), .SE(test_se), 
        .CLK(n1414), .Q(\mem1[249][11] ), .QN(n25653) );
  SDFFX1 \mem1_reg[249][10]  ( .D(n16502), .SI(\mem1[249][9] ), .SE(test_se), 
        .CLK(n1414), .Q(\mem1[249][10] ), .QN(n25654) );
  SDFFX1 \mem1_reg[249][9]  ( .D(n16501), .SI(\mem1[249][8] ), .SE(test_se), 
        .CLK(n1415), .Q(\mem1[249][9] ), .QN(n25655) );
  SDFFX1 \mem1_reg[249][8]  ( .D(n16500), .SI(\mem1[248][15] ), .SE(test_se), 
        .CLK(n1415), .Q(\mem1[249][8] ), .QN(n25656) );
  SDFFX1 \mem1_reg[248][15]  ( .D(n16499), .SI(\mem1[248][14] ), .SE(test_se), 
        .CLK(n1415), .Q(\mem1[248][15] ), .QN(n25657) );
  SDFFX1 \mem1_reg[248][14]  ( .D(n16498), .SI(\mem1[248][13] ), .SE(test_se), 
        .CLK(n1415), .Q(\mem1[248][14] ), .QN(n25658) );
  SDFFX1 \mem1_reg[248][13]  ( .D(n16497), .SI(\mem1[248][12] ), .SE(test_se), 
        .CLK(n1415), .Q(\mem1[248][13] ), .QN(n25659) );
  SDFFX1 \mem1_reg[248][12]  ( .D(n16496), .SI(\mem1[248][11] ), .SE(test_se), 
        .CLK(n1415), .Q(\mem1[248][12] ), .QN(n25660) );
  SDFFX1 \mem1_reg[248][11]  ( .D(n16495), .SI(\mem1[248][10] ), .SE(test_se), 
        .CLK(n1415), .Q(\mem1[248][11] ), .QN(n25661) );
  SDFFX1 \mem1_reg[248][10]  ( .D(n16494), .SI(\mem1[248][9] ), .SE(test_se), 
        .CLK(n1415), .Q(\mem1[248][10] ), .QN(n25662) );
  SDFFX1 \mem1_reg[248][9]  ( .D(n16493), .SI(\mem1[248][8] ), .SE(test_se), 
        .CLK(n1415), .Q(\mem1[248][9] ), .QN(n25663) );
  SDFFX1 \mem1_reg[248][8]  ( .D(n16492), .SI(\mem1[247][15] ), .SE(test_se), 
        .CLK(n1415), .Q(\mem1[248][8] ), .QN(n25664) );
  SDFFX1 \mem1_reg[247][15]  ( .D(n16491), .SI(\mem1[247][14] ), .SE(test_se), 
        .CLK(n1415), .Q(\mem1[247][15] ), .QN(n25665) );
  SDFFX1 \mem1_reg[247][14]  ( .D(n16490), .SI(\mem1[247][13] ), .SE(test_se), 
        .CLK(n1415), .Q(\mem1[247][14] ), .QN(n25666) );
  SDFFX1 \mem1_reg[247][13]  ( .D(n16489), .SI(\mem1[247][12] ), .SE(test_se), 
        .CLK(n1416), .Q(\mem1[247][13] ), .QN(n25667) );
  SDFFX1 \mem1_reg[247][12]  ( .D(n16488), .SI(\mem1[247][11] ), .SE(test_se), 
        .CLK(n1416), .Q(\mem1[247][12] ), .QN(n25668) );
  SDFFX1 \mem1_reg[247][11]  ( .D(n16487), .SI(\mem1[247][10] ), .SE(test_se), 
        .CLK(n1416), .Q(\mem1[247][11] ), .QN(n25669) );
  SDFFX1 \mem1_reg[247][10]  ( .D(n16486), .SI(\mem1[247][9] ), .SE(test_se), 
        .CLK(n1416), .Q(\mem1[247][10] ), .QN(n25670) );
  SDFFX1 \mem1_reg[247][9]  ( .D(n16485), .SI(\mem1[247][8] ), .SE(test_se), 
        .CLK(n1416), .Q(\mem1[247][9] ), .QN(n25671) );
  SDFFX1 \mem1_reg[247][8]  ( .D(n16484), .SI(\mem1[246][15] ), .SE(test_se), 
        .CLK(n1416), .Q(\mem1[247][8] ), .QN(n25672) );
  SDFFX1 \mem1_reg[246][15]  ( .D(n16483), .SI(\mem1[246][14] ), .SE(test_se), 
        .CLK(n1416), .Q(\mem1[246][15] ), .QN(n25673) );
  SDFFX1 \mem1_reg[246][14]  ( .D(n16482), .SI(\mem1[246][13] ), .SE(test_se), 
        .CLK(n1416), .Q(\mem1[246][14] ), .QN(n25674) );
  SDFFX1 \mem1_reg[246][13]  ( .D(n16481), .SI(\mem1[246][12] ), .SE(test_se), 
        .CLK(n1416), .Q(\mem1[246][13] ), .QN(n25675) );
  SDFFX1 \mem1_reg[246][12]  ( .D(n16480), .SI(\mem1[246][11] ), .SE(test_se), 
        .CLK(n1416), .Q(\mem1[246][12] ), .QN(n25676) );
  SDFFX1 \mem1_reg[246][11]  ( .D(n16479), .SI(\mem1[246][10] ), .SE(test_se), 
        .CLK(n1416), .Q(\mem1[246][11] ), .QN(n25677) );
  SDFFX1 \mem1_reg[246][10]  ( .D(n16478), .SI(\mem1[246][9] ), .SE(test_se), 
        .CLK(n1416), .Q(\mem1[246][10] ), .QN(n25678) );
  SDFFX1 \mem1_reg[246][9]  ( .D(n16477), .SI(\mem1[246][8] ), .SE(test_se), 
        .CLK(n1417), .Q(\mem1[246][9] ), .QN(n25679) );
  SDFFX1 \mem1_reg[246][8]  ( .D(n16476), .SI(\mem1[245][15] ), .SE(test_se), 
        .CLK(n1417), .Q(\mem1[246][8] ), .QN(n25680) );
  SDFFX1 \mem1_reg[245][15]  ( .D(n16475), .SI(\mem1[245][14] ), .SE(test_se), 
        .CLK(n1417), .Q(\mem1[245][15] ), .QN(n25681) );
  SDFFX1 \mem1_reg[245][14]  ( .D(n16474), .SI(\mem1[245][13] ), .SE(test_se), 
        .CLK(n1417), .Q(\mem1[245][14] ), .QN(n25682) );
  SDFFX1 \mem1_reg[245][13]  ( .D(n16473), .SI(\mem1[245][12] ), .SE(test_se), 
        .CLK(n1417), .Q(\mem1[245][13] ), .QN(n25683) );
  SDFFX1 \mem1_reg[245][12]  ( .D(n16472), .SI(\mem1[245][11] ), .SE(test_se), 
        .CLK(n1417), .Q(\mem1[245][12] ), .QN(n25684) );
  SDFFX1 \mem1_reg[245][11]  ( .D(n16471), .SI(\mem1[245][10] ), .SE(test_se), 
        .CLK(n1417), .Q(\mem1[245][11] ), .QN(n25685) );
  SDFFX1 \mem1_reg[245][10]  ( .D(n16470), .SI(\mem1[245][9] ), .SE(test_se), 
        .CLK(n1417), .Q(\mem1[245][10] ), .QN(n25686) );
  SDFFX1 \mem1_reg[245][9]  ( .D(n16469), .SI(\mem1[245][8] ), .SE(test_se), 
        .CLK(n1417), .Q(\mem1[245][9] ), .QN(n25687) );
  SDFFX1 \mem1_reg[245][8]  ( .D(n16468), .SI(\mem1[244][15] ), .SE(test_se), 
        .CLK(n1417), .Q(\mem1[245][8] ), .QN(n25688) );
  SDFFX1 \mem1_reg[244][15]  ( .D(n16467), .SI(\mem1[244][14] ), .SE(test_se), 
        .CLK(n1417), .Q(\mem1[244][15] ), .QN(n25689) );
  SDFFX1 \mem1_reg[244][14]  ( .D(n16466), .SI(\mem1[244][13] ), .SE(test_se), 
        .CLK(n1417), .Q(\mem1[244][14] ), .QN(n25690) );
  SDFFX1 \mem1_reg[244][13]  ( .D(n16465), .SI(\mem1[244][12] ), .SE(test_se), 
        .CLK(n1418), .Q(\mem1[244][13] ), .QN(n25691) );
  SDFFX1 \mem1_reg[244][12]  ( .D(n16464), .SI(\mem1[244][11] ), .SE(test_se), 
        .CLK(n1418), .Q(\mem1[244][12] ), .QN(n25692) );
  SDFFX1 \mem1_reg[244][11]  ( .D(n16463), .SI(\mem1[244][10] ), .SE(test_se), 
        .CLK(n1418), .Q(\mem1[244][11] ), .QN(n25693) );
  SDFFX1 \mem1_reg[244][10]  ( .D(n16462), .SI(\mem1[244][9] ), .SE(test_se), 
        .CLK(n1418), .Q(\mem1[244][10] ), .QN(n25694) );
  SDFFX1 \mem1_reg[244][9]  ( .D(n16461), .SI(\mem1[244][8] ), .SE(test_se), 
        .CLK(n1418), .Q(\mem1[244][9] ), .QN(n25695) );
  SDFFX1 \mem1_reg[244][8]  ( .D(n16460), .SI(\mem1[243][15] ), .SE(test_se), 
        .CLK(n1418), .Q(\mem1[244][8] ), .QN(n25696) );
  SDFFX1 \mem1_reg[243][15]  ( .D(n16459), .SI(\mem1[243][14] ), .SE(test_se), 
        .CLK(n1418), .Q(\mem1[243][15] ), .QN(n25697) );
  SDFFX1 \mem1_reg[243][14]  ( .D(n16458), .SI(\mem1[243][13] ), .SE(test_se), 
        .CLK(n1418), .Q(\mem1[243][14] ), .QN(n25698) );
  SDFFX1 \mem1_reg[243][13]  ( .D(n16457), .SI(\mem1[243][12] ), .SE(test_se), 
        .CLK(n1418), .Q(\mem1[243][13] ), .QN(n25699) );
  SDFFX1 \mem1_reg[243][12]  ( .D(n16456), .SI(\mem1[243][11] ), .SE(test_se), 
        .CLK(n1418), .Q(\mem1[243][12] ), .QN(n25700) );
  SDFFX1 \mem1_reg[243][11]  ( .D(n16455), .SI(\mem1[243][10] ), .SE(test_se), 
        .CLK(n1418), .Q(\mem1[243][11] ), .QN(n25701) );
  SDFFX1 \mem1_reg[243][10]  ( .D(n16454), .SI(\mem1[243][9] ), .SE(test_se), 
        .CLK(n1418), .Q(\mem1[243][10] ), .QN(n25702) );
  SDFFX1 \mem1_reg[243][9]  ( .D(n16453), .SI(\mem1[243][8] ), .SE(test_se), 
        .CLK(n1419), .Q(\mem1[243][9] ), .QN(n25703) );
  SDFFX1 \mem1_reg[243][8]  ( .D(n16452), .SI(\mem1[242][15] ), .SE(test_se), 
        .CLK(n1419), .Q(\mem1[243][8] ), .QN(n25704) );
  SDFFX1 \mem1_reg[242][15]  ( .D(n16451), .SI(\mem1[242][14] ), .SE(test_se), 
        .CLK(n1419), .Q(\mem1[242][15] ), .QN(n25705) );
  SDFFX1 \mem1_reg[242][14]  ( .D(n16450), .SI(\mem1[242][13] ), .SE(test_se), 
        .CLK(n1419), .Q(\mem1[242][14] ), .QN(n25706) );
  SDFFX1 \mem1_reg[242][13]  ( .D(n16449), .SI(\mem1[242][12] ), .SE(test_se), 
        .CLK(n1419), .Q(\mem1[242][13] ), .QN(n25707) );
  SDFFX1 \mem1_reg[242][12]  ( .D(n16448), .SI(\mem1[242][11] ), .SE(test_se), 
        .CLK(n1419), .Q(\mem1[242][12] ), .QN(n25708) );
  SDFFX1 \mem1_reg[242][11]  ( .D(n16447), .SI(\mem1[242][10] ), .SE(test_se), 
        .CLK(n1419), .Q(\mem1[242][11] ), .QN(n25709) );
  SDFFX1 \mem1_reg[242][10]  ( .D(n16446), .SI(\mem1[242][9] ), .SE(test_se), 
        .CLK(n1419), .Q(\mem1[242][10] ), .QN(n25710) );
  SDFFX1 \mem1_reg[242][9]  ( .D(n16445), .SI(\mem1[242][8] ), .SE(test_se), 
        .CLK(n1419), .Q(\mem1[242][9] ), .QN(n25711) );
  SDFFX1 \mem1_reg[242][8]  ( .D(n16444), .SI(\mem1[241][15] ), .SE(test_se), 
        .CLK(n1419), .Q(\mem1[242][8] ), .QN(n25712) );
  SDFFX1 \mem1_reg[241][15]  ( .D(n16443), .SI(\mem1[241][14] ), .SE(test_se), 
        .CLK(n1419), .Q(\mem1[241][15] ), .QN(n25713) );
  SDFFX1 \mem1_reg[241][14]  ( .D(n16442), .SI(\mem1[241][13] ), .SE(test_se), 
        .CLK(n1419), .Q(\mem1[241][14] ), .QN(n25714) );
  SDFFX1 \mem1_reg[241][13]  ( .D(n16441), .SI(\mem1[241][12] ), .SE(test_se), 
        .CLK(n1420), .Q(\mem1[241][13] ), .QN(n25715) );
  SDFFX1 \mem1_reg[241][12]  ( .D(n16440), .SI(\mem1[241][11] ), .SE(test_se), 
        .CLK(n1420), .Q(\mem1[241][12] ), .QN(n25716) );
  SDFFX1 \mem1_reg[241][11]  ( .D(n16439), .SI(\mem1[241][10] ), .SE(test_se), 
        .CLK(n1420), .Q(\mem1[241][11] ), .QN(n25717) );
  SDFFX1 \mem1_reg[241][10]  ( .D(n16438), .SI(\mem1[241][9] ), .SE(test_se), 
        .CLK(n1420), .Q(\mem1[241][10] ), .QN(n25718) );
  SDFFX1 \mem1_reg[241][9]  ( .D(n16437), .SI(\mem1[241][8] ), .SE(test_se), 
        .CLK(n1420), .Q(\mem1[241][9] ), .QN(n25719) );
  SDFFX1 \mem1_reg[241][8]  ( .D(n16436), .SI(\mem1[240][15] ), .SE(test_se), 
        .CLK(n1420), .Q(\mem1[241][8] ), .QN(n25720) );
  SDFFX1 \mem1_reg[240][15]  ( .D(n16435), .SI(\mem1[240][14] ), .SE(test_se), 
        .CLK(n1420), .Q(\mem1[240][15] ), .QN(n25721) );
  SDFFX1 \mem1_reg[240][14]  ( .D(n16434), .SI(\mem1[240][13] ), .SE(test_se), 
        .CLK(n1420), .Q(\mem1[240][14] ), .QN(n25722) );
  SDFFX1 \mem1_reg[240][13]  ( .D(n16433), .SI(\mem1[240][12] ), .SE(test_se), 
        .CLK(n1420), .Q(\mem1[240][13] ), .QN(n25723) );
  SDFFX1 \mem1_reg[240][12]  ( .D(n16432), .SI(\mem1[240][11] ), .SE(test_se), 
        .CLK(n1420), .Q(\mem1[240][12] ), .QN(n25724) );
  SDFFX1 \mem1_reg[240][11]  ( .D(n16431), .SI(\mem1[240][10] ), .SE(test_se), 
        .CLK(n1420), .Q(\mem1[240][11] ), .QN(n25725) );
  SDFFX1 \mem1_reg[240][10]  ( .D(n16430), .SI(\mem1[240][9] ), .SE(test_se), 
        .CLK(n1420), .Q(\mem1[240][10] ), .QN(n25726) );
  SDFFX1 \mem1_reg[240][9]  ( .D(n16429), .SI(\mem1[240][8] ), .SE(test_se), 
        .CLK(n1421), .Q(\mem1[240][9] ), .QN(n25727) );
  SDFFX1 \mem1_reg[240][8]  ( .D(n16428), .SI(\mem1[239][15] ), .SE(test_se), 
        .CLK(n1421), .Q(\mem1[240][8] ), .QN(n25728) );
  SDFFX1 \mem1_reg[239][15]  ( .D(n16427), .SI(\mem1[239][14] ), .SE(test_se), 
        .CLK(n1421), .Q(\mem1[239][15] ), .QN(n25729) );
  SDFFX1 \mem1_reg[239][14]  ( .D(n16426), .SI(\mem1[239][13] ), .SE(test_se), 
        .CLK(n1421), .Q(\mem1[239][14] ), .QN(n25730) );
  SDFFX1 \mem1_reg[239][13]  ( .D(n16425), .SI(\mem1[239][12] ), .SE(test_se), 
        .CLK(n1421), .Q(\mem1[239][13] ), .QN(n25731) );
  SDFFX1 \mem1_reg[239][12]  ( .D(n16424), .SI(\mem1[239][11] ), .SE(test_se), 
        .CLK(n1421), .Q(\mem1[239][12] ), .QN(n25732) );
  SDFFX1 \mem1_reg[239][11]  ( .D(n16423), .SI(\mem1[239][10] ), .SE(test_se), 
        .CLK(n1421), .Q(\mem1[239][11] ), .QN(n25733) );
  SDFFX1 \mem1_reg[239][10]  ( .D(n16422), .SI(\mem1[239][9] ), .SE(test_se), 
        .CLK(n1421), .Q(\mem1[239][10] ), .QN(n25734) );
  SDFFX1 \mem1_reg[239][9]  ( .D(n16421), .SI(\mem1[239][8] ), .SE(test_se), 
        .CLK(n1421), .Q(\mem1[239][9] ), .QN(n25735) );
  SDFFX1 \mem1_reg[239][8]  ( .D(n16420), .SI(\mem1[238][15] ), .SE(test_se), 
        .CLK(n1421), .Q(\mem1[239][8] ), .QN(n25736) );
  SDFFX1 \mem1_reg[238][15]  ( .D(n16419), .SI(\mem1[238][14] ), .SE(test_se), 
        .CLK(n1421), .Q(\mem1[238][15] ), .QN(n25737) );
  SDFFX1 \mem1_reg[238][14]  ( .D(n16418), .SI(\mem1[238][13] ), .SE(test_se), 
        .CLK(n1421), .Q(\mem1[238][14] ), .QN(n25738) );
  SDFFX1 \mem1_reg[238][13]  ( .D(n16417), .SI(\mem1[238][12] ), .SE(test_se), 
        .CLK(n1422), .Q(\mem1[238][13] ), .QN(n25739) );
  SDFFX1 \mem1_reg[238][12]  ( .D(n16416), .SI(\mem1[238][11] ), .SE(test_se), 
        .CLK(n1422), .Q(\mem1[238][12] ), .QN(n25740) );
  SDFFX1 \mem1_reg[238][11]  ( .D(n16415), .SI(\mem1[238][10] ), .SE(test_se), 
        .CLK(n1422), .Q(\mem1[238][11] ), .QN(n25741) );
  SDFFX1 \mem1_reg[238][10]  ( .D(n16414), .SI(\mem1[238][9] ), .SE(test_se), 
        .CLK(n1422), .Q(\mem1[238][10] ), .QN(n25742) );
  SDFFX1 \mem1_reg[238][9]  ( .D(n16413), .SI(\mem1[238][8] ), .SE(test_se), 
        .CLK(n1422), .Q(\mem1[238][9] ), .QN(n25743) );
  SDFFX1 \mem1_reg[238][8]  ( .D(n16412), .SI(\mem1[237][15] ), .SE(test_se), 
        .CLK(n1422), .Q(\mem1[238][8] ), .QN(n25744) );
  SDFFX1 \mem1_reg[237][15]  ( .D(n16411), .SI(\mem1[237][14] ), .SE(test_se), 
        .CLK(n1422), .Q(\mem1[237][15] ), .QN(n25745) );
  SDFFX1 \mem1_reg[237][14]  ( .D(n16410), .SI(\mem1[237][13] ), .SE(test_se), 
        .CLK(n1422), .Q(\mem1[237][14] ), .QN(n25746) );
  SDFFX1 \mem1_reg[237][13]  ( .D(n16409), .SI(\mem1[237][12] ), .SE(test_se), 
        .CLK(n1422), .Q(\mem1[237][13] ), .QN(n25747) );
  SDFFX1 \mem1_reg[237][12]  ( .D(n16408), .SI(\mem1[237][11] ), .SE(test_se), 
        .CLK(n1422), .Q(\mem1[237][12] ), .QN(n25748) );
  SDFFX1 \mem1_reg[237][11]  ( .D(n16407), .SI(\mem1[237][10] ), .SE(test_se), 
        .CLK(n1422), .Q(\mem1[237][11] ), .QN(n25749) );
  SDFFX1 \mem1_reg[237][10]  ( .D(n16406), .SI(\mem1[237][9] ), .SE(test_se), 
        .CLK(n1422), .Q(\mem1[237][10] ), .QN(n25750) );
  SDFFX1 \mem1_reg[237][9]  ( .D(n16405), .SI(\mem1[237][8] ), .SE(test_se), 
        .CLK(n1423), .Q(\mem1[237][9] ), .QN(n25751) );
  SDFFX1 \mem1_reg[237][8]  ( .D(n16404), .SI(\mem1[236][15] ), .SE(test_se), 
        .CLK(n1423), .Q(\mem1[237][8] ), .QN(n25752) );
  SDFFX1 \mem1_reg[236][15]  ( .D(n16403), .SI(\mem1[236][14] ), .SE(test_se), 
        .CLK(n1423), .Q(\mem1[236][15] ), .QN(n25753) );
  SDFFX1 \mem1_reg[236][14]  ( .D(n16402), .SI(\mem1[236][13] ), .SE(test_se), 
        .CLK(n1423), .Q(\mem1[236][14] ), .QN(n25754) );
  SDFFX1 \mem1_reg[236][13]  ( .D(n16401), .SI(\mem1[236][12] ), .SE(test_se), 
        .CLK(n1423), .Q(\mem1[236][13] ), .QN(n25755) );
  SDFFX1 \mem1_reg[236][12]  ( .D(n16400), .SI(\mem1[236][11] ), .SE(test_se), 
        .CLK(n1423), .Q(\mem1[236][12] ), .QN(n25756) );
  SDFFX1 \mem1_reg[236][11]  ( .D(n16399), .SI(\mem1[236][10] ), .SE(test_se), 
        .CLK(n1423), .Q(\mem1[236][11] ), .QN(n25757) );
  SDFFX1 \mem1_reg[236][10]  ( .D(n16398), .SI(\mem1[236][9] ), .SE(test_se), 
        .CLK(n1423), .Q(\mem1[236][10] ), .QN(n25758) );
  SDFFX1 \mem1_reg[236][9]  ( .D(n16397), .SI(\mem1[236][8] ), .SE(test_se), 
        .CLK(n1423), .Q(\mem1[236][9] ), .QN(n25759) );
  SDFFX1 \mem1_reg[236][8]  ( .D(n16396), .SI(\mem1[235][15] ), .SE(test_se), 
        .CLK(n1423), .Q(\mem1[236][8] ), .QN(n25760) );
  SDFFX1 \mem1_reg[235][15]  ( .D(n16395), .SI(\mem1[235][14] ), .SE(test_se), 
        .CLK(n1423), .Q(\mem1[235][15] ), .QN(n25761) );
  SDFFX1 \mem1_reg[235][14]  ( .D(n16394), .SI(\mem1[235][13] ), .SE(test_se), 
        .CLK(n1423), .Q(\mem1[235][14] ), .QN(n25762) );
  SDFFX1 \mem1_reg[235][13]  ( .D(n16393), .SI(\mem1[235][12] ), .SE(test_se), 
        .CLK(n1424), .Q(\mem1[235][13] ), .QN(n25763) );
  SDFFX1 \mem1_reg[235][12]  ( .D(n16392), .SI(\mem1[235][11] ), .SE(test_se), 
        .CLK(n1424), .Q(\mem1[235][12] ), .QN(n25764) );
  SDFFX1 \mem1_reg[235][11]  ( .D(n16391), .SI(\mem1[235][10] ), .SE(test_se), 
        .CLK(n1424), .Q(\mem1[235][11] ), .QN(n25765) );
  SDFFX1 \mem1_reg[235][10]  ( .D(n16390), .SI(\mem1[235][9] ), .SE(test_se), 
        .CLK(n1424), .Q(\mem1[235][10] ), .QN(n25766) );
  SDFFX1 \mem1_reg[235][9]  ( .D(n16389), .SI(\mem1[235][8] ), .SE(test_se), 
        .CLK(n1424), .Q(\mem1[235][9] ), .QN(n25767) );
  SDFFX1 \mem1_reg[235][8]  ( .D(n16388), .SI(\mem1[234][15] ), .SE(test_se), 
        .CLK(n1424), .Q(\mem1[235][8] ), .QN(n25768) );
  SDFFX1 \mem1_reg[234][15]  ( .D(n16387), .SI(\mem1[234][14] ), .SE(test_se), 
        .CLK(n1424), .Q(\mem1[234][15] ), .QN(n25769) );
  SDFFX1 \mem1_reg[234][14]  ( .D(n16386), .SI(\mem1[234][13] ), .SE(test_se), 
        .CLK(n1424), .Q(\mem1[234][14] ), .QN(n25770) );
  SDFFX1 \mem1_reg[234][13]  ( .D(n16385), .SI(\mem1[234][12] ), .SE(test_se), 
        .CLK(n1424), .Q(\mem1[234][13] ), .QN(n25771) );
  SDFFX1 \mem1_reg[234][12]  ( .D(n16384), .SI(\mem1[234][11] ), .SE(test_se), 
        .CLK(n1424), .Q(\mem1[234][12] ), .QN(n25772) );
  SDFFX1 \mem1_reg[234][11]  ( .D(n16383), .SI(\mem1[234][10] ), .SE(test_se), 
        .CLK(n1424), .Q(\mem1[234][11] ), .QN(n25773) );
  SDFFX1 \mem1_reg[234][10]  ( .D(n16382), .SI(\mem1[234][9] ), .SE(test_se), 
        .CLK(n1424), .Q(\mem1[234][10] ), .QN(n25774) );
  SDFFX1 \mem1_reg[234][9]  ( .D(n16381), .SI(\mem1[234][8] ), .SE(test_se), 
        .CLK(n1425), .Q(\mem1[234][9] ), .QN(n25775) );
  SDFFX1 \mem1_reg[234][8]  ( .D(n16380), .SI(\mem1[233][15] ), .SE(test_se), 
        .CLK(n1425), .Q(\mem1[234][8] ), .QN(n25776) );
  SDFFX1 \mem1_reg[233][15]  ( .D(n16379), .SI(\mem1[233][14] ), .SE(test_se), 
        .CLK(n1425), .Q(\mem1[233][15] ), .QN(n25777) );
  SDFFX1 \mem1_reg[233][14]  ( .D(n16378), .SI(\mem1[233][13] ), .SE(test_se), 
        .CLK(n1425), .Q(\mem1[233][14] ), .QN(n25778) );
  SDFFX1 \mem1_reg[233][13]  ( .D(n16377), .SI(\mem1[233][12] ), .SE(test_se), 
        .CLK(n1425), .Q(\mem1[233][13] ), .QN(n25779) );
  SDFFX1 \mem1_reg[233][12]  ( .D(n16376), .SI(\mem1[233][11] ), .SE(test_se), 
        .CLK(n1425), .Q(\mem1[233][12] ), .QN(n25780) );
  SDFFX1 \mem1_reg[233][11]  ( .D(n16375), .SI(\mem1[233][10] ), .SE(test_se), 
        .CLK(n1425), .Q(\mem1[233][11] ), .QN(n25781) );
  SDFFX1 \mem1_reg[233][10]  ( .D(n16374), .SI(\mem1[233][9] ), .SE(test_se), 
        .CLK(n1425), .Q(\mem1[233][10] ), .QN(n25782) );
  SDFFX1 \mem1_reg[233][9]  ( .D(n16373), .SI(\mem1[233][8] ), .SE(test_se), 
        .CLK(n1425), .Q(\mem1[233][9] ), .QN(n25783) );
  SDFFX1 \mem1_reg[233][8]  ( .D(n16372), .SI(\mem1[232][15] ), .SE(test_se), 
        .CLK(n1425), .Q(\mem1[233][8] ), .QN(n25784) );
  SDFFX1 \mem1_reg[232][15]  ( .D(n16371), .SI(\mem1[232][14] ), .SE(test_se), 
        .CLK(n1425), .Q(\mem1[232][15] ), .QN(n25785) );
  SDFFX1 \mem1_reg[232][14]  ( .D(n16370), .SI(\mem1[232][13] ), .SE(test_se), 
        .CLK(n1425), .Q(\mem1[232][14] ), .QN(n25786) );
  SDFFX1 \mem1_reg[232][13]  ( .D(n16369), .SI(\mem1[232][12] ), .SE(test_se), 
        .CLK(n1426), .Q(\mem1[232][13] ), .QN(n25787) );
  SDFFX1 \mem1_reg[232][12]  ( .D(n16368), .SI(\mem1[232][11] ), .SE(test_se), 
        .CLK(n1426), .Q(\mem1[232][12] ), .QN(n25788) );
  SDFFX1 \mem1_reg[232][11]  ( .D(n16367), .SI(\mem1[232][10] ), .SE(test_se), 
        .CLK(n1426), .Q(\mem1[232][11] ), .QN(n25789) );
  SDFFX1 \mem1_reg[232][10]  ( .D(n16366), .SI(\mem1[232][9] ), .SE(test_se), 
        .CLK(n1426), .Q(\mem1[232][10] ), .QN(n25790) );
  SDFFX1 \mem1_reg[232][9]  ( .D(n16365), .SI(\mem1[232][8] ), .SE(test_se), 
        .CLK(n1426), .Q(\mem1[232][9] ), .QN(n25791) );
  SDFFX1 \mem1_reg[232][8]  ( .D(n16364), .SI(\mem1[231][15] ), .SE(test_se), 
        .CLK(n1426), .Q(\mem1[232][8] ), .QN(n25792) );
  SDFFX1 \mem1_reg[231][15]  ( .D(n16363), .SI(\mem1[231][14] ), .SE(test_se), 
        .CLK(n1426), .Q(\mem1[231][15] ), .QN(n25793) );
  SDFFX1 \mem1_reg[231][14]  ( .D(n16362), .SI(\mem1[231][13] ), .SE(test_se), 
        .CLK(n1426), .Q(\mem1[231][14] ), .QN(n25794) );
  SDFFX1 \mem1_reg[231][13]  ( .D(n16361), .SI(\mem1[231][12] ), .SE(test_se), 
        .CLK(n1426), .Q(\mem1[231][13] ), .QN(n25795) );
  SDFFX1 \mem1_reg[231][12]  ( .D(n16360), .SI(\mem1[231][11] ), .SE(test_se), 
        .CLK(n1426), .Q(\mem1[231][12] ), .QN(n25796) );
  SDFFX1 \mem1_reg[231][11]  ( .D(n16359), .SI(\mem1[231][10] ), .SE(test_se), 
        .CLK(n1426), .Q(\mem1[231][11] ), .QN(n25797) );
  SDFFX1 \mem1_reg[231][10]  ( .D(n16358), .SI(\mem1[231][9] ), .SE(test_se), 
        .CLK(n1426), .Q(\mem1[231][10] ), .QN(n25798) );
  SDFFX1 \mem1_reg[231][9]  ( .D(n16357), .SI(\mem1[231][8] ), .SE(test_se), 
        .CLK(n1427), .Q(\mem1[231][9] ), .QN(n25799) );
  SDFFX1 \mem1_reg[231][8]  ( .D(n16356), .SI(\mem1[230][15] ), .SE(test_se), 
        .CLK(n1427), .Q(\mem1[231][8] ), .QN(n25800) );
  SDFFX1 \mem1_reg[230][15]  ( .D(n16355), .SI(\mem1[230][14] ), .SE(test_se), 
        .CLK(n1427), .Q(\mem1[230][15] ), .QN(n25801) );
  SDFFX1 \mem1_reg[230][14]  ( .D(n16354), .SI(\mem1[230][13] ), .SE(test_se), 
        .CLK(n1427), .Q(\mem1[230][14] ), .QN(n25802) );
  SDFFX1 \mem1_reg[230][13]  ( .D(n16353), .SI(\mem1[230][12] ), .SE(test_se), 
        .CLK(n1427), .Q(\mem1[230][13] ), .QN(n25803) );
  SDFFX1 \mem1_reg[230][12]  ( .D(n16352), .SI(\mem1[230][11] ), .SE(test_se), 
        .CLK(n1427), .Q(\mem1[230][12] ), .QN(n25804) );
  SDFFX1 \mem1_reg[230][11]  ( .D(n16351), .SI(\mem1[230][10] ), .SE(test_se), 
        .CLK(n1427), .Q(\mem1[230][11] ), .QN(n25805) );
  SDFFX1 \mem1_reg[230][10]  ( .D(n16350), .SI(\mem1[230][9] ), .SE(test_se), 
        .CLK(n1427), .Q(\mem1[230][10] ), .QN(n25806) );
  SDFFX1 \mem1_reg[230][9]  ( .D(n16349), .SI(\mem1[230][8] ), .SE(test_se), 
        .CLK(n1427), .Q(\mem1[230][9] ), .QN(n25807) );
  SDFFX1 \mem1_reg[230][8]  ( .D(n16348), .SI(\mem1[229][15] ), .SE(test_se), 
        .CLK(n1427), .Q(\mem1[230][8] ), .QN(n25808) );
  SDFFX1 \mem1_reg[229][15]  ( .D(n16347), .SI(\mem1[229][14] ), .SE(test_se), 
        .CLK(n1427), .Q(\mem1[229][15] ), .QN(n25809) );
  SDFFX1 \mem1_reg[229][14]  ( .D(n16346), .SI(\mem1[229][13] ), .SE(test_se), 
        .CLK(n1427), .Q(\mem1[229][14] ), .QN(n25810) );
  SDFFX1 \mem1_reg[229][13]  ( .D(n16345), .SI(\mem1[229][12] ), .SE(test_se), 
        .CLK(n1428), .Q(\mem1[229][13] ), .QN(n25811) );
  SDFFX1 \mem1_reg[229][12]  ( .D(n16344), .SI(\mem1[229][11] ), .SE(test_se), 
        .CLK(n1428), .Q(\mem1[229][12] ), .QN(n25812) );
  SDFFX1 \mem1_reg[229][11]  ( .D(n16343), .SI(\mem1[229][10] ), .SE(test_se), 
        .CLK(n1428), .Q(\mem1[229][11] ), .QN(n25813) );
  SDFFX1 \mem1_reg[229][10]  ( .D(n16342), .SI(\mem1[229][9] ), .SE(test_se), 
        .CLK(n1428), .Q(\mem1[229][10] ), .QN(n25814) );
  SDFFX1 \mem1_reg[229][9]  ( .D(n16341), .SI(\mem1[229][8] ), .SE(test_se), 
        .CLK(n1428), .Q(\mem1[229][9] ), .QN(n25815) );
  SDFFX1 \mem1_reg[229][8]  ( .D(n16340), .SI(\mem1[228][15] ), .SE(test_se), 
        .CLK(n1428), .Q(\mem1[229][8] ), .QN(n25816) );
  SDFFX1 \mem1_reg[228][15]  ( .D(n16339), .SI(\mem1[228][14] ), .SE(test_se), 
        .CLK(n1428), .Q(\mem1[228][15] ), .QN(n25817) );
  SDFFX1 \mem1_reg[228][14]  ( .D(n16338), .SI(\mem1[228][13] ), .SE(test_se), 
        .CLK(n1428), .Q(\mem1[228][14] ), .QN(n25818) );
  SDFFX1 \mem1_reg[228][13]  ( .D(n16337), .SI(\mem1[228][12] ), .SE(test_se), 
        .CLK(n1428), .Q(\mem1[228][13] ), .QN(n25819) );
  SDFFX1 \mem1_reg[228][12]  ( .D(n16336), .SI(\mem1[228][11] ), .SE(test_se), 
        .CLK(n1428), .Q(\mem1[228][12] ), .QN(n25820) );
  SDFFX1 \mem1_reg[228][11]  ( .D(n16335), .SI(\mem1[228][10] ), .SE(test_se), 
        .CLK(n1428), .Q(\mem1[228][11] ), .QN(n25821) );
  SDFFX1 \mem1_reg[228][10]  ( .D(n16334), .SI(\mem1[228][9] ), .SE(test_se), 
        .CLK(n1428), .Q(\mem1[228][10] ), .QN(n25822) );
  SDFFX1 \mem1_reg[228][9]  ( .D(n16333), .SI(\mem1[228][8] ), .SE(test_se), 
        .CLK(n1429), .Q(\mem1[228][9] ), .QN(n25823) );
  SDFFX1 \mem1_reg[228][8]  ( .D(n16332), .SI(\mem1[227][15] ), .SE(test_se), 
        .CLK(n1429), .Q(\mem1[228][8] ), .QN(n25824) );
  SDFFX1 \mem1_reg[227][15]  ( .D(n16331), .SI(\mem1[227][14] ), .SE(test_se), 
        .CLK(n1429), .Q(\mem1[227][15] ), .QN(n25825) );
  SDFFX1 \mem1_reg[227][14]  ( .D(n16330), .SI(\mem1[227][13] ), .SE(test_se), 
        .CLK(n1429), .Q(\mem1[227][14] ), .QN(n25826) );
  SDFFX1 \mem1_reg[227][13]  ( .D(n16329), .SI(\mem1[227][12] ), .SE(test_se), 
        .CLK(n1429), .Q(\mem1[227][13] ), .QN(n25827) );
  SDFFX1 \mem1_reg[227][12]  ( .D(n16328), .SI(\mem1[227][11] ), .SE(test_se), 
        .CLK(n1429), .Q(\mem1[227][12] ), .QN(n25828) );
  SDFFX1 \mem1_reg[227][11]  ( .D(n16327), .SI(\mem1[227][10] ), .SE(test_se), 
        .CLK(n1429), .Q(\mem1[227][11] ), .QN(n25829) );
  SDFFX1 \mem1_reg[227][10]  ( .D(n16326), .SI(\mem1[227][9] ), .SE(test_se), 
        .CLK(n1429), .Q(\mem1[227][10] ), .QN(n25830) );
  SDFFX1 \mem1_reg[227][9]  ( .D(n16325), .SI(\mem1[227][8] ), .SE(test_se), 
        .CLK(n1429), .Q(\mem1[227][9] ), .QN(n25831) );
  SDFFX1 \mem1_reg[227][8]  ( .D(n16324), .SI(\mem1[226][15] ), .SE(test_se), 
        .CLK(n1429), .Q(\mem1[227][8] ), .QN(n25832) );
  SDFFX1 \mem1_reg[226][15]  ( .D(n16323), .SI(\mem1[226][14] ), .SE(test_se), 
        .CLK(n1429), .Q(\mem1[226][15] ), .QN(n25833) );
  SDFFX1 \mem1_reg[226][14]  ( .D(n16322), .SI(\mem1[226][13] ), .SE(test_se), 
        .CLK(n1429), .Q(\mem1[226][14] ), .QN(n25834) );
  SDFFX1 \mem1_reg[226][13]  ( .D(n16321), .SI(\mem1[226][12] ), .SE(test_se), 
        .CLK(n1430), .Q(\mem1[226][13] ), .QN(n25835) );
  SDFFX1 \mem1_reg[226][12]  ( .D(n16320), .SI(\mem1[226][11] ), .SE(test_se), 
        .CLK(n1430), .Q(\mem1[226][12] ), .QN(n25836) );
  SDFFX1 \mem1_reg[226][11]  ( .D(n16319), .SI(\mem1[226][10] ), .SE(test_se), 
        .CLK(n1430), .Q(\mem1[226][11] ), .QN(n25837) );
  SDFFX1 \mem1_reg[226][10]  ( .D(n16318), .SI(\mem1[226][9] ), .SE(test_se), 
        .CLK(n1430), .Q(\mem1[226][10] ), .QN(n25838) );
  SDFFX1 \mem1_reg[226][9]  ( .D(n16317), .SI(\mem1[226][8] ), .SE(test_se), 
        .CLK(n1430), .Q(\mem1[226][9] ), .QN(n25839) );
  SDFFX1 \mem1_reg[226][8]  ( .D(n16316), .SI(\mem1[225][15] ), .SE(test_se), 
        .CLK(n1430), .Q(\mem1[226][8] ), .QN(n25840) );
  SDFFX1 \mem1_reg[225][15]  ( .D(n16315), .SI(\mem1[225][14] ), .SE(test_se), 
        .CLK(n1430), .Q(\mem1[225][15] ), .QN(n25841) );
  SDFFX1 \mem1_reg[225][14]  ( .D(n16314), .SI(\mem1[225][13] ), .SE(test_se), 
        .CLK(n1430), .Q(\mem1[225][14] ), .QN(n25842) );
  SDFFX1 \mem1_reg[225][13]  ( .D(n16313), .SI(\mem1[225][12] ), .SE(test_se), 
        .CLK(n1430), .Q(\mem1[225][13] ), .QN(n25843) );
  SDFFX1 \mem1_reg[225][12]  ( .D(n16312), .SI(\mem1[225][11] ), .SE(test_se), 
        .CLK(n1430), .Q(\mem1[225][12] ), .QN(n25844) );
  SDFFX1 \mem1_reg[225][11]  ( .D(n16311), .SI(\mem1[225][10] ), .SE(test_se), 
        .CLK(n1430), .Q(\mem1[225][11] ), .QN(n25845) );
  SDFFX1 \mem1_reg[225][10]  ( .D(n16310), .SI(\mem1[225][9] ), .SE(test_se), 
        .CLK(n1430), .Q(\mem1[225][10] ), .QN(n25846) );
  SDFFX1 \mem1_reg[225][9]  ( .D(n16309), .SI(\mem1[225][8] ), .SE(test_se), 
        .CLK(n1431), .Q(\mem1[225][9] ), .QN(n25847) );
  SDFFX1 \mem1_reg[225][8]  ( .D(n16308), .SI(\mem1[224][15] ), .SE(test_se), 
        .CLK(n1431), .Q(\mem1[225][8] ), .QN(n25848) );
  SDFFX1 \mem1_reg[224][15]  ( .D(n16307), .SI(\mem1[224][14] ), .SE(test_se), 
        .CLK(n1431), .Q(\mem1[224][15] ), .QN(n25849) );
  SDFFX1 \mem1_reg[224][14]  ( .D(n16306), .SI(\mem1[224][13] ), .SE(test_se), 
        .CLK(n1431), .Q(\mem1[224][14] ), .QN(n25850) );
  SDFFX1 \mem1_reg[224][13]  ( .D(n16305), .SI(\mem1[224][12] ), .SE(test_se), 
        .CLK(n1431), .Q(\mem1[224][13] ), .QN(n25851) );
  SDFFX1 \mem1_reg[224][12]  ( .D(n16304), .SI(\mem1[224][11] ), .SE(test_se), 
        .CLK(n1431), .Q(\mem1[224][12] ), .QN(n25852) );
  SDFFX1 \mem1_reg[224][11]  ( .D(n16303), .SI(\mem1[224][10] ), .SE(test_se), 
        .CLK(n1431), .Q(\mem1[224][11] ), .QN(n25853) );
  SDFFX1 \mem1_reg[224][10]  ( .D(n16302), .SI(\mem1[224][9] ), .SE(test_se), 
        .CLK(n1431), .Q(\mem1[224][10] ), .QN(n25854) );
  SDFFX1 \mem1_reg[224][9]  ( .D(n16301), .SI(\mem1[224][8] ), .SE(test_se), 
        .CLK(n1431), .Q(\mem1[224][9] ), .QN(n25855) );
  SDFFX1 \mem1_reg[224][8]  ( .D(n16300), .SI(\mem1[223][15] ), .SE(test_se), 
        .CLK(n1431), .Q(\mem1[224][8] ), .QN(n25856) );
  SDFFX1 \mem1_reg[223][15]  ( .D(n16299), .SI(\mem1[223][14] ), .SE(test_se), 
        .CLK(n1431), .Q(\mem1[223][15] ), .QN(n25857) );
  SDFFX1 \mem1_reg[223][14]  ( .D(n16298), .SI(\mem1[223][13] ), .SE(test_se), 
        .CLK(n1431), .Q(\mem1[223][14] ), .QN(n25858) );
  SDFFX1 \mem1_reg[223][13]  ( .D(n16297), .SI(\mem1[223][12] ), .SE(test_se), 
        .CLK(n1432), .Q(\mem1[223][13] ), .QN(n25859) );
  SDFFX1 \mem1_reg[223][12]  ( .D(n16296), .SI(\mem1[223][11] ), .SE(test_se), 
        .CLK(n1432), .Q(\mem1[223][12] ), .QN(n25860) );
  SDFFX1 \mem1_reg[223][11]  ( .D(n16295), .SI(\mem1[223][10] ), .SE(test_se), 
        .CLK(n1432), .Q(\mem1[223][11] ), .QN(n25861) );
  SDFFX1 \mem1_reg[223][10]  ( .D(n16294), .SI(\mem1[223][9] ), .SE(test_se), 
        .CLK(n1432), .Q(\mem1[223][10] ), .QN(n25862) );
  SDFFX1 \mem1_reg[223][9]  ( .D(n16293), .SI(\mem1[223][8] ), .SE(test_se), 
        .CLK(n1432), .Q(\mem1[223][9] ), .QN(n25863) );
  SDFFX1 \mem1_reg[223][8]  ( .D(n16292), .SI(\mem1[222][15] ), .SE(test_se), 
        .CLK(n1432), .Q(\mem1[223][8] ), .QN(n25864) );
  SDFFX1 \mem1_reg[222][15]  ( .D(n16291), .SI(\mem1[222][14] ), .SE(test_se), 
        .CLK(n1432), .Q(\mem1[222][15] ), .QN(n25865) );
  SDFFX1 \mem1_reg[222][14]  ( .D(n16290), .SI(\mem1[222][13] ), .SE(test_se), 
        .CLK(n1432), .Q(\mem1[222][14] ), .QN(n25866) );
  SDFFX1 \mem1_reg[222][13]  ( .D(n16289), .SI(\mem1[222][12] ), .SE(test_se), 
        .CLK(n1432), .Q(\mem1[222][13] ), .QN(n25867) );
  SDFFX1 \mem1_reg[222][12]  ( .D(n16288), .SI(\mem1[222][11] ), .SE(test_se), 
        .CLK(n1432), .Q(\mem1[222][12] ), .QN(n25868) );
  SDFFX1 \mem1_reg[222][11]  ( .D(n16287), .SI(\mem1[222][10] ), .SE(test_se), 
        .CLK(n1432), .Q(\mem1[222][11] ), .QN(n25869) );
  SDFFX1 \mem1_reg[222][10]  ( .D(n16286), .SI(\mem1[222][9] ), .SE(test_se), 
        .CLK(n1432), .Q(\mem1[222][10] ), .QN(n25870) );
  SDFFX1 \mem1_reg[222][9]  ( .D(n16285), .SI(\mem1[222][8] ), .SE(test_se), 
        .CLK(n1433), .Q(\mem1[222][9] ), .QN(n25871) );
  SDFFX1 \mem1_reg[222][8]  ( .D(n16284), .SI(\mem1[221][15] ), .SE(test_se), 
        .CLK(n1433), .Q(\mem1[222][8] ), .QN(n25872) );
  SDFFX1 \mem1_reg[221][15]  ( .D(n16283), .SI(\mem1[221][14] ), .SE(test_se), 
        .CLK(n1433), .Q(\mem1[221][15] ), .QN(n25873) );
  SDFFX1 \mem1_reg[221][14]  ( .D(n16282), .SI(\mem1[221][13] ), .SE(test_se), 
        .CLK(n1433), .Q(\mem1[221][14] ), .QN(n25874) );
  SDFFX1 \mem1_reg[221][13]  ( .D(n16281), .SI(\mem1[221][12] ), .SE(test_se), 
        .CLK(n1433), .Q(\mem1[221][13] ), .QN(n25875) );
  SDFFX1 \mem1_reg[221][12]  ( .D(n16280), .SI(\mem1[221][11] ), .SE(test_se), 
        .CLK(n1433), .Q(\mem1[221][12] ), .QN(n25876) );
  SDFFX1 \mem1_reg[221][11]  ( .D(n16279), .SI(\mem1[221][10] ), .SE(test_se), 
        .CLK(n1433), .Q(\mem1[221][11] ), .QN(n25877) );
  SDFFX1 \mem1_reg[221][10]  ( .D(n16278), .SI(\mem1[221][9] ), .SE(test_se), 
        .CLK(n1433), .Q(\mem1[221][10] ), .QN(n25878) );
  SDFFX1 \mem1_reg[221][9]  ( .D(n16277), .SI(\mem1[221][8] ), .SE(test_se), 
        .CLK(n1433), .Q(\mem1[221][9] ), .QN(n25879) );
  SDFFX1 \mem1_reg[221][8]  ( .D(n16276), .SI(\mem1[220][15] ), .SE(test_se), 
        .CLK(n1433), .Q(\mem1[221][8] ), .QN(n25880) );
  SDFFX1 \mem1_reg[220][15]  ( .D(n16275), .SI(\mem1[220][14] ), .SE(test_se), 
        .CLK(n1433), .Q(\mem1[220][15] ), .QN(n25881) );
  SDFFX1 \mem1_reg[220][14]  ( .D(n16274), .SI(\mem1[220][13] ), .SE(test_se), 
        .CLK(n1433), .Q(\mem1[220][14] ), .QN(n25882) );
  SDFFX1 \mem1_reg[220][13]  ( .D(n16273), .SI(\mem1[220][12] ), .SE(test_se), 
        .CLK(n1434), .Q(\mem1[220][13] ), .QN(n25883) );
  SDFFX1 \mem1_reg[220][12]  ( .D(n16272), .SI(\mem1[220][11] ), .SE(test_se), 
        .CLK(n1434), .Q(\mem1[220][12] ), .QN(n25884) );
  SDFFX1 \mem1_reg[220][11]  ( .D(n16271), .SI(\mem1[220][10] ), .SE(test_se), 
        .CLK(n1434), .Q(\mem1[220][11] ), .QN(n25885) );
  SDFFX1 \mem1_reg[220][10]  ( .D(n16270), .SI(\mem1[220][9] ), .SE(test_se), 
        .CLK(n1434), .Q(\mem1[220][10] ), .QN(n25886) );
  SDFFX1 \mem1_reg[220][9]  ( .D(n16269), .SI(\mem1[220][8] ), .SE(test_se), 
        .CLK(n1434), .Q(\mem1[220][9] ), .QN(n25887) );
  SDFFX1 \mem1_reg[220][8]  ( .D(n16268), .SI(\mem1[219][15] ), .SE(test_se), 
        .CLK(n1434), .Q(\mem1[220][8] ), .QN(n25888) );
  SDFFX1 \mem1_reg[219][15]  ( .D(n16267), .SI(\mem1[219][14] ), .SE(test_se), 
        .CLK(n1434), .Q(\mem1[219][15] ), .QN(n25889) );
  SDFFX1 \mem1_reg[219][14]  ( .D(n16266), .SI(\mem1[219][13] ), .SE(test_se), 
        .CLK(n1434), .Q(\mem1[219][14] ), .QN(n25890) );
  SDFFX1 \mem1_reg[219][13]  ( .D(n16265), .SI(\mem1[219][12] ), .SE(test_se), 
        .CLK(n1434), .Q(\mem1[219][13] ), .QN(n25891) );
  SDFFX1 \mem1_reg[219][12]  ( .D(n16264), .SI(\mem1[219][11] ), .SE(test_se), 
        .CLK(n1434), .Q(\mem1[219][12] ), .QN(n25892) );
  SDFFX1 \mem1_reg[219][11]  ( .D(n16263), .SI(\mem1[219][10] ), .SE(test_se), 
        .CLK(n1434), .Q(\mem1[219][11] ), .QN(n25893) );
  SDFFX1 \mem1_reg[219][10]  ( .D(n16262), .SI(\mem1[219][9] ), .SE(test_se), 
        .CLK(n1434), .Q(\mem1[219][10] ), .QN(n25894) );
  SDFFX1 \mem1_reg[219][9]  ( .D(n16261), .SI(\mem1[219][8] ), .SE(test_se), 
        .CLK(n1435), .Q(\mem1[219][9] ), .QN(n25895) );
  SDFFX1 \mem1_reg[219][8]  ( .D(n16260), .SI(\mem1[218][15] ), .SE(test_se), 
        .CLK(n1435), .Q(\mem1[219][8] ), .QN(n25896) );
  SDFFX1 \mem1_reg[218][15]  ( .D(n16259), .SI(\mem1[218][14] ), .SE(test_se), 
        .CLK(n1435), .Q(\mem1[218][15] ), .QN(n25897) );
  SDFFX1 \mem1_reg[218][14]  ( .D(n16258), .SI(\mem1[218][13] ), .SE(test_se), 
        .CLK(n1435), .Q(\mem1[218][14] ), .QN(n25898) );
  SDFFX1 \mem1_reg[218][13]  ( .D(n16257), .SI(\mem1[218][12] ), .SE(test_se), 
        .CLK(n1435), .Q(\mem1[218][13] ), .QN(n25899) );
  SDFFX1 \mem1_reg[218][12]  ( .D(n16256), .SI(\mem1[218][11] ), .SE(test_se), 
        .CLK(n1435), .Q(\mem1[218][12] ), .QN(n25900) );
  SDFFX1 \mem1_reg[218][11]  ( .D(n16255), .SI(\mem1[218][10] ), .SE(test_se), 
        .CLK(n1435), .Q(\mem1[218][11] ), .QN(n25901) );
  SDFFX1 \mem1_reg[218][10]  ( .D(n16254), .SI(\mem1[218][9] ), .SE(test_se), 
        .CLK(n1435), .Q(\mem1[218][10] ), .QN(n25902) );
  SDFFX1 \mem1_reg[218][9]  ( .D(n16253), .SI(\mem1[218][8] ), .SE(test_se), 
        .CLK(n1435), .Q(\mem1[218][9] ), .QN(n25903) );
  SDFFX1 \mem1_reg[218][8]  ( .D(n16252), .SI(\mem1[217][15] ), .SE(test_se), 
        .CLK(n1435), .Q(\mem1[218][8] ), .QN(n25904) );
  SDFFX1 \mem1_reg[217][15]  ( .D(n16251), .SI(\mem1[217][14] ), .SE(test_se), 
        .CLK(n1435), .Q(\mem1[217][15] ), .QN(n25905) );
  SDFFX1 \mem1_reg[217][14]  ( .D(n16250), .SI(\mem1[217][13] ), .SE(test_se), 
        .CLK(n1435), .Q(\mem1[217][14] ), .QN(n25906) );
  SDFFX1 \mem1_reg[217][13]  ( .D(n16249), .SI(\mem1[217][12] ), .SE(test_se), 
        .CLK(n1436), .Q(\mem1[217][13] ), .QN(n25907) );
  SDFFX1 \mem1_reg[217][12]  ( .D(n16248), .SI(\mem1[217][11] ), .SE(test_se), 
        .CLK(n1436), .Q(\mem1[217][12] ), .QN(n25908) );
  SDFFX1 \mem1_reg[217][11]  ( .D(n16247), .SI(\mem1[217][10] ), .SE(test_se), 
        .CLK(n1436), .Q(\mem1[217][11] ), .QN(n25909) );
  SDFFX1 \mem1_reg[217][10]  ( .D(n16246), .SI(\mem1[217][9] ), .SE(test_se), 
        .CLK(n1436), .Q(\mem1[217][10] ), .QN(n25910) );
  SDFFX1 \mem1_reg[217][9]  ( .D(n16245), .SI(\mem1[217][8] ), .SE(test_se), 
        .CLK(n1436), .Q(\mem1[217][9] ), .QN(n25911) );
  SDFFX1 \mem1_reg[217][8]  ( .D(n16244), .SI(\mem1[216][15] ), .SE(test_se), 
        .CLK(n1436), .Q(\mem1[217][8] ), .QN(n25912) );
  SDFFX1 \mem1_reg[216][15]  ( .D(n16243), .SI(\mem1[216][14] ), .SE(test_se), 
        .CLK(n1436), .Q(\mem1[216][15] ), .QN(n25913) );
  SDFFX1 \mem1_reg[216][14]  ( .D(n16242), .SI(\mem1[216][13] ), .SE(test_se), 
        .CLK(n1436), .Q(\mem1[216][14] ), .QN(n25914) );
  SDFFX1 \mem1_reg[216][13]  ( .D(n16241), .SI(\mem1[216][12] ), .SE(test_se), 
        .CLK(n1436), .Q(\mem1[216][13] ), .QN(n25915) );
  SDFFX1 \mem1_reg[216][12]  ( .D(n16240), .SI(\mem1[216][11] ), .SE(test_se), 
        .CLK(n1436), .Q(\mem1[216][12] ), .QN(n25916) );
  SDFFX1 \mem1_reg[216][11]  ( .D(n16239), .SI(\mem1[216][10] ), .SE(test_se), 
        .CLK(n1436), .Q(\mem1[216][11] ), .QN(n25917) );
  SDFFX1 \mem1_reg[216][10]  ( .D(n16238), .SI(\mem1[216][9] ), .SE(test_se), 
        .CLK(n1436), .Q(\mem1[216][10] ), .QN(n25918) );
  SDFFX1 \mem1_reg[216][9]  ( .D(n16237), .SI(\mem1[216][8] ), .SE(test_se), 
        .CLK(n1437), .Q(\mem1[216][9] ), .QN(n25919) );
  SDFFX1 \mem1_reg[216][8]  ( .D(n16236), .SI(\mem1[215][15] ), .SE(test_se), 
        .CLK(n1437), .Q(\mem1[216][8] ), .QN(n25920) );
  SDFFX1 \mem1_reg[215][15]  ( .D(n16235), .SI(\mem1[215][14] ), .SE(test_se), 
        .CLK(n1437), .Q(\mem1[215][15] ), .QN(n25921) );
  SDFFX1 \mem1_reg[215][14]  ( .D(n16234), .SI(\mem1[215][13] ), .SE(test_se), 
        .CLK(n1437), .Q(\mem1[215][14] ), .QN(n25922) );
  SDFFX1 \mem1_reg[215][13]  ( .D(n16233), .SI(\mem1[215][12] ), .SE(test_se), 
        .CLK(n1437), .Q(\mem1[215][13] ), .QN(n25923) );
  SDFFX1 \mem1_reg[215][12]  ( .D(n16232), .SI(\mem1[215][11] ), .SE(test_se), 
        .CLK(n1437), .Q(\mem1[215][12] ), .QN(n25924) );
  SDFFX1 \mem1_reg[215][11]  ( .D(n16231), .SI(\mem1[215][10] ), .SE(test_se), 
        .CLK(n1437), .Q(\mem1[215][11] ), .QN(n25925) );
  SDFFX1 \mem1_reg[215][10]  ( .D(n16230), .SI(\mem1[215][9] ), .SE(test_se), 
        .CLK(n1437), .Q(\mem1[215][10] ), .QN(n25926) );
  SDFFX1 \mem1_reg[215][9]  ( .D(n16229), .SI(\mem1[215][8] ), .SE(test_se), 
        .CLK(n1437), .Q(\mem1[215][9] ), .QN(n25927) );
  SDFFX1 \mem1_reg[215][8]  ( .D(n16228), .SI(\mem1[214][15] ), .SE(test_se), 
        .CLK(n1437), .Q(\mem1[215][8] ), .QN(n25928) );
  SDFFX1 \mem1_reg[214][15]  ( .D(n16227), .SI(\mem1[214][14] ), .SE(test_se), 
        .CLK(n1437), .Q(\mem1[214][15] ), .QN(n25929) );
  SDFFX1 \mem1_reg[214][14]  ( .D(n16226), .SI(\mem1[214][13] ), .SE(test_se), 
        .CLK(n1437), .Q(\mem1[214][14] ), .QN(n25930) );
  SDFFX1 \mem1_reg[214][13]  ( .D(n16225), .SI(\mem1[214][12] ), .SE(test_se), 
        .CLK(n1438), .Q(\mem1[214][13] ), .QN(n25931) );
  SDFFX1 \mem1_reg[214][12]  ( .D(n16224), .SI(\mem1[214][11] ), .SE(test_se), 
        .CLK(n1438), .Q(\mem1[214][12] ), .QN(n25932) );
  SDFFX1 \mem1_reg[214][11]  ( .D(n16223), .SI(\mem1[214][10] ), .SE(test_se), 
        .CLK(n1438), .Q(\mem1[214][11] ), .QN(n25933) );
  SDFFX1 \mem1_reg[214][10]  ( .D(n16222), .SI(\mem1[214][9] ), .SE(test_se), 
        .CLK(n1438), .Q(\mem1[214][10] ), .QN(n25934) );
  SDFFX1 \mem1_reg[214][9]  ( .D(n16221), .SI(\mem1[214][8] ), .SE(test_se), 
        .CLK(n1438), .Q(\mem1[214][9] ), .QN(n25935) );
  SDFFX1 \mem1_reg[214][8]  ( .D(n16220), .SI(\mem1[213][15] ), .SE(test_se), 
        .CLK(n1438), .Q(\mem1[214][8] ), .QN(n25936) );
  SDFFX1 \mem1_reg[213][15]  ( .D(n16219), .SI(\mem1[213][14] ), .SE(test_se), 
        .CLK(n1438), .Q(\mem1[213][15] ), .QN(n25937) );
  SDFFX1 \mem1_reg[213][14]  ( .D(n16218), .SI(\mem1[213][13] ), .SE(test_se), 
        .CLK(n1438), .Q(\mem1[213][14] ), .QN(n25938) );
  SDFFX1 \mem1_reg[213][13]  ( .D(n16217), .SI(\mem1[213][12] ), .SE(test_se), 
        .CLK(n1438), .Q(\mem1[213][13] ), .QN(n25939) );
  SDFFX1 \mem1_reg[213][12]  ( .D(n16216), .SI(\mem1[213][11] ), .SE(test_se), 
        .CLK(n1438), .Q(\mem1[213][12] ), .QN(n25940) );
  SDFFX1 \mem1_reg[213][11]  ( .D(n16215), .SI(\mem1[213][10] ), .SE(test_se), 
        .CLK(n1438), .Q(\mem1[213][11] ), .QN(n25941) );
  SDFFX1 \mem1_reg[213][10]  ( .D(n16214), .SI(\mem1[213][9] ), .SE(test_se), 
        .CLK(n1438), .Q(\mem1[213][10] ), .QN(n25942) );
  SDFFX1 \mem1_reg[213][9]  ( .D(n16213), .SI(\mem1[213][8] ), .SE(test_se), 
        .CLK(n1439), .Q(\mem1[213][9] ), .QN(n25943) );
  SDFFX1 \mem1_reg[213][8]  ( .D(n16212), .SI(\mem1[212][15] ), .SE(test_se), 
        .CLK(n1439), .Q(\mem1[213][8] ), .QN(n25944) );
  SDFFX1 \mem1_reg[212][15]  ( .D(n16211), .SI(\mem1[212][14] ), .SE(test_se), 
        .CLK(n1439), .Q(\mem1[212][15] ), .QN(n25945) );
  SDFFX1 \mem1_reg[212][14]  ( .D(n16210), .SI(\mem1[212][13] ), .SE(test_se), 
        .CLK(n1439), .Q(\mem1[212][14] ), .QN(n25946) );
  SDFFX1 \mem1_reg[212][13]  ( .D(n16209), .SI(\mem1[212][12] ), .SE(test_se), 
        .CLK(n1439), .Q(\mem1[212][13] ), .QN(n25947) );
  SDFFX1 \mem1_reg[212][12]  ( .D(n16208), .SI(\mem1[212][11] ), .SE(test_se), 
        .CLK(n1439), .Q(\mem1[212][12] ), .QN(n25948) );
  SDFFX1 \mem1_reg[212][11]  ( .D(n16207), .SI(\mem1[212][10] ), .SE(test_se), 
        .CLK(n1439), .Q(\mem1[212][11] ), .QN(n25949) );
  SDFFX1 \mem1_reg[212][10]  ( .D(n16206), .SI(\mem1[212][9] ), .SE(test_se), 
        .CLK(n1439), .Q(\mem1[212][10] ), .QN(n25950) );
  SDFFX1 \mem1_reg[212][9]  ( .D(n16205), .SI(\mem1[212][8] ), .SE(test_se), 
        .CLK(n1439), .Q(\mem1[212][9] ), .QN(n25951) );
  SDFFX1 \mem1_reg[212][8]  ( .D(n16204), .SI(\mem1[211][15] ), .SE(test_se), 
        .CLK(n1439), .Q(\mem1[212][8] ), .QN(n25952) );
  SDFFX1 \mem1_reg[211][15]  ( .D(n16203), .SI(\mem1[211][14] ), .SE(test_se), 
        .CLK(n1439), .Q(\mem1[211][15] ), .QN(n25953) );
  SDFFX1 \mem1_reg[211][14]  ( .D(n16202), .SI(\mem1[211][13] ), .SE(test_se), 
        .CLK(n1439), .Q(\mem1[211][14] ), .QN(n25954) );
  SDFFX1 \mem1_reg[211][13]  ( .D(n16201), .SI(\mem1[211][12] ), .SE(test_se), 
        .CLK(n1440), .Q(\mem1[211][13] ), .QN(n25955) );
  SDFFX1 \mem1_reg[211][12]  ( .D(n16200), .SI(\mem1[211][11] ), .SE(test_se), 
        .CLK(n1440), .Q(\mem1[211][12] ), .QN(n25956) );
  SDFFX1 \mem1_reg[211][11]  ( .D(n16199), .SI(\mem1[211][10] ), .SE(test_se), 
        .CLK(n1440), .Q(\mem1[211][11] ), .QN(n25957) );
  SDFFX1 \mem1_reg[211][10]  ( .D(n16198), .SI(\mem1[211][9] ), .SE(test_se), 
        .CLK(n1440), .Q(\mem1[211][10] ), .QN(n25958) );
  SDFFX1 \mem1_reg[211][9]  ( .D(n16197), .SI(\mem1[211][8] ), .SE(test_se), 
        .CLK(n1440), .Q(\mem1[211][9] ), .QN(n25959) );
  SDFFX1 \mem1_reg[211][8]  ( .D(n16196), .SI(\mem1[210][15] ), .SE(test_se), 
        .CLK(n1440), .Q(\mem1[211][8] ), .QN(n25960) );
  SDFFX1 \mem1_reg[210][15]  ( .D(n16195), .SI(\mem1[210][14] ), .SE(test_se), 
        .CLK(n1440), .Q(\mem1[210][15] ), .QN(n25961) );
  SDFFX1 \mem1_reg[210][14]  ( .D(n16194), .SI(\mem1[210][13] ), .SE(test_se), 
        .CLK(n1440), .Q(\mem1[210][14] ), .QN(n25962) );
  SDFFX1 \mem1_reg[210][13]  ( .D(n16193), .SI(\mem1[210][12] ), .SE(test_se), 
        .CLK(n1440), .Q(\mem1[210][13] ), .QN(n25963) );
  SDFFX1 \mem1_reg[210][12]  ( .D(n16192), .SI(\mem1[210][11] ), .SE(test_se), 
        .CLK(n1440), .Q(\mem1[210][12] ), .QN(n25964) );
  SDFFX1 \mem1_reg[210][11]  ( .D(n16191), .SI(\mem1[210][10] ), .SE(test_se), 
        .CLK(n1440), .Q(\mem1[210][11] ), .QN(n25965) );
  SDFFX1 \mem1_reg[210][10]  ( .D(n16190), .SI(\mem1[210][9] ), .SE(test_se), 
        .CLK(n1440), .Q(\mem1[210][10] ), .QN(n25966) );
  SDFFX1 \mem1_reg[210][9]  ( .D(n16189), .SI(\mem1[210][8] ), .SE(test_se), 
        .CLK(n1441), .Q(\mem1[210][9] ), .QN(n25967) );
  SDFFX1 \mem1_reg[210][8]  ( .D(n16188), .SI(\mem1[209][15] ), .SE(test_se), 
        .CLK(n1441), .Q(\mem1[210][8] ), .QN(n25968) );
  SDFFX1 \mem1_reg[209][15]  ( .D(n16187), .SI(\mem1[209][14] ), .SE(test_se), 
        .CLK(n1441), .Q(\mem1[209][15] ), .QN(n25969) );
  SDFFX1 \mem1_reg[209][14]  ( .D(n16186), .SI(\mem1[209][13] ), .SE(test_se), 
        .CLK(n1441), .Q(\mem1[209][14] ), .QN(n25970) );
  SDFFX1 \mem1_reg[209][13]  ( .D(n16185), .SI(\mem1[209][12] ), .SE(test_se), 
        .CLK(n1441), .Q(\mem1[209][13] ), .QN(n25971) );
  SDFFX1 \mem1_reg[209][12]  ( .D(n16184), .SI(\mem1[209][11] ), .SE(test_se), 
        .CLK(n1441), .Q(\mem1[209][12] ), .QN(n25972) );
  SDFFX1 \mem1_reg[209][11]  ( .D(n16183), .SI(\mem1[209][10] ), .SE(test_se), 
        .CLK(n1441), .Q(\mem1[209][11] ), .QN(n25973) );
  SDFFX1 \mem1_reg[209][10]  ( .D(n16182), .SI(\mem1[209][9] ), .SE(test_se), 
        .CLK(n1441), .Q(\mem1[209][10] ), .QN(n25974) );
  SDFFX1 \mem1_reg[209][9]  ( .D(n16181), .SI(\mem1[209][8] ), .SE(test_se), 
        .CLK(n1441), .Q(\mem1[209][9] ), .QN(n25975) );
  SDFFX1 \mem1_reg[209][8]  ( .D(n16180), .SI(\mem1[208][15] ), .SE(test_se), 
        .CLK(n1441), .Q(\mem1[209][8] ), .QN(n25976) );
  SDFFX1 \mem1_reg[208][15]  ( .D(n16179), .SI(\mem1[208][14] ), .SE(test_se), 
        .CLK(n1441), .Q(\mem1[208][15] ), .QN(n25977) );
  SDFFX1 \mem1_reg[208][14]  ( .D(n16178), .SI(\mem1[208][13] ), .SE(test_se), 
        .CLK(n1441), .Q(\mem1[208][14] ), .QN(n25978) );
  SDFFX1 \mem1_reg[208][13]  ( .D(n16177), .SI(\mem1[208][12] ), .SE(test_se), 
        .CLK(n1442), .Q(\mem1[208][13] ), .QN(n25979) );
  SDFFX1 \mem1_reg[208][12]  ( .D(n16176), .SI(\mem1[208][11] ), .SE(test_se), 
        .CLK(n1442), .Q(\mem1[208][12] ), .QN(n25980) );
  SDFFX1 \mem1_reg[208][11]  ( .D(n16175), .SI(\mem1[208][10] ), .SE(test_se), 
        .CLK(n1442), .Q(\mem1[208][11] ), .QN(n25981) );
  SDFFX1 \mem1_reg[208][10]  ( .D(n16174), .SI(\mem1[208][9] ), .SE(test_se), 
        .CLK(n1442), .Q(\mem1[208][10] ), .QN(n25982) );
  SDFFX1 \mem1_reg[208][9]  ( .D(n16173), .SI(\mem1[208][8] ), .SE(test_se), 
        .CLK(n1442), .Q(\mem1[208][9] ), .QN(n25983) );
  SDFFX1 \mem1_reg[208][8]  ( .D(n16172), .SI(\mem1[207][15] ), .SE(test_se), 
        .CLK(n1442), .Q(\mem1[208][8] ), .QN(n25984) );
  SDFFX1 \mem1_reg[207][15]  ( .D(n16171), .SI(\mem1[207][14] ), .SE(test_se), 
        .CLK(n1442), .Q(\mem1[207][15] ), .QN(n25985) );
  SDFFX1 \mem1_reg[207][14]  ( .D(n16170), .SI(\mem1[207][13] ), .SE(test_se), 
        .CLK(n1442), .Q(\mem1[207][14] ), .QN(n25986) );
  SDFFX1 \mem1_reg[207][13]  ( .D(n16169), .SI(\mem1[207][12] ), .SE(test_se), 
        .CLK(n1442), .Q(\mem1[207][13] ), .QN(n25987) );
  SDFFX1 \mem1_reg[207][12]  ( .D(n16168), .SI(\mem1[207][11] ), .SE(test_se), 
        .CLK(n1442), .Q(\mem1[207][12] ), .QN(n25988) );
  SDFFX1 \mem1_reg[207][11]  ( .D(n16167), .SI(\mem1[207][10] ), .SE(test_se), 
        .CLK(n1442), .Q(\mem1[207][11] ), .QN(n25989) );
  SDFFX1 \mem1_reg[207][10]  ( .D(n16166), .SI(\mem1[207][9] ), .SE(test_se), 
        .CLK(n1442), .Q(\mem1[207][10] ), .QN(n25990) );
  SDFFX1 \mem1_reg[207][9]  ( .D(n16165), .SI(\mem1[207][8] ), .SE(test_se), 
        .CLK(n1443), .Q(\mem1[207][9] ), .QN(n25991) );
  SDFFX1 \mem1_reg[207][8]  ( .D(n16164), .SI(\mem1[206][15] ), .SE(test_se), 
        .CLK(n1443), .Q(\mem1[207][8] ), .QN(n25992) );
  SDFFX1 \mem1_reg[206][15]  ( .D(n16163), .SI(\mem1[206][14] ), .SE(test_se), 
        .CLK(n1443), .Q(\mem1[206][15] ), .QN(n25993) );
  SDFFX1 \mem1_reg[206][14]  ( .D(n16162), .SI(\mem1[206][13] ), .SE(test_se), 
        .CLK(n1443), .Q(\mem1[206][14] ), .QN(n25994) );
  SDFFX1 \mem1_reg[206][13]  ( .D(n16161), .SI(\mem1[206][12] ), .SE(test_se), 
        .CLK(n1443), .Q(\mem1[206][13] ), .QN(n25995) );
  SDFFX1 \mem1_reg[206][12]  ( .D(n16160), .SI(\mem1[206][11] ), .SE(test_se), 
        .CLK(n1443), .Q(\mem1[206][12] ), .QN(n25996) );
  SDFFX1 \mem1_reg[206][11]  ( .D(n16159), .SI(\mem1[206][10] ), .SE(test_se), 
        .CLK(n1443), .Q(\mem1[206][11] ), .QN(n25997) );
  SDFFX1 \mem1_reg[206][10]  ( .D(n16158), .SI(\mem1[206][9] ), .SE(test_se), 
        .CLK(n1443), .Q(\mem1[206][10] ), .QN(n25998) );
  SDFFX1 \mem1_reg[206][9]  ( .D(n16157), .SI(\mem1[206][8] ), .SE(test_se), 
        .CLK(n1443), .Q(\mem1[206][9] ), .QN(n25999) );
  SDFFX1 \mem1_reg[206][8]  ( .D(n16156), .SI(\mem1[205][15] ), .SE(test_se), 
        .CLK(n1443), .Q(\mem1[206][8] ), .QN(n26000) );
  SDFFX1 \mem1_reg[205][15]  ( .D(n16155), .SI(\mem1[205][14] ), .SE(test_se), 
        .CLK(n1443), .Q(\mem1[205][15] ), .QN(n26001) );
  SDFFX1 \mem1_reg[205][14]  ( .D(n16154), .SI(\mem1[205][13] ), .SE(test_se), 
        .CLK(n1443), .Q(\mem1[205][14] ), .QN(n26002) );
  SDFFX1 \mem1_reg[205][13]  ( .D(n16153), .SI(\mem1[205][12] ), .SE(test_se), 
        .CLK(n1444), .Q(\mem1[205][13] ), .QN(n26003) );
  SDFFX1 \mem1_reg[205][12]  ( .D(n16152), .SI(\mem1[205][11] ), .SE(test_se), 
        .CLK(n1444), .Q(\mem1[205][12] ), .QN(n26004) );
  SDFFX1 \mem1_reg[205][11]  ( .D(n16151), .SI(\mem1[205][10] ), .SE(test_se), 
        .CLK(n1444), .Q(\mem1[205][11] ), .QN(n26005) );
  SDFFX1 \mem1_reg[205][10]  ( .D(n16150), .SI(\mem1[205][9] ), .SE(test_se), 
        .CLK(n1444), .Q(\mem1[205][10] ), .QN(n26006) );
  SDFFX1 \mem1_reg[205][9]  ( .D(n16149), .SI(\mem1[205][8] ), .SE(test_se), 
        .CLK(n1444), .Q(\mem1[205][9] ), .QN(n26007) );
  SDFFX1 \mem1_reg[205][8]  ( .D(n16148), .SI(\mem1[204][15] ), .SE(test_se), 
        .CLK(n1444), .Q(\mem1[205][8] ), .QN(n26008) );
  SDFFX1 \mem1_reg[204][15]  ( .D(n16147), .SI(\mem1[204][14] ), .SE(test_se), 
        .CLK(n1444), .Q(\mem1[204][15] ), .QN(n26009) );
  SDFFX1 \mem1_reg[204][14]  ( .D(n16146), .SI(\mem1[204][13] ), .SE(test_se), 
        .CLK(n1444), .Q(\mem1[204][14] ), .QN(n26010) );
  SDFFX1 \mem1_reg[204][13]  ( .D(n16145), .SI(\mem1[204][12] ), .SE(test_se), 
        .CLK(n1444), .Q(\mem1[204][13] ), .QN(n26011) );
  SDFFX1 \mem1_reg[204][12]  ( .D(n16144), .SI(\mem1[204][11] ), .SE(test_se), 
        .CLK(n1444), .Q(\mem1[204][12] ), .QN(n26012) );
  SDFFX1 \mem1_reg[204][11]  ( .D(n16143), .SI(\mem1[204][10] ), .SE(test_se), 
        .CLK(n1444), .Q(\mem1[204][11] ), .QN(n26013) );
  SDFFX1 \mem1_reg[204][10]  ( .D(n16142), .SI(\mem1[204][9] ), .SE(test_se), 
        .CLK(n1444), .Q(\mem1[204][10] ), .QN(n26014) );
  SDFFX1 \mem1_reg[204][9]  ( .D(n16141), .SI(\mem1[204][8] ), .SE(test_se), 
        .CLK(n1445), .Q(\mem1[204][9] ), .QN(n26015) );
  SDFFX1 \mem1_reg[204][8]  ( .D(n16140), .SI(\mem1[203][15] ), .SE(test_se), 
        .CLK(n1445), .Q(\mem1[204][8] ), .QN(n26016) );
  SDFFX1 \mem1_reg[203][15]  ( .D(n16139), .SI(\mem1[203][14] ), .SE(test_se), 
        .CLK(n1445), .Q(\mem1[203][15] ), .QN(n26017) );
  SDFFX1 \mem1_reg[203][14]  ( .D(n16138), .SI(\mem1[203][13] ), .SE(test_se), 
        .CLK(n1445), .Q(\mem1[203][14] ), .QN(n26018) );
  SDFFX1 \mem1_reg[203][13]  ( .D(n16137), .SI(\mem1[203][12] ), .SE(test_se), 
        .CLK(n1445), .Q(\mem1[203][13] ), .QN(n26019) );
  SDFFX1 \mem1_reg[203][12]  ( .D(n16136), .SI(\mem1[203][11] ), .SE(test_se), 
        .CLK(n1445), .Q(\mem1[203][12] ), .QN(n26020) );
  SDFFX1 \mem1_reg[203][11]  ( .D(n16135), .SI(\mem1[203][10] ), .SE(test_se), 
        .CLK(n1445), .Q(\mem1[203][11] ), .QN(n26021) );
  SDFFX1 \mem1_reg[203][10]  ( .D(n16134), .SI(\mem1[203][9] ), .SE(test_se), 
        .CLK(n1445), .Q(\mem1[203][10] ), .QN(n26022) );
  SDFFX1 \mem1_reg[203][9]  ( .D(n16133), .SI(\mem1[203][8] ), .SE(test_se), 
        .CLK(n1445), .Q(\mem1[203][9] ), .QN(n26023) );
  SDFFX1 \mem1_reg[203][8]  ( .D(n16132), .SI(\mem1[202][15] ), .SE(test_se), 
        .CLK(n1445), .Q(\mem1[203][8] ), .QN(n26024) );
  SDFFX1 \mem1_reg[202][15]  ( .D(n16131), .SI(\mem1[202][14] ), .SE(test_se), 
        .CLK(n1445), .Q(\mem1[202][15] ), .QN(n26025) );
  SDFFX1 \mem1_reg[202][14]  ( .D(n16130), .SI(\mem1[202][13] ), .SE(test_se), 
        .CLK(n1445), .Q(\mem1[202][14] ), .QN(n26026) );
  SDFFX1 \mem1_reg[202][13]  ( .D(n16129), .SI(\mem1[202][12] ), .SE(test_se), 
        .CLK(n1446), .Q(\mem1[202][13] ), .QN(n26027) );
  SDFFX1 \mem1_reg[202][12]  ( .D(n16128), .SI(\mem1[202][11] ), .SE(test_se), 
        .CLK(n1446), .Q(\mem1[202][12] ), .QN(n26028) );
  SDFFX1 \mem1_reg[202][11]  ( .D(n16127), .SI(\mem1[202][10] ), .SE(test_se), 
        .CLK(n1446), .Q(\mem1[202][11] ), .QN(n26029) );
  SDFFX1 \mem1_reg[202][10]  ( .D(n16126), .SI(\mem1[202][9] ), .SE(test_se), 
        .CLK(n1446), .Q(\mem1[202][10] ), .QN(n26030) );
  SDFFX1 \mem1_reg[202][9]  ( .D(n16125), .SI(\mem1[202][8] ), .SE(test_se), 
        .CLK(n1446), .Q(\mem1[202][9] ), .QN(n26031) );
  SDFFX1 \mem1_reg[202][8]  ( .D(n16124), .SI(\mem1[201][15] ), .SE(test_se), 
        .CLK(n1446), .Q(\mem1[202][8] ), .QN(n26032) );
  SDFFX1 \mem1_reg[201][15]  ( .D(n16123), .SI(\mem1[201][14] ), .SE(test_se), 
        .CLK(n1446), .Q(\mem1[201][15] ), .QN(n26033) );
  SDFFX1 \mem1_reg[201][14]  ( .D(n16122), .SI(\mem1[201][13] ), .SE(test_se), 
        .CLK(n1446), .Q(\mem1[201][14] ), .QN(n26034) );
  SDFFX1 \mem1_reg[201][13]  ( .D(n16121), .SI(\mem1[201][12] ), .SE(test_se), 
        .CLK(n1446), .Q(\mem1[201][13] ), .QN(n26035) );
  SDFFX1 \mem1_reg[201][12]  ( .D(n16120), .SI(\mem1[201][11] ), .SE(test_se), 
        .CLK(n1446), .Q(\mem1[201][12] ), .QN(n26036) );
  SDFFX1 \mem1_reg[201][11]  ( .D(n16119), .SI(\mem1[201][10] ), .SE(test_se), 
        .CLK(n1446), .Q(\mem1[201][11] ), .QN(n26037) );
  SDFFX1 \mem1_reg[201][10]  ( .D(n16118), .SI(\mem1[201][9] ), .SE(test_se), 
        .CLK(n1446), .Q(\mem1[201][10] ), .QN(n26038) );
  SDFFX1 \mem1_reg[201][9]  ( .D(n16117), .SI(\mem1[201][8] ), .SE(test_se), 
        .CLK(n1447), .Q(\mem1[201][9] ), .QN(n26039) );
  SDFFX1 \mem1_reg[201][8]  ( .D(n16116), .SI(\mem1[200][15] ), .SE(test_se), 
        .CLK(n1447), .Q(\mem1[201][8] ), .QN(n26040) );
  SDFFX1 \mem1_reg[200][15]  ( .D(n16115), .SI(\mem1[200][14] ), .SE(test_se), 
        .CLK(n1447), .Q(\mem1[200][15] ), .QN(n26041) );
  SDFFX1 \mem1_reg[200][14]  ( .D(n16114), .SI(\mem1[200][13] ), .SE(test_se), 
        .CLK(n1447), .Q(\mem1[200][14] ), .QN(n26042) );
  SDFFX1 \mem1_reg[200][13]  ( .D(n16113), .SI(\mem1[200][12] ), .SE(test_se), 
        .CLK(n1447), .Q(\mem1[200][13] ), .QN(n26043) );
  SDFFX1 \mem1_reg[200][12]  ( .D(n16112), .SI(\mem1[200][11] ), .SE(test_se), 
        .CLK(n1447), .Q(\mem1[200][12] ), .QN(n26044) );
  SDFFX1 \mem1_reg[200][11]  ( .D(n16111), .SI(\mem1[200][10] ), .SE(test_se), 
        .CLK(n1447), .Q(\mem1[200][11] ), .QN(n26045) );
  SDFFX1 \mem1_reg[200][10]  ( .D(n16110), .SI(\mem1[200][9] ), .SE(test_se), 
        .CLK(n1447), .Q(\mem1[200][10] ), .QN(n26046) );
  SDFFX1 \mem1_reg[200][9]  ( .D(n16109), .SI(\mem1[200][8] ), .SE(test_se), 
        .CLK(n1447), .Q(\mem1[200][9] ), .QN(n26047) );
  SDFFX1 \mem1_reg[200][8]  ( .D(n16108), .SI(\mem1[199][15] ), .SE(test_se), 
        .CLK(n1447), .Q(\mem1[200][8] ), .QN(n26048) );
  SDFFX1 \mem1_reg[199][15]  ( .D(n16107), .SI(\mem1[199][14] ), .SE(test_se), 
        .CLK(n1447), .Q(\mem1[199][15] ), .QN(n26049) );
  SDFFX1 \mem1_reg[199][14]  ( .D(n16106), .SI(\mem1[199][13] ), .SE(test_se), 
        .CLK(n1447), .Q(\mem1[199][14] ), .QN(n26050) );
  SDFFX1 \mem1_reg[199][13]  ( .D(n16105), .SI(\mem1[199][12] ), .SE(test_se), 
        .CLK(n1448), .Q(\mem1[199][13] ), .QN(n26051) );
  SDFFX1 \mem1_reg[199][12]  ( .D(n16104), .SI(\mem1[199][11] ), .SE(test_se), 
        .CLK(n1448), .Q(\mem1[199][12] ), .QN(n26052) );
  SDFFX1 \mem1_reg[199][11]  ( .D(n16103), .SI(\mem1[199][10] ), .SE(test_se), 
        .CLK(n1448), .Q(\mem1[199][11] ), .QN(n26053) );
  SDFFX1 \mem1_reg[199][10]  ( .D(n16102), .SI(\mem1[199][9] ), .SE(test_se), 
        .CLK(n1448), .Q(\mem1[199][10] ), .QN(n26054) );
  SDFFX1 \mem1_reg[199][9]  ( .D(n16101), .SI(\mem1[199][8] ), .SE(test_se), 
        .CLK(n1448), .Q(\mem1[199][9] ), .QN(n26055) );
  SDFFX1 \mem1_reg[199][8]  ( .D(n16100), .SI(\mem1[198][15] ), .SE(test_se), 
        .CLK(n1448), .Q(\mem1[199][8] ), .QN(n26056) );
  SDFFX1 \mem1_reg[198][15]  ( .D(n16099), .SI(\mem1[198][14] ), .SE(test_se), 
        .CLK(n1448), .Q(\mem1[198][15] ), .QN(n26057) );
  SDFFX1 \mem1_reg[198][14]  ( .D(n16098), .SI(\mem1[198][13] ), .SE(test_se), 
        .CLK(n1448), .Q(\mem1[198][14] ), .QN(n26058) );
  SDFFX1 \mem1_reg[198][13]  ( .D(n16097), .SI(\mem1[198][12] ), .SE(test_se), 
        .CLK(n1448), .Q(\mem1[198][13] ), .QN(n26059) );
  SDFFX1 \mem1_reg[198][12]  ( .D(n16096), .SI(\mem1[198][11] ), .SE(test_se), 
        .CLK(n1448), .Q(\mem1[198][12] ), .QN(n26060) );
  SDFFX1 \mem1_reg[198][11]  ( .D(n16095), .SI(\mem1[198][10] ), .SE(test_se), 
        .CLK(n1448), .Q(\mem1[198][11] ), .QN(n26061) );
  SDFFX1 \mem1_reg[198][10]  ( .D(n16094), .SI(\mem1[198][9] ), .SE(test_se), 
        .CLK(n1448), .Q(\mem1[198][10] ), .QN(n26062) );
  SDFFX1 \mem1_reg[198][9]  ( .D(n16093), .SI(\mem1[198][8] ), .SE(test_se), 
        .CLK(n1449), .Q(\mem1[198][9] ), .QN(n26063) );
  SDFFX1 \mem1_reg[198][8]  ( .D(n16092), .SI(\mem1[197][15] ), .SE(test_se), 
        .CLK(n1449), .Q(\mem1[198][8] ), .QN(n26064) );
  SDFFX1 \mem1_reg[197][15]  ( .D(n16091), .SI(\mem1[197][14] ), .SE(test_se), 
        .CLK(n1449), .Q(\mem1[197][15] ), .QN(n26065) );
  SDFFX1 \mem1_reg[197][14]  ( .D(n16090), .SI(\mem1[197][13] ), .SE(test_se), 
        .CLK(n1449), .Q(\mem1[197][14] ), .QN(n26066) );
  SDFFX1 \mem1_reg[197][13]  ( .D(n16089), .SI(\mem1[197][12] ), .SE(test_se), 
        .CLK(n1449), .Q(\mem1[197][13] ), .QN(n26067) );
  SDFFX1 \mem1_reg[197][12]  ( .D(n16088), .SI(\mem1[197][11] ), .SE(test_se), 
        .CLK(n1449), .Q(\mem1[197][12] ), .QN(n26068) );
  SDFFX1 \mem1_reg[197][11]  ( .D(n16087), .SI(\mem1[197][10] ), .SE(test_se), 
        .CLK(n1449), .Q(\mem1[197][11] ), .QN(n26069) );
  SDFFX1 \mem1_reg[197][10]  ( .D(n16086), .SI(\mem1[197][9] ), .SE(test_se), 
        .CLK(n1449), .Q(\mem1[197][10] ), .QN(n26070) );
  SDFFX1 \mem1_reg[197][9]  ( .D(n16085), .SI(\mem1[197][8] ), .SE(test_se), 
        .CLK(n1449), .Q(\mem1[197][9] ), .QN(n26071) );
  SDFFX1 \mem1_reg[197][8]  ( .D(n16084), .SI(\mem1[196][15] ), .SE(test_se), 
        .CLK(n1449), .Q(\mem1[197][8] ), .QN(n26072) );
  SDFFX1 \mem1_reg[196][15]  ( .D(n16083), .SI(\mem1[196][14] ), .SE(test_se), 
        .CLK(n1449), .Q(\mem1[196][15] ), .QN(n26073) );
  SDFFX1 \mem1_reg[196][14]  ( .D(n16082), .SI(\mem1[196][13] ), .SE(test_se), 
        .CLK(n1449), .Q(\mem1[196][14] ), .QN(n26074) );
  SDFFX1 \mem1_reg[196][13]  ( .D(n16081), .SI(\mem1[196][12] ), .SE(test_se), 
        .CLK(n1450), .Q(\mem1[196][13] ), .QN(n26075) );
  SDFFX1 \mem1_reg[196][12]  ( .D(n16080), .SI(\mem1[196][11] ), .SE(test_se), 
        .CLK(n1450), .Q(\mem1[196][12] ), .QN(n26076) );
  SDFFX1 \mem1_reg[196][11]  ( .D(n16079), .SI(\mem1[196][10] ), .SE(test_se), 
        .CLK(n1450), .Q(\mem1[196][11] ), .QN(n26077) );
  SDFFX1 \mem1_reg[196][10]  ( .D(n16078), .SI(\mem1[196][9] ), .SE(test_se), 
        .CLK(n1450), .Q(\mem1[196][10] ), .QN(n26078) );
  SDFFX1 \mem1_reg[196][9]  ( .D(n16077), .SI(\mem1[196][8] ), .SE(test_se), 
        .CLK(n1450), .Q(\mem1[196][9] ), .QN(n26079) );
  SDFFX1 \mem1_reg[196][8]  ( .D(n16076), .SI(\mem1[195][15] ), .SE(test_se), 
        .CLK(n1450), .Q(\mem1[196][8] ), .QN(n26080) );
  SDFFX1 \mem1_reg[195][15]  ( .D(n16075), .SI(\mem1[195][14] ), .SE(test_se), 
        .CLK(n1450), .Q(\mem1[195][15] ), .QN(n26081) );
  SDFFX1 \mem1_reg[195][14]  ( .D(n16074), .SI(\mem1[195][13] ), .SE(test_se), 
        .CLK(n1450), .Q(\mem1[195][14] ), .QN(n26082) );
  SDFFX1 \mem1_reg[195][13]  ( .D(n16073), .SI(\mem1[195][12] ), .SE(test_se), 
        .CLK(n1450), .Q(\mem1[195][13] ), .QN(n26083) );
  SDFFX1 \mem1_reg[195][12]  ( .D(n16072), .SI(\mem1[195][11] ), .SE(test_se), 
        .CLK(n1450), .Q(\mem1[195][12] ), .QN(n26084) );
  SDFFX1 \mem1_reg[195][11]  ( .D(n16071), .SI(\mem1[195][10] ), .SE(test_se), 
        .CLK(n1450), .Q(\mem1[195][11] ), .QN(n26085) );
  SDFFX1 \mem1_reg[195][10]  ( .D(n16070), .SI(\mem1[195][9] ), .SE(test_se), 
        .CLK(n1450), .Q(\mem1[195][10] ), .QN(n26086) );
  SDFFX1 \mem1_reg[195][9]  ( .D(n16069), .SI(\mem1[195][8] ), .SE(test_se), 
        .CLK(n1451), .Q(\mem1[195][9] ), .QN(n26087) );
  SDFFX1 \mem1_reg[195][8]  ( .D(n16068), .SI(\mem1[194][15] ), .SE(test_se), 
        .CLK(n1451), .Q(\mem1[195][8] ), .QN(n26088) );
  SDFFX1 \mem1_reg[194][15]  ( .D(n16067), .SI(\mem1[194][14] ), .SE(test_se), 
        .CLK(n1451), .Q(\mem1[194][15] ), .QN(n26089) );
  SDFFX1 \mem1_reg[194][14]  ( .D(n16066), .SI(\mem1[194][13] ), .SE(test_se), 
        .CLK(n1451), .Q(\mem1[194][14] ), .QN(n26090) );
  SDFFX1 \mem1_reg[194][13]  ( .D(n16065), .SI(\mem1[194][12] ), .SE(test_se), 
        .CLK(n1451), .Q(\mem1[194][13] ), .QN(n26091) );
  SDFFX1 \mem1_reg[194][12]  ( .D(n16064), .SI(\mem1[194][11] ), .SE(test_se), 
        .CLK(n1451), .Q(\mem1[194][12] ), .QN(n26092) );
  SDFFX1 \mem1_reg[194][11]  ( .D(n16063), .SI(\mem1[194][10] ), .SE(test_se), 
        .CLK(n1451), .Q(\mem1[194][11] ), .QN(n26093) );
  SDFFX1 \mem1_reg[194][10]  ( .D(n16062), .SI(\mem1[194][9] ), .SE(test_se), 
        .CLK(n1451), .Q(\mem1[194][10] ), .QN(n26094) );
  SDFFX1 \mem1_reg[194][9]  ( .D(n16061), .SI(\mem1[194][8] ), .SE(test_se), 
        .CLK(n1451), .Q(\mem1[194][9] ), .QN(n26095) );
  SDFFX1 \mem1_reg[194][8]  ( .D(n16060), .SI(\mem1[193][15] ), .SE(test_se), 
        .CLK(n1451), .Q(\mem1[194][8] ), .QN(n26096) );
  SDFFX1 \mem1_reg[193][15]  ( .D(n16059), .SI(\mem1[193][14] ), .SE(test_se), 
        .CLK(n1451), .Q(\mem1[193][15] ), .QN(n26097) );
  SDFFX1 \mem1_reg[193][14]  ( .D(n16058), .SI(\mem1[193][13] ), .SE(test_se), 
        .CLK(n1451), .Q(\mem1[193][14] ), .QN(n26098) );
  SDFFX1 \mem1_reg[193][13]  ( .D(n16057), .SI(\mem1[193][12] ), .SE(test_se), 
        .CLK(n1452), .Q(\mem1[193][13] ), .QN(n26099) );
  SDFFX1 \mem1_reg[193][12]  ( .D(n16056), .SI(\mem1[193][11] ), .SE(test_se), 
        .CLK(n1452), .Q(\mem1[193][12] ), .QN(n26100) );
  SDFFX1 \mem1_reg[193][11]  ( .D(n16055), .SI(\mem1[193][10] ), .SE(test_se), 
        .CLK(n1452), .Q(\mem1[193][11] ), .QN(n26101) );
  SDFFX1 \mem1_reg[193][10]  ( .D(n16054), .SI(\mem1[193][9] ), .SE(test_se), 
        .CLK(n1452), .Q(\mem1[193][10] ), .QN(n26102) );
  SDFFX1 \mem1_reg[193][9]  ( .D(n16053), .SI(\mem1[193][8] ), .SE(test_se), 
        .CLK(n1452), .Q(\mem1[193][9] ), .QN(n26103) );
  SDFFX1 \mem1_reg[193][8]  ( .D(n16052), .SI(\mem1[192][15] ), .SE(test_se), 
        .CLK(n1452), .Q(\mem1[193][8] ), .QN(n26104) );
  SDFFX1 \mem1_reg[192][15]  ( .D(n16051), .SI(\mem1[192][14] ), .SE(test_se), 
        .CLK(n1452), .Q(\mem1[192][15] ), .QN(n26105) );
  SDFFX1 \mem1_reg[192][14]  ( .D(n16050), .SI(\mem1[192][13] ), .SE(test_se), 
        .CLK(n1452), .Q(\mem1[192][14] ), .QN(n26106) );
  SDFFX1 \mem1_reg[192][13]  ( .D(n16049), .SI(\mem1[192][12] ), .SE(test_se), 
        .CLK(n1452), .Q(\mem1[192][13] ), .QN(n26107) );
  SDFFX1 \mem1_reg[192][12]  ( .D(n16048), .SI(\mem1[192][11] ), .SE(test_se), 
        .CLK(n1452), .Q(\mem1[192][12] ), .QN(n26108) );
  SDFFX1 \mem1_reg[192][11]  ( .D(n16047), .SI(\mem1[192][10] ), .SE(test_se), 
        .CLK(n1452), .Q(\mem1[192][11] ), .QN(n26109) );
  SDFFX1 \mem1_reg[192][10]  ( .D(n16046), .SI(\mem1[192][9] ), .SE(test_se), 
        .CLK(n1452), .Q(\mem1[192][10] ), .QN(n26110) );
  SDFFX1 \mem1_reg[192][9]  ( .D(n16045), .SI(\mem1[192][8] ), .SE(test_se), 
        .CLK(n1453), .Q(\mem1[192][9] ), .QN(n26111) );
  SDFFX1 \mem1_reg[192][8]  ( .D(n16044), .SI(\mem1[191][15] ), .SE(test_se), 
        .CLK(n1453), .Q(\mem1[192][8] ), .QN(n26112) );
  SDFFX1 \mem1_reg[191][15]  ( .D(n16043), .SI(\mem1[191][14] ), .SE(test_se), 
        .CLK(n1453), .Q(\mem1[191][15] ), .QN(n26113) );
  SDFFX1 \mem1_reg[191][14]  ( .D(n16042), .SI(\mem1[191][13] ), .SE(test_se), 
        .CLK(n1453), .Q(\mem1[191][14] ), .QN(n26114) );
  SDFFX1 \mem1_reg[191][13]  ( .D(n16041), .SI(\mem1[191][12] ), .SE(test_se), 
        .CLK(n1453), .Q(\mem1[191][13] ), .QN(n26115) );
  SDFFX1 \mem1_reg[191][12]  ( .D(n16040), .SI(\mem1[191][11] ), .SE(test_se), 
        .CLK(n1453), .Q(\mem1[191][12] ), .QN(n26116) );
  SDFFX1 \mem1_reg[191][11]  ( .D(n16039), .SI(\mem1[191][10] ), .SE(test_se), 
        .CLK(n1453), .Q(\mem1[191][11] ), .QN(n26117) );
  SDFFX1 \mem1_reg[191][10]  ( .D(n16038), .SI(\mem1[191][9] ), .SE(test_se), 
        .CLK(n1453), .Q(\mem1[191][10] ), .QN(n26118) );
  SDFFX1 \mem1_reg[191][9]  ( .D(n16037), .SI(\mem1[191][8] ), .SE(test_se), 
        .CLK(n1453), .Q(\mem1[191][9] ), .QN(n26119) );
  SDFFX1 \mem1_reg[191][8]  ( .D(n16036), .SI(\mem1[190][15] ), .SE(test_se), 
        .CLK(n1453), .Q(\mem1[191][8] ), .QN(n26120) );
  SDFFX1 \mem1_reg[190][15]  ( .D(n16035), .SI(\mem1[190][14] ), .SE(test_se), 
        .CLK(n1453), .Q(\mem1[190][15] ), .QN(n26121) );
  SDFFX1 \mem1_reg[190][14]  ( .D(n16034), .SI(\mem1[190][13] ), .SE(test_se), 
        .CLK(n1453), .Q(\mem1[190][14] ), .QN(n26122) );
  SDFFX1 \mem1_reg[190][13]  ( .D(n16033), .SI(\mem1[190][12] ), .SE(test_se), 
        .CLK(n1454), .Q(\mem1[190][13] ), .QN(n26123) );
  SDFFX1 \mem1_reg[190][12]  ( .D(n16032), .SI(\mem1[190][11] ), .SE(test_se), 
        .CLK(n1454), .Q(\mem1[190][12] ), .QN(n26124) );
  SDFFX1 \mem1_reg[190][11]  ( .D(n16031), .SI(\mem1[190][10] ), .SE(test_se), 
        .CLK(n1454), .Q(\mem1[190][11] ), .QN(n26125) );
  SDFFX1 \mem1_reg[190][10]  ( .D(n16030), .SI(\mem1[190][9] ), .SE(test_se), 
        .CLK(n1454), .Q(\mem1[190][10] ), .QN(n26126) );
  SDFFX1 \mem1_reg[190][9]  ( .D(n16029), .SI(\mem1[190][8] ), .SE(test_se), 
        .CLK(n1454), .Q(\mem1[190][9] ), .QN(n26127) );
  SDFFX1 \mem1_reg[190][8]  ( .D(n16028), .SI(\mem1[189][15] ), .SE(test_se), 
        .CLK(n1454), .Q(\mem1[190][8] ), .QN(n26128) );
  SDFFX1 \mem1_reg[189][15]  ( .D(n16027), .SI(\mem1[189][14] ), .SE(test_se), 
        .CLK(n1454), .Q(\mem1[189][15] ), .QN(n26129) );
  SDFFX1 \mem1_reg[189][14]  ( .D(n16026), .SI(\mem1[189][13] ), .SE(test_se), 
        .CLK(n1454), .Q(\mem1[189][14] ), .QN(n26130) );
  SDFFX1 \mem1_reg[189][13]  ( .D(n16025), .SI(\mem1[189][12] ), .SE(test_se), 
        .CLK(n1454), .Q(\mem1[189][13] ), .QN(n26131) );
  SDFFX1 \mem1_reg[189][12]  ( .D(n16024), .SI(\mem1[189][11] ), .SE(test_se), 
        .CLK(n1454), .Q(\mem1[189][12] ), .QN(n26132) );
  SDFFX1 \mem1_reg[189][11]  ( .D(n16023), .SI(\mem1[189][10] ), .SE(test_se), 
        .CLK(n1454), .Q(\mem1[189][11] ), .QN(n26133) );
  SDFFX1 \mem1_reg[189][10]  ( .D(n16022), .SI(\mem1[189][9] ), .SE(test_se), 
        .CLK(n1454), .Q(\mem1[189][10] ), .QN(n26134) );
  SDFFX1 \mem1_reg[189][9]  ( .D(n16021), .SI(\mem1[189][8] ), .SE(test_se), 
        .CLK(n1455), .Q(\mem1[189][9] ), .QN(n26135) );
  SDFFX1 \mem1_reg[189][8]  ( .D(n16020), .SI(\mem1[188][15] ), .SE(test_se), 
        .CLK(n1455), .Q(\mem1[189][8] ), .QN(n26136) );
  SDFFX1 \mem1_reg[188][15]  ( .D(n16019), .SI(\mem1[188][14] ), .SE(test_se), 
        .CLK(n1455), .Q(\mem1[188][15] ), .QN(n26137) );
  SDFFX1 \mem1_reg[188][14]  ( .D(n16018), .SI(\mem1[188][13] ), .SE(test_se), 
        .CLK(n1455), .Q(\mem1[188][14] ), .QN(n26138) );
  SDFFX1 \mem1_reg[188][13]  ( .D(n16017), .SI(\mem1[188][12] ), .SE(test_se), 
        .CLK(n1455), .Q(\mem1[188][13] ), .QN(n26139) );
  SDFFX1 \mem1_reg[188][12]  ( .D(n16016), .SI(\mem1[188][11] ), .SE(test_se), 
        .CLK(n1455), .Q(\mem1[188][12] ), .QN(n26140) );
  SDFFX1 \mem1_reg[188][11]  ( .D(n16015), .SI(\mem1[188][10] ), .SE(test_se), 
        .CLK(n1455), .Q(\mem1[188][11] ), .QN(n26141) );
  SDFFX1 \mem1_reg[188][10]  ( .D(n16014), .SI(\mem1[188][9] ), .SE(test_se), 
        .CLK(n1455), .Q(\mem1[188][10] ), .QN(n26142) );
  SDFFX1 \mem1_reg[188][9]  ( .D(n16013), .SI(\mem1[188][8] ), .SE(test_se), 
        .CLK(n1455), .Q(\mem1[188][9] ), .QN(n26143) );
  SDFFX1 \mem1_reg[188][8]  ( .D(n16012), .SI(\mem1[187][15] ), .SE(test_se), 
        .CLK(n1455), .Q(\mem1[188][8] ), .QN(n26144) );
  SDFFX1 \mem1_reg[187][15]  ( .D(n16011), .SI(\mem1[187][14] ), .SE(test_se), 
        .CLK(n1455), .Q(\mem1[187][15] ), .QN(n26145) );
  SDFFX1 \mem1_reg[187][14]  ( .D(n16010), .SI(\mem1[187][13] ), .SE(test_se), 
        .CLK(n1455), .Q(\mem1[187][14] ), .QN(n26146) );
  SDFFX1 \mem1_reg[187][13]  ( .D(n16009), .SI(\mem1[187][12] ), .SE(test_se), 
        .CLK(n1456), .Q(\mem1[187][13] ), .QN(n26147) );
  SDFFX1 \mem1_reg[187][12]  ( .D(n16008), .SI(\mem1[187][11] ), .SE(test_se), 
        .CLK(n1456), .Q(\mem1[187][12] ), .QN(n26148) );
  SDFFX1 \mem1_reg[187][11]  ( .D(n16007), .SI(\mem1[187][10] ), .SE(test_se), 
        .CLK(n1456), .Q(\mem1[187][11] ), .QN(n26149) );
  SDFFX1 \mem1_reg[187][10]  ( .D(n16006), .SI(\mem1[187][9] ), .SE(test_se), 
        .CLK(n1456), .Q(\mem1[187][10] ), .QN(n26150) );
  SDFFX1 \mem1_reg[187][9]  ( .D(n16005), .SI(\mem1[187][8] ), .SE(test_se), 
        .CLK(n1456), .Q(\mem1[187][9] ), .QN(n26151) );
  SDFFX1 \mem1_reg[187][8]  ( .D(n16004), .SI(\mem1[186][15] ), .SE(test_se), 
        .CLK(n1456), .Q(\mem1[187][8] ), .QN(n26152) );
  SDFFX1 \mem1_reg[186][15]  ( .D(n16003), .SI(\mem1[186][14] ), .SE(test_se), 
        .CLK(n1456), .Q(\mem1[186][15] ), .QN(n26153) );
  SDFFX1 \mem1_reg[186][14]  ( .D(n16002), .SI(\mem1[186][13] ), .SE(test_se), 
        .CLK(n1456), .Q(\mem1[186][14] ), .QN(n26154) );
  SDFFX1 \mem1_reg[186][13]  ( .D(n16001), .SI(\mem1[186][12] ), .SE(test_se), 
        .CLK(n1456), .Q(\mem1[186][13] ), .QN(n26155) );
  SDFFX1 \mem1_reg[186][12]  ( .D(n16000), .SI(\mem1[186][11] ), .SE(test_se), 
        .CLK(n1456), .Q(\mem1[186][12] ), .QN(n26156) );
  SDFFX1 \mem1_reg[186][11]  ( .D(n15999), .SI(\mem1[186][10] ), .SE(test_se), 
        .CLK(n1456), .Q(\mem1[186][11] ), .QN(n26157) );
  SDFFX1 \mem1_reg[186][10]  ( .D(n15998), .SI(\mem1[186][9] ), .SE(test_se), 
        .CLK(n1456), .Q(\mem1[186][10] ), .QN(n26158) );
  SDFFX1 \mem1_reg[186][9]  ( .D(n15997), .SI(\mem1[186][8] ), .SE(test_se), 
        .CLK(n1457), .Q(\mem1[186][9] ), .QN(n26159) );
  SDFFX1 \mem1_reg[186][8]  ( .D(n15996), .SI(\mem1[185][15] ), .SE(test_se), 
        .CLK(n1457), .Q(\mem1[186][8] ), .QN(n26160) );
  SDFFX1 \mem1_reg[185][15]  ( .D(n15995), .SI(\mem1[185][14] ), .SE(test_se), 
        .CLK(n1457), .Q(\mem1[185][15] ), .QN(n26161) );
  SDFFX1 \mem1_reg[185][14]  ( .D(n15994), .SI(\mem1[185][13] ), .SE(test_se), 
        .CLK(n1457), .Q(\mem1[185][14] ), .QN(n26162) );
  SDFFX1 \mem1_reg[185][13]  ( .D(n15993), .SI(\mem1[185][12] ), .SE(test_se), 
        .CLK(n1457), .Q(\mem1[185][13] ), .QN(n26163) );
  SDFFX1 \mem1_reg[185][12]  ( .D(n15992), .SI(\mem1[185][11] ), .SE(test_se), 
        .CLK(n1457), .Q(\mem1[185][12] ), .QN(n26164) );
  SDFFX1 \mem1_reg[185][11]  ( .D(n15991), .SI(\mem1[185][10] ), .SE(test_se), 
        .CLK(n1457), .Q(\mem1[185][11] ), .QN(n26165) );
  SDFFX1 \mem1_reg[185][10]  ( .D(n15990), .SI(\mem1[185][9] ), .SE(test_se), 
        .CLK(n1457), .Q(\mem1[185][10] ), .QN(n26166) );
  SDFFX1 \mem1_reg[185][9]  ( .D(n15989), .SI(\mem1[185][8] ), .SE(test_se), 
        .CLK(n1457), .Q(\mem1[185][9] ), .QN(n26167) );
  SDFFX1 \mem1_reg[185][8]  ( .D(n15988), .SI(\mem1[184][15] ), .SE(test_se), 
        .CLK(n1457), .Q(\mem1[185][8] ), .QN(n26168) );
  SDFFX1 \mem1_reg[184][15]  ( .D(n15987), .SI(\mem1[184][14] ), .SE(test_se), 
        .CLK(n1457), .Q(\mem1[184][15] ), .QN(n26169) );
  SDFFX1 \mem1_reg[184][14]  ( .D(n15986), .SI(\mem1[184][13] ), .SE(test_se), 
        .CLK(n1457), .Q(\mem1[184][14] ), .QN(n26170) );
  SDFFX1 \mem1_reg[184][13]  ( .D(n15985), .SI(\mem1[184][12] ), .SE(test_se), 
        .CLK(n1458), .Q(\mem1[184][13] ), .QN(n26171) );
  SDFFX1 \mem1_reg[184][12]  ( .D(n15984), .SI(\mem1[184][11] ), .SE(test_se), 
        .CLK(n1458), .Q(\mem1[184][12] ), .QN(n26172) );
  SDFFX1 \mem1_reg[184][11]  ( .D(n15983), .SI(\mem1[184][10] ), .SE(test_se), 
        .CLK(n1458), .Q(\mem1[184][11] ), .QN(n26173) );
  SDFFX1 \mem1_reg[184][10]  ( .D(n15982), .SI(\mem1[184][9] ), .SE(test_se), 
        .CLK(n1458), .Q(\mem1[184][10] ), .QN(n26174) );
  SDFFX1 \mem1_reg[184][9]  ( .D(n15981), .SI(\mem1[184][8] ), .SE(test_se), 
        .CLK(n1458), .Q(\mem1[184][9] ), .QN(n26175) );
  SDFFX1 \mem1_reg[184][8]  ( .D(n15980), .SI(\mem1[183][15] ), .SE(test_se), 
        .CLK(n1458), .Q(\mem1[184][8] ), .QN(n26176) );
  SDFFX1 \mem1_reg[183][15]  ( .D(n15979), .SI(\mem1[183][14] ), .SE(test_se), 
        .CLK(n1458), .Q(\mem1[183][15] ), .QN(n26177) );
  SDFFX1 \mem1_reg[183][14]  ( .D(n15978), .SI(\mem1[183][13] ), .SE(test_se), 
        .CLK(n1458), .Q(\mem1[183][14] ), .QN(n26178) );
  SDFFX1 \mem1_reg[183][13]  ( .D(n15977), .SI(\mem1[183][12] ), .SE(test_se), 
        .CLK(n1458), .Q(\mem1[183][13] ), .QN(n26179) );
  SDFFX1 \mem1_reg[183][12]  ( .D(n15976), .SI(\mem1[183][11] ), .SE(test_se), 
        .CLK(n1458), .Q(\mem1[183][12] ), .QN(n26180) );
  SDFFX1 \mem1_reg[183][11]  ( .D(n15975), .SI(\mem1[183][10] ), .SE(test_se), 
        .CLK(n1458), .Q(\mem1[183][11] ), .QN(n26181) );
  SDFFX1 \mem1_reg[183][10]  ( .D(n15974), .SI(\mem1[183][9] ), .SE(test_se), 
        .CLK(n1458), .Q(\mem1[183][10] ), .QN(n26182) );
  SDFFX1 \mem1_reg[183][9]  ( .D(n15973), .SI(\mem1[183][8] ), .SE(test_se), 
        .CLK(n1459), .Q(\mem1[183][9] ), .QN(n26183) );
  SDFFX1 \mem1_reg[183][8]  ( .D(n15972), .SI(\mem1[182][15] ), .SE(test_se), 
        .CLK(n1459), .Q(\mem1[183][8] ), .QN(n26184) );
  SDFFX1 \mem1_reg[182][15]  ( .D(n15971), .SI(\mem1[182][14] ), .SE(test_se), 
        .CLK(n1459), .Q(\mem1[182][15] ), .QN(n26185) );
  SDFFX1 \mem1_reg[182][14]  ( .D(n15970), .SI(\mem1[182][13] ), .SE(test_se), 
        .CLK(n1459), .Q(\mem1[182][14] ), .QN(n26186) );
  SDFFX1 \mem1_reg[182][13]  ( .D(n15969), .SI(\mem1[182][12] ), .SE(test_se), 
        .CLK(n1459), .Q(\mem1[182][13] ), .QN(n26187) );
  SDFFX1 \mem1_reg[182][12]  ( .D(n15968), .SI(\mem1[182][11] ), .SE(test_se), 
        .CLK(n1459), .Q(\mem1[182][12] ), .QN(n26188) );
  SDFFX1 \mem1_reg[182][11]  ( .D(n15967), .SI(\mem1[182][10] ), .SE(test_se), 
        .CLK(n1459), .Q(\mem1[182][11] ), .QN(n26189) );
  SDFFX1 \mem1_reg[182][10]  ( .D(n15966), .SI(\mem1[182][9] ), .SE(test_se), 
        .CLK(n1459), .Q(\mem1[182][10] ), .QN(n26190) );
  SDFFX1 \mem1_reg[182][9]  ( .D(n15965), .SI(\mem1[182][8] ), .SE(test_se), 
        .CLK(n1459), .Q(\mem1[182][9] ), .QN(n26191) );
  SDFFX1 \mem1_reg[182][8]  ( .D(n15964), .SI(\mem1[181][15] ), .SE(test_se), 
        .CLK(n1459), .Q(\mem1[182][8] ), .QN(n26192) );
  SDFFX1 \mem1_reg[181][15]  ( .D(n15963), .SI(\mem1[181][14] ), .SE(test_se), 
        .CLK(n1459), .Q(\mem1[181][15] ), .QN(n26193) );
  SDFFX1 \mem1_reg[181][14]  ( .D(n15962), .SI(\mem1[181][13] ), .SE(test_se), 
        .CLK(n1459), .Q(\mem1[181][14] ), .QN(n26194) );
  SDFFX1 \mem1_reg[181][13]  ( .D(n15961), .SI(\mem1[181][12] ), .SE(test_se), 
        .CLK(n1460), .Q(\mem1[181][13] ), .QN(n26195) );
  SDFFX1 \mem1_reg[181][12]  ( .D(n15960), .SI(\mem1[181][11] ), .SE(test_se), 
        .CLK(n1460), .Q(\mem1[181][12] ), .QN(n26196) );
  SDFFX1 \mem1_reg[181][11]  ( .D(n15959), .SI(\mem1[181][10] ), .SE(test_se), 
        .CLK(n1460), .Q(\mem1[181][11] ), .QN(n26197) );
  SDFFX1 \mem1_reg[181][10]  ( .D(n15958), .SI(\mem1[181][9] ), .SE(test_se), 
        .CLK(n1460), .Q(\mem1[181][10] ), .QN(n26198) );
  SDFFX1 \mem1_reg[181][9]  ( .D(n15957), .SI(\mem1[181][8] ), .SE(test_se), 
        .CLK(n1460), .Q(\mem1[181][9] ), .QN(n26199) );
  SDFFX1 \mem1_reg[181][8]  ( .D(n15956), .SI(\mem1[180][15] ), .SE(test_se), 
        .CLK(n1460), .Q(\mem1[181][8] ), .QN(n26200) );
  SDFFX1 \mem1_reg[180][15]  ( .D(n15955), .SI(\mem1[180][14] ), .SE(test_se), 
        .CLK(n1460), .Q(\mem1[180][15] ), .QN(n26201) );
  SDFFX1 \mem1_reg[180][14]  ( .D(n15954), .SI(\mem1[180][13] ), .SE(test_se), 
        .CLK(n1460), .Q(\mem1[180][14] ), .QN(n26202) );
  SDFFX1 \mem1_reg[180][13]  ( .D(n15953), .SI(\mem1[180][12] ), .SE(test_se), 
        .CLK(n1460), .Q(\mem1[180][13] ), .QN(n26203) );
  SDFFX1 \mem1_reg[180][12]  ( .D(n15952), .SI(\mem1[180][11] ), .SE(test_se), 
        .CLK(n1460), .Q(\mem1[180][12] ), .QN(n26204) );
  SDFFX1 \mem1_reg[180][11]  ( .D(n15951), .SI(\mem1[180][10] ), .SE(test_se), 
        .CLK(n1460), .Q(\mem1[180][11] ), .QN(n26205) );
  SDFFX1 \mem1_reg[180][10]  ( .D(n15950), .SI(\mem1[180][9] ), .SE(test_se), 
        .CLK(n1460), .Q(\mem1[180][10] ), .QN(n26206) );
  SDFFX1 \mem1_reg[180][9]  ( .D(n15949), .SI(\mem1[180][8] ), .SE(test_se), 
        .CLK(n1461), .Q(\mem1[180][9] ), .QN(n26207) );
  SDFFX1 \mem1_reg[180][8]  ( .D(n15948), .SI(\mem1[179][15] ), .SE(test_se), 
        .CLK(n1461), .Q(\mem1[180][8] ), .QN(n26208) );
  SDFFX1 \mem1_reg[179][15]  ( .D(n15947), .SI(\mem1[179][14] ), .SE(test_se), 
        .CLK(n1461), .Q(\mem1[179][15] ), .QN(n26209) );
  SDFFX1 \mem1_reg[179][14]  ( .D(n15946), .SI(\mem1[179][13] ), .SE(test_se), 
        .CLK(n1461), .Q(\mem1[179][14] ), .QN(n26210) );
  SDFFX1 \mem1_reg[179][13]  ( .D(n15945), .SI(\mem1[179][12] ), .SE(test_se), 
        .CLK(n1461), .Q(\mem1[179][13] ), .QN(n26211) );
  SDFFX1 \mem1_reg[179][12]  ( .D(n15944), .SI(\mem1[179][11] ), .SE(test_se), 
        .CLK(n1461), .Q(\mem1[179][12] ), .QN(n26212) );
  SDFFX1 \mem1_reg[179][11]  ( .D(n15943), .SI(\mem1[179][10] ), .SE(test_se), 
        .CLK(n1461), .Q(\mem1[179][11] ), .QN(n26213) );
  SDFFX1 \mem1_reg[179][10]  ( .D(n15942), .SI(\mem1[179][9] ), .SE(test_se), 
        .CLK(n1461), .Q(\mem1[179][10] ), .QN(n26214) );
  SDFFX1 \mem1_reg[179][9]  ( .D(n15941), .SI(\mem1[179][8] ), .SE(test_se), 
        .CLK(n1461), .Q(\mem1[179][9] ), .QN(n26215) );
  SDFFX1 \mem1_reg[179][8]  ( .D(n15940), .SI(\mem1[178][15] ), .SE(test_se), 
        .CLK(n1461), .Q(\mem1[179][8] ), .QN(n26216) );
  SDFFX1 \mem1_reg[178][15]  ( .D(n15939), .SI(\mem1[178][14] ), .SE(test_se), 
        .CLK(n1461), .Q(\mem1[178][15] ), .QN(n26217) );
  SDFFX1 \mem1_reg[178][14]  ( .D(n15938), .SI(\mem1[178][13] ), .SE(test_se), 
        .CLK(n1461), .Q(\mem1[178][14] ), .QN(n26218) );
  SDFFX1 \mem1_reg[178][13]  ( .D(n15937), .SI(\mem1[178][12] ), .SE(test_se), 
        .CLK(n1462), .Q(\mem1[178][13] ), .QN(n26219) );
  SDFFX1 \mem1_reg[178][12]  ( .D(n15936), .SI(\mem1[178][11] ), .SE(test_se), 
        .CLK(n1462), .Q(\mem1[178][12] ), .QN(n26220) );
  SDFFX1 \mem1_reg[178][11]  ( .D(n15935), .SI(\mem1[178][10] ), .SE(test_se), 
        .CLK(n1462), .Q(\mem1[178][11] ), .QN(n26221) );
  SDFFX1 \mem1_reg[178][10]  ( .D(n15934), .SI(\mem1[178][9] ), .SE(test_se), 
        .CLK(n1462), .Q(\mem1[178][10] ), .QN(n26222) );
  SDFFX1 \mem1_reg[178][9]  ( .D(n15933), .SI(\mem1[178][8] ), .SE(test_se), 
        .CLK(n1462), .Q(\mem1[178][9] ), .QN(n26223) );
  SDFFX1 \mem1_reg[178][8]  ( .D(n15932), .SI(\mem1[177][15] ), .SE(test_se), 
        .CLK(n1462), .Q(\mem1[178][8] ), .QN(n26224) );
  SDFFX1 \mem1_reg[177][15]  ( .D(n15931), .SI(\mem1[177][14] ), .SE(test_se), 
        .CLK(n1462), .Q(\mem1[177][15] ), .QN(n26225) );
  SDFFX1 \mem1_reg[177][14]  ( .D(n15930), .SI(\mem1[177][13] ), .SE(test_se), 
        .CLK(n1462), .Q(\mem1[177][14] ), .QN(n26226) );
  SDFFX1 \mem1_reg[177][13]  ( .D(n15929), .SI(\mem1[177][12] ), .SE(test_se), 
        .CLK(n1462), .Q(\mem1[177][13] ), .QN(n26227) );
  SDFFX1 \mem1_reg[177][12]  ( .D(n15928), .SI(\mem1[177][11] ), .SE(test_se), 
        .CLK(n1462), .Q(\mem1[177][12] ), .QN(n26228) );
  SDFFX1 \mem1_reg[177][11]  ( .D(n15927), .SI(\mem1[177][10] ), .SE(test_se), 
        .CLK(n1462), .Q(\mem1[177][11] ), .QN(n26229) );
  SDFFX1 \mem1_reg[177][10]  ( .D(n15926), .SI(\mem1[177][9] ), .SE(test_se), 
        .CLK(n1462), .Q(\mem1[177][10] ), .QN(n26230) );
  SDFFX1 \mem1_reg[177][9]  ( .D(n15925), .SI(\mem1[177][8] ), .SE(test_se), 
        .CLK(n1463), .Q(\mem1[177][9] ), .QN(n26231) );
  SDFFX1 \mem1_reg[177][8]  ( .D(n15924), .SI(\mem1[176][15] ), .SE(test_se), 
        .CLK(n1463), .Q(\mem1[177][8] ), .QN(n26232) );
  SDFFX1 \mem1_reg[176][15]  ( .D(n15923), .SI(\mem1[176][14] ), .SE(test_se), 
        .CLK(n1463), .Q(\mem1[176][15] ), .QN(n26233) );
  SDFFX1 \mem1_reg[176][14]  ( .D(n15922), .SI(\mem1[176][13] ), .SE(test_se), 
        .CLK(n1463), .Q(\mem1[176][14] ), .QN(n26234) );
  SDFFX1 \mem1_reg[176][13]  ( .D(n15921), .SI(\mem1[176][12] ), .SE(test_se), 
        .CLK(n1463), .Q(\mem1[176][13] ), .QN(n26235) );
  SDFFX1 \mem1_reg[176][12]  ( .D(n15920), .SI(\mem1[176][11] ), .SE(test_se), 
        .CLK(n1463), .Q(\mem1[176][12] ), .QN(n26236) );
  SDFFX1 \mem1_reg[176][11]  ( .D(n15919), .SI(\mem1[176][10] ), .SE(test_se), 
        .CLK(n1463), .Q(\mem1[176][11] ), .QN(n26237) );
  SDFFX1 \mem1_reg[176][10]  ( .D(n15918), .SI(\mem1[176][9] ), .SE(test_se), 
        .CLK(n1463), .Q(\mem1[176][10] ), .QN(n26238) );
  SDFFX1 \mem1_reg[176][9]  ( .D(n15917), .SI(\mem1[176][8] ), .SE(test_se), 
        .CLK(n1463), .Q(\mem1[176][9] ), .QN(n26239) );
  SDFFX1 \mem1_reg[176][8]  ( .D(n15916), .SI(\mem1[175][15] ), .SE(test_se), 
        .CLK(n1463), .Q(\mem1[176][8] ), .QN(n26240) );
  SDFFX1 \mem1_reg[175][15]  ( .D(n15915), .SI(\mem1[175][14] ), .SE(test_se), 
        .CLK(n1463), .Q(\mem1[175][15] ), .QN(n26241) );
  SDFFX1 \mem1_reg[175][14]  ( .D(n15914), .SI(\mem1[175][13] ), .SE(test_se), 
        .CLK(n1463), .Q(\mem1[175][14] ), .QN(n26242) );
  SDFFX1 \mem1_reg[175][13]  ( .D(n15913), .SI(\mem1[175][12] ), .SE(test_se), 
        .CLK(n1464), .Q(\mem1[175][13] ), .QN(n26243) );
  SDFFX1 \mem1_reg[175][12]  ( .D(n15912), .SI(\mem1[175][11] ), .SE(test_se), 
        .CLK(n1464), .Q(\mem1[175][12] ), .QN(n26244) );
  SDFFX1 \mem1_reg[175][11]  ( .D(n15911), .SI(\mem1[175][10] ), .SE(test_se), 
        .CLK(n1464), .Q(\mem1[175][11] ), .QN(n26245) );
  SDFFX1 \mem1_reg[175][10]  ( .D(n15910), .SI(\mem1[175][9] ), .SE(test_se), 
        .CLK(n1464), .Q(\mem1[175][10] ), .QN(n26246) );
  SDFFX1 \mem1_reg[175][9]  ( .D(n15909), .SI(\mem1[175][8] ), .SE(test_se), 
        .CLK(n1464), .Q(\mem1[175][9] ), .QN(n26247) );
  SDFFX1 \mem1_reg[175][8]  ( .D(n15908), .SI(\mem1[174][15] ), .SE(test_se), 
        .CLK(n1464), .Q(\mem1[175][8] ), .QN(n26248) );
  SDFFX1 \mem1_reg[174][15]  ( .D(n15907), .SI(\mem1[174][14] ), .SE(test_se), 
        .CLK(n1464), .Q(\mem1[174][15] ), .QN(n26249) );
  SDFFX1 \mem1_reg[174][14]  ( .D(n15906), .SI(\mem1[174][13] ), .SE(test_se), 
        .CLK(n1464), .Q(\mem1[174][14] ), .QN(n26250) );
  SDFFX1 \mem1_reg[174][13]  ( .D(n15905), .SI(\mem1[174][12] ), .SE(test_se), 
        .CLK(n1464), .Q(\mem1[174][13] ), .QN(n26251) );
  SDFFX1 \mem1_reg[174][12]  ( .D(n15904), .SI(\mem1[174][11] ), .SE(test_se), 
        .CLK(n1464), .Q(\mem1[174][12] ), .QN(n26252) );
  SDFFX1 \mem1_reg[174][11]  ( .D(n15903), .SI(\mem1[174][10] ), .SE(test_se), 
        .CLK(n1464), .Q(\mem1[174][11] ), .QN(n26253) );
  SDFFX1 \mem1_reg[174][10]  ( .D(n15902), .SI(\mem1[174][9] ), .SE(test_se), 
        .CLK(n1464), .Q(\mem1[174][10] ), .QN(n26254) );
  SDFFX1 \mem1_reg[174][9]  ( .D(n15901), .SI(\mem1[174][8] ), .SE(test_se), 
        .CLK(n1465), .Q(\mem1[174][9] ), .QN(n26255) );
  SDFFX1 \mem1_reg[174][8]  ( .D(n15900), .SI(\mem1[173][15] ), .SE(test_se), 
        .CLK(n1465), .Q(\mem1[174][8] ), .QN(n26256) );
  SDFFX1 \mem1_reg[173][15]  ( .D(n15899), .SI(\mem1[173][14] ), .SE(test_se), 
        .CLK(n1465), .Q(\mem1[173][15] ), .QN(n26257) );
  SDFFX1 \mem1_reg[173][14]  ( .D(n15898), .SI(\mem1[173][13] ), .SE(test_se), 
        .CLK(n1465), .Q(\mem1[173][14] ), .QN(n26258) );
  SDFFX1 \mem1_reg[173][13]  ( .D(n15897), .SI(\mem1[173][12] ), .SE(test_se), 
        .CLK(n1465), .Q(\mem1[173][13] ), .QN(n26259) );
  SDFFX1 \mem1_reg[173][12]  ( .D(n15896), .SI(\mem1[173][11] ), .SE(test_se), 
        .CLK(n1465), .Q(\mem1[173][12] ), .QN(n26260) );
  SDFFX1 \mem1_reg[173][11]  ( .D(n15895), .SI(\mem1[173][10] ), .SE(test_se), 
        .CLK(n1465), .Q(\mem1[173][11] ), .QN(n26261) );
  SDFFX1 \mem1_reg[173][10]  ( .D(n15894), .SI(\mem1[173][9] ), .SE(test_se), 
        .CLK(n1465), .Q(\mem1[173][10] ), .QN(n26262) );
  SDFFX1 \mem1_reg[173][9]  ( .D(n15893), .SI(\mem1[173][8] ), .SE(test_se), 
        .CLK(n1465), .Q(\mem1[173][9] ), .QN(n26263) );
  SDFFX1 \mem1_reg[173][8]  ( .D(n15892), .SI(\mem1[172][15] ), .SE(test_se), 
        .CLK(n1465), .Q(\mem1[173][8] ), .QN(n26264) );
  SDFFX1 \mem1_reg[172][15]  ( .D(n15891), .SI(\mem1[172][14] ), .SE(test_se), 
        .CLK(n1465), .Q(\mem1[172][15] ), .QN(n26265) );
  SDFFX1 \mem1_reg[172][14]  ( .D(n15890), .SI(\mem1[172][13] ), .SE(test_se), 
        .CLK(n1465), .Q(\mem1[172][14] ), .QN(n26266) );
  SDFFX1 \mem1_reg[172][13]  ( .D(n15889), .SI(\mem1[172][12] ), .SE(test_se), 
        .CLK(n1466), .Q(\mem1[172][13] ), .QN(n26267) );
  SDFFX1 \mem1_reg[172][12]  ( .D(n15888), .SI(\mem1[172][11] ), .SE(test_se), 
        .CLK(n1466), .Q(\mem1[172][12] ), .QN(n26268) );
  SDFFX1 \mem1_reg[172][11]  ( .D(n15887), .SI(\mem1[172][10] ), .SE(test_se), 
        .CLK(n1466), .Q(\mem1[172][11] ), .QN(n26269) );
  SDFFX1 \mem1_reg[172][10]  ( .D(n15886), .SI(\mem1[172][9] ), .SE(test_se), 
        .CLK(n1466), .Q(\mem1[172][10] ), .QN(n26270) );
  SDFFX1 \mem1_reg[172][9]  ( .D(n15885), .SI(\mem1[172][8] ), .SE(test_se), 
        .CLK(n1466), .Q(\mem1[172][9] ), .QN(n26271) );
  SDFFX1 \mem1_reg[172][8]  ( .D(n15884), .SI(\mem1[171][15] ), .SE(test_se), 
        .CLK(n1466), .Q(\mem1[172][8] ), .QN(n26272) );
  SDFFX1 \mem1_reg[171][15]  ( .D(n15883), .SI(\mem1[171][14] ), .SE(test_se), 
        .CLK(n1466), .Q(\mem1[171][15] ), .QN(n26273) );
  SDFFX1 \mem1_reg[171][14]  ( .D(n15882), .SI(\mem1[171][13] ), .SE(test_se), 
        .CLK(n1466), .Q(\mem1[171][14] ), .QN(n26274) );
  SDFFX1 \mem1_reg[171][13]  ( .D(n15881), .SI(\mem1[171][12] ), .SE(test_se), 
        .CLK(n1466), .Q(\mem1[171][13] ), .QN(n26275) );
  SDFFX1 \mem1_reg[171][12]  ( .D(n15880), .SI(\mem1[171][11] ), .SE(test_se), 
        .CLK(n1466), .Q(\mem1[171][12] ), .QN(n26276) );
  SDFFX1 \mem1_reg[171][11]  ( .D(n15879), .SI(\mem1[171][10] ), .SE(test_se), 
        .CLK(n1466), .Q(\mem1[171][11] ), .QN(n26277) );
  SDFFX1 \mem1_reg[171][10]  ( .D(n15878), .SI(\mem1[171][9] ), .SE(test_se), 
        .CLK(n1466), .Q(\mem1[171][10] ), .QN(n26278) );
  SDFFX1 \mem1_reg[171][9]  ( .D(n15877), .SI(\mem1[171][8] ), .SE(test_se), 
        .CLK(n1467), .Q(\mem1[171][9] ), .QN(n26279) );
  SDFFX1 \mem1_reg[171][8]  ( .D(n15876), .SI(\mem1[170][15] ), .SE(test_se), 
        .CLK(n1467), .Q(\mem1[171][8] ), .QN(n26280) );
  SDFFX1 \mem1_reg[170][15]  ( .D(n15875), .SI(\mem1[170][14] ), .SE(test_se), 
        .CLK(n1467), .Q(\mem1[170][15] ), .QN(n26281) );
  SDFFX1 \mem1_reg[170][14]  ( .D(n15874), .SI(\mem1[170][13] ), .SE(test_se), 
        .CLK(n1467), .Q(\mem1[170][14] ), .QN(n26282) );
  SDFFX1 \mem1_reg[170][13]  ( .D(n15873), .SI(\mem1[170][12] ), .SE(test_se), 
        .CLK(n1467), .Q(\mem1[170][13] ), .QN(n26283) );
  SDFFX1 \mem1_reg[170][12]  ( .D(n15872), .SI(\mem1[170][11] ), .SE(test_se), 
        .CLK(n1467), .Q(\mem1[170][12] ), .QN(n26284) );
  SDFFX1 \mem1_reg[170][11]  ( .D(n15871), .SI(\mem1[170][10] ), .SE(test_se), 
        .CLK(n1467), .Q(\mem1[170][11] ), .QN(n26285) );
  SDFFX1 \mem1_reg[170][10]  ( .D(n15870), .SI(\mem1[170][9] ), .SE(test_se), 
        .CLK(n1467), .Q(\mem1[170][10] ), .QN(n26286) );
  SDFFX1 \mem1_reg[170][9]  ( .D(n15869), .SI(\mem1[170][8] ), .SE(test_se), 
        .CLK(n1467), .Q(\mem1[170][9] ), .QN(n26287) );
  SDFFX1 \mem1_reg[170][8]  ( .D(n15868), .SI(\mem1[169][15] ), .SE(test_se), 
        .CLK(n1467), .Q(\mem1[170][8] ), .QN(n26288) );
  SDFFX1 \mem1_reg[169][15]  ( .D(n15867), .SI(\mem1[169][14] ), .SE(test_se), 
        .CLK(n1467), .Q(\mem1[169][15] ), .QN(n26289) );
  SDFFX1 \mem1_reg[169][14]  ( .D(n15866), .SI(\mem1[169][13] ), .SE(test_se), 
        .CLK(n1467), .Q(\mem1[169][14] ), .QN(n26290) );
  SDFFX1 \mem1_reg[169][13]  ( .D(n15865), .SI(\mem1[169][12] ), .SE(test_se), 
        .CLK(n1468), .Q(\mem1[169][13] ), .QN(n26291) );
  SDFFX1 \mem1_reg[169][12]  ( .D(n15864), .SI(\mem1[169][11] ), .SE(test_se), 
        .CLK(n1468), .Q(\mem1[169][12] ), .QN(n26292) );
  SDFFX1 \mem1_reg[169][11]  ( .D(n15863), .SI(\mem1[169][10] ), .SE(test_se), 
        .CLK(n1468), .Q(\mem1[169][11] ), .QN(n26293) );
  SDFFX1 \mem1_reg[169][10]  ( .D(n15862), .SI(\mem1[169][9] ), .SE(test_se), 
        .CLK(n1468), .Q(\mem1[169][10] ), .QN(n26294) );
  SDFFX1 \mem1_reg[169][9]  ( .D(n15861), .SI(\mem1[169][8] ), .SE(test_se), 
        .CLK(n1468), .Q(\mem1[169][9] ), .QN(n26295) );
  SDFFX1 \mem1_reg[169][8]  ( .D(n15860), .SI(\mem1[168][15] ), .SE(test_se), 
        .CLK(n1468), .Q(\mem1[169][8] ), .QN(n26296) );
  SDFFX1 \mem1_reg[168][15]  ( .D(n15859), .SI(\mem1[168][14] ), .SE(test_se), 
        .CLK(n1468), .Q(\mem1[168][15] ), .QN(n26297) );
  SDFFX1 \mem1_reg[168][14]  ( .D(n15858), .SI(\mem1[168][13] ), .SE(test_se), 
        .CLK(n1468), .Q(\mem1[168][14] ), .QN(n26298) );
  SDFFX1 \mem1_reg[168][13]  ( .D(n15857), .SI(\mem1[168][12] ), .SE(test_se), 
        .CLK(n1468), .Q(\mem1[168][13] ), .QN(n26299) );
  SDFFX1 \mem1_reg[168][12]  ( .D(n15856), .SI(\mem1[168][11] ), .SE(test_se), 
        .CLK(n1468), .Q(\mem1[168][12] ), .QN(n26300) );
  SDFFX1 \mem1_reg[168][11]  ( .D(n15855), .SI(\mem1[168][10] ), .SE(test_se), 
        .CLK(n1468), .Q(\mem1[168][11] ), .QN(n26301) );
  SDFFX1 \mem1_reg[168][10]  ( .D(n15854), .SI(\mem1[168][9] ), .SE(test_se), 
        .CLK(n1468), .Q(\mem1[168][10] ), .QN(n26302) );
  SDFFX1 \mem1_reg[168][9]  ( .D(n15853), .SI(\mem1[168][8] ), .SE(test_se), 
        .CLK(n1469), .Q(\mem1[168][9] ), .QN(n26303) );
  SDFFX1 \mem1_reg[168][8]  ( .D(n15852), .SI(\mem1[167][15] ), .SE(test_se), 
        .CLK(n1469), .Q(\mem1[168][8] ), .QN(n26304) );
  SDFFX1 \mem1_reg[167][15]  ( .D(n15851), .SI(\mem1[167][14] ), .SE(test_se), 
        .CLK(n1469), .Q(\mem1[167][15] ), .QN(n26305) );
  SDFFX1 \mem1_reg[167][14]  ( .D(n15850), .SI(\mem1[167][13] ), .SE(test_se), 
        .CLK(n1469), .Q(\mem1[167][14] ), .QN(n26306) );
  SDFFX1 \mem1_reg[167][13]  ( .D(n15849), .SI(\mem1[167][12] ), .SE(test_se), 
        .CLK(n1469), .Q(\mem1[167][13] ), .QN(n26307) );
  SDFFX1 \mem1_reg[167][12]  ( .D(n15848), .SI(\mem1[167][11] ), .SE(test_se), 
        .CLK(n1469), .Q(\mem1[167][12] ), .QN(n26308) );
  SDFFX1 \mem1_reg[167][11]  ( .D(n15847), .SI(\mem1[167][10] ), .SE(test_se), 
        .CLK(n1469), .Q(\mem1[167][11] ), .QN(n26309) );
  SDFFX1 \mem1_reg[167][10]  ( .D(n15846), .SI(\mem1[167][9] ), .SE(test_se), 
        .CLK(n1469), .Q(\mem1[167][10] ), .QN(n26310) );
  SDFFX1 \mem1_reg[167][9]  ( .D(n15845), .SI(\mem1[167][8] ), .SE(test_se), 
        .CLK(n1469), .Q(\mem1[167][9] ), .QN(n26311) );
  SDFFX1 \mem1_reg[167][8]  ( .D(n15844), .SI(\mem1[166][15] ), .SE(test_se), 
        .CLK(n1469), .Q(\mem1[167][8] ), .QN(n26312) );
  SDFFX1 \mem1_reg[166][15]  ( .D(n15843), .SI(\mem1[166][14] ), .SE(test_se), 
        .CLK(n1469), .Q(\mem1[166][15] ), .QN(n26313) );
  SDFFX1 \mem1_reg[166][14]  ( .D(n15842), .SI(\mem1[166][13] ), .SE(test_se), 
        .CLK(n1469), .Q(\mem1[166][14] ), .QN(n26314) );
  SDFFX1 \mem1_reg[166][13]  ( .D(n15841), .SI(\mem1[166][12] ), .SE(test_se), 
        .CLK(n1470), .Q(\mem1[166][13] ), .QN(n26315) );
  SDFFX1 \mem1_reg[166][12]  ( .D(n15840), .SI(\mem1[166][11] ), .SE(test_se), 
        .CLK(n1470), .Q(\mem1[166][12] ), .QN(n26316) );
  SDFFX1 \mem1_reg[166][11]  ( .D(n15839), .SI(\mem1[166][10] ), .SE(test_se), 
        .CLK(n1470), .Q(\mem1[166][11] ), .QN(n26317) );
  SDFFX1 \mem1_reg[166][10]  ( .D(n15838), .SI(\mem1[166][9] ), .SE(test_se), 
        .CLK(n1470), .Q(\mem1[166][10] ), .QN(n26318) );
  SDFFX1 \mem1_reg[166][9]  ( .D(n15837), .SI(\mem1[166][8] ), .SE(test_se), 
        .CLK(n1470), .Q(\mem1[166][9] ), .QN(n26319) );
  SDFFX1 \mem1_reg[166][8]  ( .D(n15836), .SI(\mem1[165][15] ), .SE(test_se), 
        .CLK(n1470), .Q(\mem1[166][8] ), .QN(n26320) );
  SDFFX1 \mem1_reg[165][15]  ( .D(n15835), .SI(\mem1[165][14] ), .SE(test_se), 
        .CLK(n1470), .Q(\mem1[165][15] ), .QN(n26321) );
  SDFFX1 \mem1_reg[165][14]  ( .D(n15834), .SI(\mem1[165][13] ), .SE(test_se), 
        .CLK(n1470), .Q(\mem1[165][14] ), .QN(n26322) );
  SDFFX1 \mem1_reg[165][13]  ( .D(n15833), .SI(\mem1[165][12] ), .SE(test_se), 
        .CLK(n1470), .Q(\mem1[165][13] ), .QN(n26323) );
  SDFFX1 \mem1_reg[165][12]  ( .D(n15832), .SI(\mem1[165][11] ), .SE(test_se), 
        .CLK(n1470), .Q(\mem1[165][12] ), .QN(n26324) );
  SDFFX1 \mem1_reg[165][11]  ( .D(n15831), .SI(\mem1[165][10] ), .SE(test_se), 
        .CLK(n1470), .Q(\mem1[165][11] ), .QN(n26325) );
  SDFFX1 \mem1_reg[165][10]  ( .D(n15830), .SI(\mem1[165][9] ), .SE(test_se), 
        .CLK(n1470), .Q(\mem1[165][10] ), .QN(n26326) );
  SDFFX1 \mem1_reg[165][9]  ( .D(n15829), .SI(\mem1[165][8] ), .SE(test_se), 
        .CLK(n1471), .Q(\mem1[165][9] ), .QN(n26327) );
  SDFFX1 \mem1_reg[165][8]  ( .D(n15828), .SI(\mem1[164][15] ), .SE(test_se), 
        .CLK(n1471), .Q(\mem1[165][8] ), .QN(n26328) );
  SDFFX1 \mem1_reg[164][15]  ( .D(n15827), .SI(\mem1[164][14] ), .SE(test_se), 
        .CLK(n1471), .Q(\mem1[164][15] ), .QN(n26329) );
  SDFFX1 \mem1_reg[164][14]  ( .D(n15826), .SI(\mem1[164][13] ), .SE(test_se), 
        .CLK(n1471), .Q(\mem1[164][14] ), .QN(n26330) );
  SDFFX1 \mem1_reg[164][13]  ( .D(n15825), .SI(\mem1[164][12] ), .SE(test_se), 
        .CLK(n1471), .Q(\mem1[164][13] ), .QN(n26331) );
  SDFFX1 \mem1_reg[164][12]  ( .D(n15824), .SI(\mem1[164][11] ), .SE(test_se), 
        .CLK(n1471), .Q(\mem1[164][12] ), .QN(n26332) );
  SDFFX1 \mem1_reg[164][11]  ( .D(n15823), .SI(\mem1[164][10] ), .SE(test_se), 
        .CLK(n1471), .Q(\mem1[164][11] ), .QN(n26333) );
  SDFFX1 \mem1_reg[164][10]  ( .D(n15822), .SI(\mem1[164][9] ), .SE(test_se), 
        .CLK(n1471), .Q(\mem1[164][10] ), .QN(n26334) );
  SDFFX1 \mem1_reg[164][9]  ( .D(n15821), .SI(\mem1[164][8] ), .SE(test_se), 
        .CLK(n1471), .Q(\mem1[164][9] ), .QN(n26335) );
  SDFFX1 \mem1_reg[164][8]  ( .D(n15820), .SI(\mem1[163][15] ), .SE(test_se), 
        .CLK(n1471), .Q(\mem1[164][8] ), .QN(n26336) );
  SDFFX1 \mem1_reg[163][15]  ( .D(n15819), .SI(\mem1[163][14] ), .SE(test_se), 
        .CLK(n1471), .Q(\mem1[163][15] ), .QN(n26337) );
  SDFFX1 \mem1_reg[163][14]  ( .D(n15818), .SI(\mem1[163][13] ), .SE(test_se), 
        .CLK(n1471), .Q(\mem1[163][14] ), .QN(n26338) );
  SDFFX1 \mem1_reg[163][13]  ( .D(n15817), .SI(\mem1[163][12] ), .SE(test_se), 
        .CLK(n1472), .Q(\mem1[163][13] ), .QN(n26339) );
  SDFFX1 \mem1_reg[163][12]  ( .D(n15816), .SI(\mem1[163][11] ), .SE(test_se), 
        .CLK(n1472), .Q(\mem1[163][12] ), .QN(n26340) );
  SDFFX1 \mem1_reg[163][11]  ( .D(n15815), .SI(\mem1[163][10] ), .SE(test_se), 
        .CLK(n1472), .Q(\mem1[163][11] ), .QN(n26341) );
  SDFFX1 \mem1_reg[163][10]  ( .D(n15814), .SI(\mem1[163][9] ), .SE(test_se), 
        .CLK(n1472), .Q(\mem1[163][10] ), .QN(n26342) );
  SDFFX1 \mem1_reg[163][9]  ( .D(n15813), .SI(\mem1[163][8] ), .SE(test_se), 
        .CLK(n1472), .Q(\mem1[163][9] ), .QN(n26343) );
  SDFFX1 \mem1_reg[163][8]  ( .D(n15812), .SI(\mem1[162][15] ), .SE(test_se), 
        .CLK(n1472), .Q(\mem1[163][8] ), .QN(n26344) );
  SDFFX1 \mem1_reg[162][15]  ( .D(n15811), .SI(\mem1[162][14] ), .SE(test_se), 
        .CLK(n1472), .Q(\mem1[162][15] ), .QN(n26345) );
  SDFFX1 \mem1_reg[162][14]  ( .D(n15810), .SI(\mem1[162][13] ), .SE(test_se), 
        .CLK(n1472), .Q(\mem1[162][14] ), .QN(n26346) );
  SDFFX1 \mem1_reg[162][13]  ( .D(n15809), .SI(\mem1[162][12] ), .SE(test_se), 
        .CLK(n1472), .Q(\mem1[162][13] ), .QN(n26347) );
  SDFFX1 \mem1_reg[162][12]  ( .D(n15808), .SI(\mem1[162][11] ), .SE(test_se), 
        .CLK(n1472), .Q(\mem1[162][12] ), .QN(n26348) );
  SDFFX1 \mem1_reg[162][11]  ( .D(n15807), .SI(\mem1[162][10] ), .SE(test_se), 
        .CLK(n1472), .Q(\mem1[162][11] ), .QN(n26349) );
  SDFFX1 \mem1_reg[162][10]  ( .D(n15806), .SI(\mem1[162][9] ), .SE(test_se), 
        .CLK(n1472), .Q(\mem1[162][10] ), .QN(n26350) );
  SDFFX1 \mem1_reg[162][9]  ( .D(n15805), .SI(\mem1[162][8] ), .SE(test_se), 
        .CLK(n1473), .Q(\mem1[162][9] ), .QN(n26351) );
  SDFFX1 \mem1_reg[162][8]  ( .D(n15804), .SI(\mem1[161][15] ), .SE(test_se), 
        .CLK(n1473), .Q(\mem1[162][8] ), .QN(n26352) );
  SDFFX1 \mem1_reg[161][15]  ( .D(n15803), .SI(\mem1[161][14] ), .SE(test_se), 
        .CLK(n1473), .Q(\mem1[161][15] ), .QN(n26353) );
  SDFFX1 \mem1_reg[161][14]  ( .D(n15802), .SI(\mem1[161][13] ), .SE(test_se), 
        .CLK(n1473), .Q(\mem1[161][14] ), .QN(n26354) );
  SDFFX1 \mem1_reg[161][13]  ( .D(n15801), .SI(\mem1[161][12] ), .SE(test_se), 
        .CLK(n1473), .Q(\mem1[161][13] ), .QN(n26355) );
  SDFFX1 \mem1_reg[161][12]  ( .D(n15800), .SI(\mem1[161][11] ), .SE(test_se), 
        .CLK(n1473), .Q(\mem1[161][12] ), .QN(n26356) );
  SDFFX1 \mem1_reg[161][11]  ( .D(n15799), .SI(\mem1[161][10] ), .SE(test_se), 
        .CLK(n1473), .Q(\mem1[161][11] ), .QN(n26357) );
  SDFFX1 \mem1_reg[161][10]  ( .D(n15798), .SI(\mem1[161][9] ), .SE(test_se), 
        .CLK(n1473), .Q(\mem1[161][10] ), .QN(n26358) );
  SDFFX1 \mem1_reg[161][9]  ( .D(n15797), .SI(\mem1[161][8] ), .SE(test_se), 
        .CLK(n1473), .Q(\mem1[161][9] ), .QN(n26359) );
  SDFFX1 \mem1_reg[161][8]  ( .D(n15796), .SI(\mem1[160][15] ), .SE(test_se), 
        .CLK(n1473), .Q(\mem1[161][8] ), .QN(n26360) );
  SDFFX1 \mem1_reg[160][15]  ( .D(n15795), .SI(\mem1[160][14] ), .SE(test_se), 
        .CLK(n1473), .Q(\mem1[160][15] ), .QN(n26361) );
  SDFFX1 \mem1_reg[160][14]  ( .D(n15794), .SI(\mem1[160][13] ), .SE(test_se), 
        .CLK(n1473), .Q(\mem1[160][14] ), .QN(n26362) );
  SDFFX1 \mem1_reg[160][13]  ( .D(n15793), .SI(\mem1[160][12] ), .SE(test_se), 
        .CLK(n1474), .Q(\mem1[160][13] ), .QN(n26363) );
  SDFFX1 \mem1_reg[160][12]  ( .D(n15792), .SI(\mem1[160][11] ), .SE(test_se), 
        .CLK(n1474), .Q(\mem1[160][12] ), .QN(n26364) );
  SDFFX1 \mem1_reg[160][11]  ( .D(n15791), .SI(\mem1[160][10] ), .SE(test_se), 
        .CLK(n1474), .Q(\mem1[160][11] ), .QN(n26365) );
  SDFFX1 \mem1_reg[160][10]  ( .D(n15790), .SI(\mem1[160][9] ), .SE(test_se), 
        .CLK(n1474), .Q(\mem1[160][10] ), .QN(n26366) );
  SDFFX1 \mem1_reg[160][9]  ( .D(n15789), .SI(\mem1[160][8] ), .SE(test_se), 
        .CLK(n1474), .Q(\mem1[160][9] ), .QN(n26367) );
  SDFFX1 \mem1_reg[160][8]  ( .D(n15788), .SI(\mem1[159][15] ), .SE(test_se), 
        .CLK(n1474), .Q(\mem1[160][8] ), .QN(n26368) );
  SDFFX1 \mem1_reg[159][15]  ( .D(n15787), .SI(\mem1[159][14] ), .SE(test_se), 
        .CLK(n1474), .Q(\mem1[159][15] ), .QN(n26369) );
  SDFFX1 \mem1_reg[159][14]  ( .D(n15786), .SI(\mem1[159][13] ), .SE(test_se), 
        .CLK(n1474), .Q(\mem1[159][14] ), .QN(n26370) );
  SDFFX1 \mem1_reg[159][13]  ( .D(n15785), .SI(\mem1[159][12] ), .SE(test_se), 
        .CLK(n1474), .Q(\mem1[159][13] ), .QN(n26371) );
  SDFFX1 \mem1_reg[159][12]  ( .D(n15784), .SI(\mem1[159][11] ), .SE(test_se), 
        .CLK(n1474), .Q(\mem1[159][12] ), .QN(n26372) );
  SDFFX1 \mem1_reg[159][11]  ( .D(n15783), .SI(\mem1[159][10] ), .SE(test_se), 
        .CLK(n1474), .Q(\mem1[159][11] ), .QN(n26373) );
  SDFFX1 \mem1_reg[159][10]  ( .D(n15782), .SI(\mem1[159][9] ), .SE(test_se), 
        .CLK(n1474), .Q(\mem1[159][10] ), .QN(n26374) );
  SDFFX1 \mem1_reg[159][9]  ( .D(n15781), .SI(\mem1[159][8] ), .SE(test_se), 
        .CLK(n1475), .Q(\mem1[159][9] ), .QN(n26375) );
  SDFFX1 \mem1_reg[159][8]  ( .D(n15780), .SI(\mem1[158][15] ), .SE(test_se), 
        .CLK(n1475), .Q(\mem1[159][8] ), .QN(n26376) );
  SDFFX1 \mem1_reg[158][15]  ( .D(n15779), .SI(\mem1[158][14] ), .SE(test_se), 
        .CLK(n1475), .Q(\mem1[158][15] ), .QN(n26377) );
  SDFFX1 \mem1_reg[158][14]  ( .D(n15778), .SI(\mem1[158][13] ), .SE(test_se), 
        .CLK(n1475), .Q(\mem1[158][14] ), .QN(n26378) );
  SDFFX1 \mem1_reg[158][13]  ( .D(n15777), .SI(\mem1[158][12] ), .SE(test_se), 
        .CLK(n1475), .Q(\mem1[158][13] ), .QN(n26379) );
  SDFFX1 \mem1_reg[158][12]  ( .D(n15776), .SI(\mem1[158][11] ), .SE(test_se), 
        .CLK(n1475), .Q(\mem1[158][12] ), .QN(n26380) );
  SDFFX1 \mem1_reg[158][11]  ( .D(n15775), .SI(\mem1[158][10] ), .SE(test_se), 
        .CLK(n1475), .Q(\mem1[158][11] ), .QN(n26381) );
  SDFFX1 \mem1_reg[158][10]  ( .D(n15774), .SI(\mem1[158][9] ), .SE(test_se), 
        .CLK(n1475), .Q(\mem1[158][10] ), .QN(n26382) );
  SDFFX1 \mem1_reg[158][9]  ( .D(n15773), .SI(\mem1[158][8] ), .SE(test_se), 
        .CLK(n1475), .Q(\mem1[158][9] ), .QN(n26383) );
  SDFFX1 \mem1_reg[158][8]  ( .D(n15772), .SI(\mem1[157][15] ), .SE(test_se), 
        .CLK(n1475), .Q(\mem1[158][8] ), .QN(n26384) );
  SDFFX1 \mem1_reg[157][15]  ( .D(n15771), .SI(\mem1[157][14] ), .SE(test_se), 
        .CLK(n1475), .Q(\mem1[157][15] ), .QN(n26385) );
  SDFFX1 \mem1_reg[157][14]  ( .D(n15770), .SI(\mem1[157][13] ), .SE(test_se), 
        .CLK(n1475), .Q(\mem1[157][14] ), .QN(n26386) );
  SDFFX1 \mem1_reg[157][13]  ( .D(n15769), .SI(\mem1[157][12] ), .SE(test_se), 
        .CLK(n1476), .Q(\mem1[157][13] ), .QN(n26387) );
  SDFFX1 \mem1_reg[157][12]  ( .D(n15768), .SI(\mem1[157][11] ), .SE(test_se), 
        .CLK(n1476), .Q(\mem1[157][12] ), .QN(n26388) );
  SDFFX1 \mem1_reg[157][11]  ( .D(n15767), .SI(\mem1[157][10] ), .SE(test_se), 
        .CLK(n1476), .Q(\mem1[157][11] ), .QN(n26389) );
  SDFFX1 \mem1_reg[157][10]  ( .D(n15766), .SI(\mem1[157][9] ), .SE(test_se), 
        .CLK(n1476), .Q(\mem1[157][10] ), .QN(n26390) );
  SDFFX1 \mem1_reg[157][9]  ( .D(n15765), .SI(\mem1[157][8] ), .SE(test_se), 
        .CLK(n1476), .Q(\mem1[157][9] ), .QN(n26391) );
  SDFFX1 \mem1_reg[157][8]  ( .D(n15764), .SI(\mem1[156][15] ), .SE(test_se), 
        .CLK(n1476), .Q(\mem1[157][8] ), .QN(n26392) );
  SDFFX1 \mem1_reg[156][15]  ( .D(n15763), .SI(\mem1[156][14] ), .SE(test_se), 
        .CLK(n1476), .Q(\mem1[156][15] ), .QN(n26393) );
  SDFFX1 \mem1_reg[156][14]  ( .D(n15762), .SI(\mem1[156][13] ), .SE(test_se), 
        .CLK(n1476), .Q(\mem1[156][14] ), .QN(n26394) );
  SDFFX1 \mem1_reg[156][13]  ( .D(n15761), .SI(\mem1[156][12] ), .SE(test_se), 
        .CLK(n1476), .Q(\mem1[156][13] ), .QN(n26395) );
  SDFFX1 \mem1_reg[156][12]  ( .D(n15760), .SI(\mem1[156][11] ), .SE(test_se), 
        .CLK(n1476), .Q(\mem1[156][12] ), .QN(n26396) );
  SDFFX1 \mem1_reg[156][11]  ( .D(n15759), .SI(\mem1[156][10] ), .SE(test_se), 
        .CLK(n1476), .Q(\mem1[156][11] ), .QN(n26397) );
  SDFFX1 \mem1_reg[156][10]  ( .D(n15758), .SI(\mem1[156][9] ), .SE(test_se), 
        .CLK(n1476), .Q(\mem1[156][10] ), .QN(n26398) );
  SDFFX1 \mem1_reg[156][9]  ( .D(n15757), .SI(\mem1[156][8] ), .SE(test_se), 
        .CLK(n1477), .Q(\mem1[156][9] ), .QN(n26399) );
  SDFFX1 \mem1_reg[156][8]  ( .D(n15756), .SI(\mem1[155][15] ), .SE(test_se), 
        .CLK(n1477), .Q(\mem1[156][8] ), .QN(n26400) );
  SDFFX1 \mem1_reg[155][15]  ( .D(n15755), .SI(\mem1[155][14] ), .SE(test_se), 
        .CLK(n1477), .Q(\mem1[155][15] ), .QN(n26401) );
  SDFFX1 \mem1_reg[155][14]  ( .D(n15754), .SI(\mem1[155][13] ), .SE(test_se), 
        .CLK(n1477), .Q(\mem1[155][14] ), .QN(n26402) );
  SDFFX1 \mem1_reg[155][13]  ( .D(n15753), .SI(\mem1[155][12] ), .SE(test_se), 
        .CLK(n1477), .Q(\mem1[155][13] ), .QN(n26403) );
  SDFFX1 \mem1_reg[155][12]  ( .D(n15752), .SI(\mem1[155][11] ), .SE(test_se), 
        .CLK(n1477), .Q(\mem1[155][12] ), .QN(n26404) );
  SDFFX1 \mem1_reg[155][11]  ( .D(n15751), .SI(\mem1[155][10] ), .SE(test_se), 
        .CLK(n1477), .Q(\mem1[155][11] ), .QN(n26405) );
  SDFFX1 \mem1_reg[155][10]  ( .D(n15750), .SI(\mem1[155][9] ), .SE(test_se), 
        .CLK(n1477), .Q(\mem1[155][10] ), .QN(n26406) );
  SDFFX1 \mem1_reg[155][9]  ( .D(n15749), .SI(\mem1[155][8] ), .SE(test_se), 
        .CLK(n1477), .Q(\mem1[155][9] ), .QN(n26407) );
  SDFFX1 \mem1_reg[155][8]  ( .D(n15748), .SI(\mem1[154][15] ), .SE(test_se), 
        .CLK(n1477), .Q(\mem1[155][8] ), .QN(n26408) );
  SDFFX1 \mem1_reg[154][15]  ( .D(n15747), .SI(\mem1[154][14] ), .SE(test_se), 
        .CLK(n1477), .Q(\mem1[154][15] ), .QN(n26409) );
  SDFFX1 \mem1_reg[154][14]  ( .D(n15746), .SI(\mem1[154][13] ), .SE(test_se), 
        .CLK(n1477), .Q(\mem1[154][14] ), .QN(n26410) );
  SDFFX1 \mem1_reg[154][13]  ( .D(n15745), .SI(\mem1[154][12] ), .SE(test_se), 
        .CLK(n1478), .Q(\mem1[154][13] ), .QN(n26411) );
  SDFFX1 \mem1_reg[154][12]  ( .D(n15744), .SI(\mem1[154][11] ), .SE(test_se), 
        .CLK(n1478), .Q(\mem1[154][12] ), .QN(n26412) );
  SDFFX1 \mem1_reg[154][11]  ( .D(n15743), .SI(\mem1[154][10] ), .SE(test_se), 
        .CLK(n1478), .Q(\mem1[154][11] ), .QN(n26413) );
  SDFFX1 \mem1_reg[154][10]  ( .D(n15742), .SI(\mem1[154][9] ), .SE(test_se), 
        .CLK(n1478), .Q(\mem1[154][10] ), .QN(n26414) );
  SDFFX1 \mem1_reg[154][9]  ( .D(n15741), .SI(\mem1[154][8] ), .SE(test_se), 
        .CLK(n1478), .Q(\mem1[154][9] ), .QN(n26415) );
  SDFFX1 \mem1_reg[154][8]  ( .D(n15740), .SI(\mem1[153][15] ), .SE(test_se), 
        .CLK(n1478), .Q(\mem1[154][8] ), .QN(n26416) );
  SDFFX1 \mem1_reg[153][15]  ( .D(n15739), .SI(\mem1[153][14] ), .SE(test_se), 
        .CLK(n1478), .Q(\mem1[153][15] ), .QN(n26417) );
  SDFFX1 \mem1_reg[153][14]  ( .D(n15738), .SI(\mem1[153][13] ), .SE(test_se), 
        .CLK(n1478), .Q(\mem1[153][14] ), .QN(n26418) );
  SDFFX1 \mem1_reg[153][13]  ( .D(n15737), .SI(\mem1[153][12] ), .SE(test_se), 
        .CLK(n1478), .Q(\mem1[153][13] ), .QN(n26419) );
  SDFFX1 \mem1_reg[153][12]  ( .D(n15736), .SI(\mem1[153][11] ), .SE(test_se), 
        .CLK(n1478), .Q(\mem1[153][12] ), .QN(n26420) );
  SDFFX1 \mem1_reg[153][11]  ( .D(n15735), .SI(\mem1[153][10] ), .SE(test_se), 
        .CLK(n1478), .Q(\mem1[153][11] ), .QN(n26421) );
  SDFFX1 \mem1_reg[153][10]  ( .D(n15734), .SI(\mem1[153][9] ), .SE(test_se), 
        .CLK(n1478), .Q(\mem1[153][10] ), .QN(n26422) );
  SDFFX1 \mem1_reg[153][9]  ( .D(n15733), .SI(\mem1[153][8] ), .SE(test_se), 
        .CLK(n1479), .Q(\mem1[153][9] ), .QN(n26423) );
  SDFFX1 \mem1_reg[153][8]  ( .D(n15732), .SI(\mem1[152][15] ), .SE(test_se), 
        .CLK(n1479), .Q(\mem1[153][8] ), .QN(n26424) );
  SDFFX1 \mem1_reg[152][15]  ( .D(n15731), .SI(\mem1[152][14] ), .SE(test_se), 
        .CLK(n1479), .Q(\mem1[152][15] ), .QN(n26425) );
  SDFFX1 \mem1_reg[152][14]  ( .D(n15730), .SI(\mem1[152][13] ), .SE(test_se), 
        .CLK(n1479), .Q(\mem1[152][14] ), .QN(n26426) );
  SDFFX1 \mem1_reg[152][13]  ( .D(n15729), .SI(\mem1[152][12] ), .SE(test_se), 
        .CLK(n1479), .Q(\mem1[152][13] ), .QN(n26427) );
  SDFFX1 \mem1_reg[152][12]  ( .D(n15728), .SI(\mem1[152][11] ), .SE(test_se), 
        .CLK(n1479), .Q(\mem1[152][12] ), .QN(n26428) );
  SDFFX1 \mem1_reg[152][11]  ( .D(n15727), .SI(\mem1[152][10] ), .SE(test_se), 
        .CLK(n1479), .Q(\mem1[152][11] ), .QN(n26429) );
  SDFFX1 \mem1_reg[152][10]  ( .D(n15726), .SI(\mem1[152][9] ), .SE(test_se), 
        .CLK(n1479), .Q(\mem1[152][10] ), .QN(n26430) );
  SDFFX1 \mem1_reg[152][9]  ( .D(n15725), .SI(\mem1[152][8] ), .SE(test_se), 
        .CLK(n1479), .Q(\mem1[152][9] ), .QN(n26431) );
  SDFFX1 \mem1_reg[152][8]  ( .D(n15724), .SI(\mem1[151][15] ), .SE(test_se), 
        .CLK(n1479), .Q(\mem1[152][8] ), .QN(n26432) );
  SDFFX1 \mem1_reg[151][15]  ( .D(n15723), .SI(\mem1[151][14] ), .SE(test_se), 
        .CLK(n1479), .Q(\mem1[151][15] ), .QN(n26433) );
  SDFFX1 \mem1_reg[151][14]  ( .D(n15722), .SI(\mem1[151][13] ), .SE(test_se), 
        .CLK(n1479), .Q(\mem1[151][14] ), .QN(n26434) );
  SDFFX1 \mem1_reg[151][13]  ( .D(n15721), .SI(\mem1[151][12] ), .SE(test_se), 
        .CLK(n1480), .Q(\mem1[151][13] ), .QN(n26435) );
  SDFFX1 \mem1_reg[151][12]  ( .D(n15720), .SI(\mem1[151][11] ), .SE(test_se), 
        .CLK(n1480), .Q(\mem1[151][12] ), .QN(n26436) );
  SDFFX1 \mem1_reg[151][11]  ( .D(n15719), .SI(\mem1[151][10] ), .SE(test_se), 
        .CLK(n1480), .Q(\mem1[151][11] ), .QN(n26437) );
  SDFFX1 \mem1_reg[151][10]  ( .D(n15718), .SI(\mem1[151][9] ), .SE(test_se), 
        .CLK(n1480), .Q(\mem1[151][10] ), .QN(n26438) );
  SDFFX1 \mem1_reg[151][9]  ( .D(n15717), .SI(\mem1[151][8] ), .SE(test_se), 
        .CLK(n1480), .Q(\mem1[151][9] ), .QN(n26439) );
  SDFFX1 \mem1_reg[151][8]  ( .D(n15716), .SI(\mem1[150][15] ), .SE(test_se), 
        .CLK(n1480), .Q(\mem1[151][8] ), .QN(n26440) );
  SDFFX1 \mem1_reg[150][15]  ( .D(n15715), .SI(\mem1[150][14] ), .SE(test_se), 
        .CLK(n1480), .Q(\mem1[150][15] ), .QN(n26441) );
  SDFFX1 \mem1_reg[150][14]  ( .D(n15714), .SI(\mem1[150][13] ), .SE(test_se), 
        .CLK(n1480), .Q(\mem1[150][14] ), .QN(n26442) );
  SDFFX1 \mem1_reg[150][13]  ( .D(n15713), .SI(\mem1[150][12] ), .SE(test_se), 
        .CLK(n1480), .Q(\mem1[150][13] ), .QN(n26443) );
  SDFFX1 \mem1_reg[150][12]  ( .D(n15712), .SI(\mem1[150][11] ), .SE(test_se), 
        .CLK(n1480), .Q(\mem1[150][12] ), .QN(n26444) );
  SDFFX1 \mem1_reg[150][11]  ( .D(n15711), .SI(\mem1[150][10] ), .SE(test_se), 
        .CLK(n1480), .Q(\mem1[150][11] ), .QN(n26445) );
  SDFFX1 \mem1_reg[150][10]  ( .D(n15710), .SI(\mem1[150][9] ), .SE(test_se), 
        .CLK(n1480), .Q(\mem1[150][10] ), .QN(n26446) );
  SDFFX1 \mem1_reg[150][9]  ( .D(n15709), .SI(\mem1[150][8] ), .SE(test_se), 
        .CLK(n1481), .Q(\mem1[150][9] ), .QN(n26447) );
  SDFFX1 \mem1_reg[150][8]  ( .D(n15708), .SI(\mem1[149][15] ), .SE(test_se), 
        .CLK(n1481), .Q(\mem1[150][8] ), .QN(n26448) );
  SDFFX1 \mem1_reg[149][15]  ( .D(n15707), .SI(\mem1[149][14] ), .SE(test_se), 
        .CLK(n1481), .Q(\mem1[149][15] ), .QN(n26449) );
  SDFFX1 \mem1_reg[149][14]  ( .D(n15706), .SI(\mem1[149][13] ), .SE(test_se), 
        .CLK(n1481), .Q(\mem1[149][14] ), .QN(n26450) );
  SDFFX1 \mem1_reg[149][13]  ( .D(n15705), .SI(\mem1[149][12] ), .SE(test_se), 
        .CLK(n1481), .Q(\mem1[149][13] ), .QN(n26451) );
  SDFFX1 \mem1_reg[149][12]  ( .D(n15704), .SI(\mem1[149][11] ), .SE(test_se), 
        .CLK(n1481), .Q(\mem1[149][12] ), .QN(n26452) );
  SDFFX1 \mem1_reg[149][11]  ( .D(n15703), .SI(\mem1[149][10] ), .SE(test_se), 
        .CLK(n1481), .Q(\mem1[149][11] ), .QN(n26453) );
  SDFFX1 \mem1_reg[149][10]  ( .D(n15702), .SI(\mem1[149][9] ), .SE(test_se), 
        .CLK(n1481), .Q(\mem1[149][10] ), .QN(n26454) );
  SDFFX1 \mem1_reg[149][9]  ( .D(n15701), .SI(\mem1[149][8] ), .SE(test_se), 
        .CLK(n1481), .Q(\mem1[149][9] ), .QN(n26455) );
  SDFFX1 \mem1_reg[149][8]  ( .D(n15700), .SI(\mem1[148][15] ), .SE(test_se), 
        .CLK(n1481), .Q(\mem1[149][8] ), .QN(n26456) );
  SDFFX1 \mem1_reg[148][15]  ( .D(n15699), .SI(\mem1[148][14] ), .SE(test_se), 
        .CLK(n1481), .Q(\mem1[148][15] ), .QN(n26457) );
  SDFFX1 \mem1_reg[148][14]  ( .D(n15698), .SI(\mem1[148][13] ), .SE(test_se), 
        .CLK(n1481), .Q(\mem1[148][14] ), .QN(n26458) );
  SDFFX1 \mem1_reg[148][13]  ( .D(n15697), .SI(\mem1[148][12] ), .SE(test_se), 
        .CLK(n1482), .Q(\mem1[148][13] ), .QN(n26459) );
  SDFFX1 \mem1_reg[148][12]  ( .D(n15696), .SI(\mem1[148][11] ), .SE(test_se), 
        .CLK(n1482), .Q(\mem1[148][12] ), .QN(n26460) );
  SDFFX1 \mem1_reg[148][11]  ( .D(n15695), .SI(\mem1[148][10] ), .SE(test_se), 
        .CLK(n1482), .Q(\mem1[148][11] ), .QN(n26461) );
  SDFFX1 \mem1_reg[148][10]  ( .D(n15694), .SI(\mem1[148][9] ), .SE(test_se), 
        .CLK(n1482), .Q(\mem1[148][10] ), .QN(n26462) );
  SDFFX1 \mem1_reg[148][9]  ( .D(n15693), .SI(\mem1[148][8] ), .SE(test_se), 
        .CLK(n1482), .Q(\mem1[148][9] ), .QN(n26463) );
  SDFFX1 \mem1_reg[148][8]  ( .D(n15692), .SI(\mem1[147][15] ), .SE(test_se), 
        .CLK(n1482), .Q(\mem1[148][8] ), .QN(n26464) );
  SDFFX1 \mem1_reg[147][15]  ( .D(n15691), .SI(\mem1[147][14] ), .SE(test_se), 
        .CLK(n1482), .Q(\mem1[147][15] ), .QN(n26465) );
  SDFFX1 \mem1_reg[147][14]  ( .D(n15690), .SI(\mem1[147][13] ), .SE(test_se), 
        .CLK(n1482), .Q(\mem1[147][14] ), .QN(n26466) );
  SDFFX1 \mem1_reg[147][13]  ( .D(n15689), .SI(\mem1[147][12] ), .SE(test_se), 
        .CLK(n1482), .Q(\mem1[147][13] ), .QN(n26467) );
  SDFFX1 \mem1_reg[147][12]  ( .D(n15688), .SI(\mem1[147][11] ), .SE(test_se), 
        .CLK(n1482), .Q(\mem1[147][12] ), .QN(n26468) );
  SDFFX1 \mem1_reg[147][11]  ( .D(n15687), .SI(\mem1[147][10] ), .SE(test_se), 
        .CLK(n1482), .Q(\mem1[147][11] ), .QN(n26469) );
  SDFFX1 \mem1_reg[147][10]  ( .D(n15686), .SI(\mem1[147][9] ), .SE(test_se), 
        .CLK(n1482), .Q(\mem1[147][10] ), .QN(n26470) );
  SDFFX1 \mem1_reg[147][9]  ( .D(n15685), .SI(\mem1[147][8] ), .SE(test_se), 
        .CLK(n1483), .Q(\mem1[147][9] ), .QN(n26471) );
  SDFFX1 \mem1_reg[147][8]  ( .D(n15684), .SI(\mem1[146][15] ), .SE(test_se), 
        .CLK(n1483), .Q(\mem1[147][8] ), .QN(n26472) );
  SDFFX1 \mem1_reg[146][15]  ( .D(n15683), .SI(\mem1[146][14] ), .SE(test_se), 
        .CLK(n1483), .Q(\mem1[146][15] ), .QN(n26473) );
  SDFFX1 \mem1_reg[146][14]  ( .D(n15682), .SI(\mem1[146][13] ), .SE(test_se), 
        .CLK(n1483), .Q(\mem1[146][14] ), .QN(n26474) );
  SDFFX1 \mem1_reg[146][13]  ( .D(n15681), .SI(\mem1[146][12] ), .SE(test_se), 
        .CLK(n1483), .Q(\mem1[146][13] ), .QN(n26475) );
  SDFFX1 \mem1_reg[146][12]  ( .D(n15680), .SI(\mem1[146][11] ), .SE(test_se), 
        .CLK(n1483), .Q(\mem1[146][12] ), .QN(n26476) );
  SDFFX1 \mem1_reg[146][11]  ( .D(n15679), .SI(\mem1[146][10] ), .SE(test_se), 
        .CLK(n1483), .Q(\mem1[146][11] ), .QN(n26477) );
  SDFFX1 \mem1_reg[146][10]  ( .D(n15678), .SI(\mem1[146][9] ), .SE(test_se), 
        .CLK(n1483), .Q(\mem1[146][10] ), .QN(n26478) );
  SDFFX1 \mem1_reg[146][9]  ( .D(n15677), .SI(\mem1[146][8] ), .SE(test_se), 
        .CLK(n1483), .Q(\mem1[146][9] ), .QN(n26479) );
  SDFFX1 \mem1_reg[146][8]  ( .D(n15676), .SI(\mem1[145][15] ), .SE(test_se), 
        .CLK(n1483), .Q(\mem1[146][8] ), .QN(n26480) );
  SDFFX1 \mem1_reg[145][15]  ( .D(n15675), .SI(\mem1[145][14] ), .SE(test_se), 
        .CLK(n1483), .Q(\mem1[145][15] ), .QN(n26481) );
  SDFFX1 \mem1_reg[145][14]  ( .D(n15674), .SI(\mem1[145][13] ), .SE(test_se), 
        .CLK(n1483), .Q(\mem1[145][14] ), .QN(n26482) );
  SDFFX1 \mem1_reg[145][13]  ( .D(n15673), .SI(\mem1[145][12] ), .SE(test_se), 
        .CLK(n1484), .Q(\mem1[145][13] ), .QN(n26483) );
  SDFFX1 \mem1_reg[145][12]  ( .D(n15672), .SI(\mem1[145][11] ), .SE(test_se), 
        .CLK(n1484), .Q(\mem1[145][12] ), .QN(n26484) );
  SDFFX1 \mem1_reg[145][11]  ( .D(n15671), .SI(\mem1[145][10] ), .SE(test_se), 
        .CLK(n1484), .Q(\mem1[145][11] ), .QN(n26485) );
  SDFFX1 \mem1_reg[145][10]  ( .D(n15670), .SI(\mem1[145][9] ), .SE(test_se), 
        .CLK(n1484), .Q(\mem1[145][10] ), .QN(n26486) );
  SDFFX1 \mem1_reg[145][9]  ( .D(n15669), .SI(\mem1[145][8] ), .SE(test_se), 
        .CLK(n1484), .Q(\mem1[145][9] ), .QN(n26487) );
  SDFFX1 \mem1_reg[145][8]  ( .D(n15668), .SI(\mem1[144][15] ), .SE(test_se), 
        .CLK(n1484), .Q(\mem1[145][8] ), .QN(n26488) );
  SDFFX1 \mem1_reg[144][15]  ( .D(n15667), .SI(\mem1[144][14] ), .SE(test_se), 
        .CLK(n1484), .Q(\mem1[144][15] ), .QN(n26489) );
  SDFFX1 \mem1_reg[144][14]  ( .D(n15666), .SI(\mem1[144][13] ), .SE(test_se), 
        .CLK(n1484), .Q(\mem1[144][14] ), .QN(n26490) );
  SDFFX1 \mem1_reg[144][13]  ( .D(n15665), .SI(\mem1[144][12] ), .SE(test_se), 
        .CLK(n1484), .Q(\mem1[144][13] ), .QN(n26491) );
  SDFFX1 \mem1_reg[144][12]  ( .D(n15664), .SI(\mem1[144][11] ), .SE(test_se), 
        .CLK(n1484), .Q(\mem1[144][12] ), .QN(n26492) );
  SDFFX1 \mem1_reg[144][11]  ( .D(n15663), .SI(\mem1[144][10] ), .SE(test_se), 
        .CLK(n1484), .Q(\mem1[144][11] ), .QN(n26493) );
  SDFFX1 \mem1_reg[144][10]  ( .D(n15662), .SI(\mem1[144][9] ), .SE(test_se), 
        .CLK(n1484), .Q(\mem1[144][10] ), .QN(n26494) );
  SDFFX1 \mem1_reg[144][9]  ( .D(n15661), .SI(\mem1[144][8] ), .SE(test_se), 
        .CLK(n1485), .Q(\mem1[144][9] ), .QN(n26495) );
  SDFFX1 \mem1_reg[144][8]  ( .D(n15660), .SI(\mem1[143][15] ), .SE(test_se), 
        .CLK(n1485), .Q(\mem1[144][8] ), .QN(n26496) );
  SDFFX1 \mem1_reg[143][15]  ( .D(n15659), .SI(\mem1[143][14] ), .SE(test_se), 
        .CLK(n1485), .Q(\mem1[143][15] ), .QN(n26497) );
  SDFFX1 \mem1_reg[143][14]  ( .D(n15658), .SI(\mem1[143][13] ), .SE(test_se), 
        .CLK(n1485), .Q(\mem1[143][14] ), .QN(n26498) );
  SDFFX1 \mem1_reg[143][13]  ( .D(n15657), .SI(\mem1[143][12] ), .SE(test_se), 
        .CLK(n1485), .Q(\mem1[143][13] ), .QN(n26499) );
  SDFFX1 \mem1_reg[143][12]  ( .D(n15656), .SI(\mem1[143][11] ), .SE(test_se), 
        .CLK(n1485), .Q(\mem1[143][12] ), .QN(n26500) );
  SDFFX1 \mem1_reg[143][11]  ( .D(n15655), .SI(\mem1[143][10] ), .SE(test_se), 
        .CLK(n1485), .Q(\mem1[143][11] ), .QN(n26501) );
  SDFFX1 \mem1_reg[143][10]  ( .D(n15654), .SI(\mem1[143][9] ), .SE(test_se), 
        .CLK(n1485), .Q(\mem1[143][10] ), .QN(n26502) );
  SDFFX1 \mem1_reg[143][9]  ( .D(n15653), .SI(\mem1[143][8] ), .SE(test_se), 
        .CLK(n1485), .Q(\mem1[143][9] ), .QN(n26503) );
  SDFFX1 \mem1_reg[143][8]  ( .D(n15652), .SI(\mem1[142][15] ), .SE(test_se), 
        .CLK(n1485), .Q(\mem1[143][8] ), .QN(n26504) );
  SDFFX1 \mem1_reg[142][15]  ( .D(n15651), .SI(\mem1[142][14] ), .SE(test_se), 
        .CLK(n1485), .Q(\mem1[142][15] ), .QN(n26505) );
  SDFFX1 \mem1_reg[142][14]  ( .D(n15650), .SI(\mem1[142][13] ), .SE(test_se), 
        .CLK(n1485), .Q(\mem1[142][14] ), .QN(n26506) );
  SDFFX1 \mem1_reg[142][13]  ( .D(n15649), .SI(\mem1[142][12] ), .SE(test_se), 
        .CLK(n1486), .Q(\mem1[142][13] ), .QN(n26507) );
  SDFFX1 \mem1_reg[142][12]  ( .D(n15648), .SI(\mem1[142][11] ), .SE(test_se), 
        .CLK(n1486), .Q(\mem1[142][12] ), .QN(n26508) );
  SDFFX1 \mem1_reg[142][11]  ( .D(n15647), .SI(\mem1[142][10] ), .SE(test_se), 
        .CLK(n1486), .Q(\mem1[142][11] ), .QN(n26509) );
  SDFFX1 \mem1_reg[142][10]  ( .D(n15646), .SI(\mem1[142][9] ), .SE(test_se), 
        .CLK(n1486), .Q(\mem1[142][10] ), .QN(n26510) );
  SDFFX1 \mem1_reg[142][9]  ( .D(n15645), .SI(\mem1[142][8] ), .SE(test_se), 
        .CLK(n1486), .Q(\mem1[142][9] ), .QN(n26511) );
  SDFFX1 \mem1_reg[142][8]  ( .D(n15644), .SI(\mem1[141][15] ), .SE(test_se), 
        .CLK(n1486), .Q(\mem1[142][8] ), .QN(n26512) );
  SDFFX1 \mem1_reg[141][15]  ( .D(n15643), .SI(\mem1[141][14] ), .SE(test_se), 
        .CLK(n1486), .Q(\mem1[141][15] ), .QN(n26513) );
  SDFFX1 \mem1_reg[141][14]  ( .D(n15642), .SI(\mem1[141][13] ), .SE(test_se), 
        .CLK(n1486), .Q(\mem1[141][14] ), .QN(n26514) );
  SDFFX1 \mem1_reg[141][13]  ( .D(n15641), .SI(\mem1[141][12] ), .SE(test_se), 
        .CLK(n1486), .Q(\mem1[141][13] ), .QN(n26515) );
  SDFFX1 \mem1_reg[141][12]  ( .D(n15640), .SI(\mem1[141][11] ), .SE(test_se), 
        .CLK(n1486), .Q(\mem1[141][12] ), .QN(n26516) );
  SDFFX1 \mem1_reg[141][11]  ( .D(n15639), .SI(\mem1[141][10] ), .SE(test_se), 
        .CLK(n1486), .Q(\mem1[141][11] ), .QN(n26517) );
  SDFFX1 \mem1_reg[141][10]  ( .D(n15638), .SI(\mem1[141][9] ), .SE(test_se), 
        .CLK(n1486), .Q(\mem1[141][10] ), .QN(n26518) );
  SDFFX1 \mem1_reg[141][9]  ( .D(n15637), .SI(\mem1[141][8] ), .SE(test_se), 
        .CLK(n1487), .Q(\mem1[141][9] ), .QN(n26519) );
  SDFFX1 \mem1_reg[141][8]  ( .D(n15636), .SI(\mem1[140][15] ), .SE(test_se), 
        .CLK(n1487), .Q(\mem1[141][8] ), .QN(n26520) );
  SDFFX1 \mem1_reg[140][15]  ( .D(n15635), .SI(\mem1[140][14] ), .SE(test_se), 
        .CLK(n1487), .Q(\mem1[140][15] ), .QN(n26521) );
  SDFFX1 \mem1_reg[140][14]  ( .D(n15634), .SI(\mem1[140][13] ), .SE(test_se), 
        .CLK(n1487), .Q(\mem1[140][14] ), .QN(n26522) );
  SDFFX1 \mem1_reg[140][13]  ( .D(n15633), .SI(\mem1[140][12] ), .SE(test_se), 
        .CLK(n1487), .Q(\mem1[140][13] ), .QN(n26523) );
  SDFFX1 \mem1_reg[140][12]  ( .D(n15632), .SI(\mem1[140][11] ), .SE(test_se), 
        .CLK(n1487), .Q(\mem1[140][12] ), .QN(n26524) );
  SDFFX1 \mem1_reg[140][11]  ( .D(n15631), .SI(\mem1[140][10] ), .SE(test_se), 
        .CLK(n1487), .Q(\mem1[140][11] ), .QN(n26525) );
  SDFFX1 \mem1_reg[140][10]  ( .D(n15630), .SI(\mem1[140][9] ), .SE(test_se), 
        .CLK(n1487), .Q(\mem1[140][10] ), .QN(n26526) );
  SDFFX1 \mem1_reg[140][9]  ( .D(n15629), .SI(\mem1[140][8] ), .SE(test_se), 
        .CLK(n1487), .Q(\mem1[140][9] ), .QN(n26527) );
  SDFFX1 \mem1_reg[140][8]  ( .D(n15628), .SI(\mem1[139][15] ), .SE(test_se), 
        .CLK(n1487), .Q(\mem1[140][8] ), .QN(n26528) );
  SDFFX1 \mem1_reg[139][15]  ( .D(n15627), .SI(\mem1[139][14] ), .SE(test_se), 
        .CLK(n1487), .Q(\mem1[139][15] ), .QN(n26529) );
  SDFFX1 \mem1_reg[139][14]  ( .D(n15626), .SI(\mem1[139][13] ), .SE(test_se), 
        .CLK(n1487), .Q(\mem1[139][14] ), .QN(n26530) );
  SDFFX1 \mem1_reg[139][13]  ( .D(n15625), .SI(\mem1[139][12] ), .SE(test_se), 
        .CLK(n1488), .Q(\mem1[139][13] ), .QN(n26531) );
  SDFFX1 \mem1_reg[139][12]  ( .D(n15624), .SI(\mem1[139][11] ), .SE(test_se), 
        .CLK(n1488), .Q(\mem1[139][12] ), .QN(n26532) );
  SDFFX1 \mem1_reg[139][11]  ( .D(n15623), .SI(\mem1[139][10] ), .SE(test_se), 
        .CLK(n1488), .Q(\mem1[139][11] ), .QN(n26533) );
  SDFFX1 \mem1_reg[139][10]  ( .D(n15622), .SI(\mem1[139][9] ), .SE(test_se), 
        .CLK(n1488), .Q(\mem1[139][10] ), .QN(n26534) );
  SDFFX1 \mem1_reg[139][9]  ( .D(n15621), .SI(\mem1[139][8] ), .SE(test_se), 
        .CLK(n1488), .Q(\mem1[139][9] ), .QN(n26535) );
  SDFFX1 \mem1_reg[139][8]  ( .D(n15620), .SI(\mem1[138][15] ), .SE(test_se), 
        .CLK(n1488), .Q(\mem1[139][8] ), .QN(n26536) );
  SDFFX1 \mem1_reg[138][15]  ( .D(n15619), .SI(\mem1[138][14] ), .SE(test_se), 
        .CLK(n1488), .Q(\mem1[138][15] ), .QN(n26537) );
  SDFFX1 \mem1_reg[138][14]  ( .D(n15618), .SI(\mem1[138][13] ), .SE(test_se), 
        .CLK(n1488), .Q(\mem1[138][14] ), .QN(n26538) );
  SDFFX1 \mem1_reg[138][13]  ( .D(n15617), .SI(\mem1[138][12] ), .SE(test_se), 
        .CLK(n1488), .Q(\mem1[138][13] ), .QN(n26539) );
  SDFFX1 \mem1_reg[138][12]  ( .D(n15616), .SI(\mem1[138][11] ), .SE(test_se), 
        .CLK(n1488), .Q(\mem1[138][12] ), .QN(n26540) );
  SDFFX1 \mem1_reg[138][11]  ( .D(n15615), .SI(\mem1[138][10] ), .SE(test_se), 
        .CLK(n1488), .Q(\mem1[138][11] ), .QN(n26541) );
  SDFFX1 \mem1_reg[138][10]  ( .D(n15614), .SI(\mem1[138][9] ), .SE(test_se), 
        .CLK(n1488), .Q(\mem1[138][10] ), .QN(n26542) );
  SDFFX1 \mem1_reg[138][9]  ( .D(n15613), .SI(\mem1[138][8] ), .SE(test_se), 
        .CLK(n1489), .Q(\mem1[138][9] ), .QN(n26543) );
  SDFFX1 \mem1_reg[138][8]  ( .D(n15612), .SI(\mem1[137][15] ), .SE(test_se), 
        .CLK(n1489), .Q(\mem1[138][8] ), .QN(n26544) );
  SDFFX1 \mem1_reg[137][15]  ( .D(n15611), .SI(\mem1[137][14] ), .SE(test_se), 
        .CLK(n1489), .Q(\mem1[137][15] ), .QN(n26545) );
  SDFFX1 \mem1_reg[137][14]  ( .D(n15610), .SI(\mem1[137][13] ), .SE(test_se), 
        .CLK(n1489), .Q(\mem1[137][14] ), .QN(n26546) );
  SDFFX1 \mem1_reg[137][13]  ( .D(n15609), .SI(\mem1[137][12] ), .SE(test_se), 
        .CLK(n1489), .Q(\mem1[137][13] ), .QN(n26547) );
  SDFFX1 \mem1_reg[137][12]  ( .D(n15608), .SI(\mem1[137][11] ), .SE(test_se), 
        .CLK(n1489), .Q(\mem1[137][12] ), .QN(n26548) );
  SDFFX1 \mem1_reg[137][11]  ( .D(n15607), .SI(\mem1[137][10] ), .SE(test_se), 
        .CLK(n1489), .Q(\mem1[137][11] ), .QN(n26549) );
  SDFFX1 \mem1_reg[137][10]  ( .D(n15606), .SI(\mem1[137][9] ), .SE(test_se), 
        .CLK(n1489), .Q(\mem1[137][10] ), .QN(n26550) );
  SDFFX1 \mem1_reg[137][9]  ( .D(n15605), .SI(\mem1[137][8] ), .SE(test_se), 
        .CLK(n1489), .Q(\mem1[137][9] ), .QN(n26551) );
  SDFFX1 \mem1_reg[137][8]  ( .D(n15604), .SI(\mem1[136][15] ), .SE(test_se), 
        .CLK(n1489), .Q(\mem1[137][8] ), .QN(n26552) );
  SDFFX1 \mem1_reg[136][15]  ( .D(n15603), .SI(\mem1[136][14] ), .SE(test_se), 
        .CLK(n1489), .Q(\mem1[136][15] ), .QN(n26553) );
  SDFFX1 \mem1_reg[136][14]  ( .D(n15602), .SI(\mem1[136][13] ), .SE(test_se), 
        .CLK(n1489), .Q(\mem1[136][14] ), .QN(n26554) );
  SDFFX1 \mem1_reg[136][13]  ( .D(n15601), .SI(\mem1[136][12] ), .SE(test_se), 
        .CLK(n1490), .Q(\mem1[136][13] ), .QN(n26555) );
  SDFFX1 \mem1_reg[136][12]  ( .D(n15600), .SI(\mem1[136][11] ), .SE(test_se), 
        .CLK(n1490), .Q(\mem1[136][12] ), .QN(n26556) );
  SDFFX1 \mem1_reg[136][11]  ( .D(n15599), .SI(\mem1[136][10] ), .SE(test_se), 
        .CLK(n1490), .Q(\mem1[136][11] ), .QN(n26557) );
  SDFFX1 \mem1_reg[136][10]  ( .D(n15598), .SI(\mem1[136][9] ), .SE(test_se), 
        .CLK(n1490), .Q(\mem1[136][10] ), .QN(n26558) );
  SDFFX1 \mem1_reg[136][9]  ( .D(n15597), .SI(\mem1[136][8] ), .SE(test_se), 
        .CLK(n1490), .Q(\mem1[136][9] ), .QN(n26559) );
  SDFFX1 \mem1_reg[136][8]  ( .D(n15596), .SI(\mem1[135][15] ), .SE(test_se), 
        .CLK(n1490), .Q(\mem1[136][8] ), .QN(n26560) );
  SDFFX1 \mem1_reg[135][15]  ( .D(n15595), .SI(\mem1[135][14] ), .SE(test_se), 
        .CLK(n1490), .Q(\mem1[135][15] ), .QN(n26561) );
  SDFFX1 \mem1_reg[135][14]  ( .D(n15594), .SI(\mem1[135][13] ), .SE(test_se), 
        .CLK(n1490), .Q(\mem1[135][14] ), .QN(n26562) );
  SDFFX1 \mem1_reg[135][13]  ( .D(n15593), .SI(\mem1[135][12] ), .SE(test_se), 
        .CLK(n1490), .Q(\mem1[135][13] ), .QN(n26563) );
  SDFFX1 \mem1_reg[135][12]  ( .D(n15592), .SI(\mem1[135][11] ), .SE(test_se), 
        .CLK(n1490), .Q(\mem1[135][12] ), .QN(n26564) );
  SDFFX1 \mem1_reg[135][11]  ( .D(n15591), .SI(\mem1[135][10] ), .SE(test_se), 
        .CLK(n1490), .Q(\mem1[135][11] ), .QN(n26565) );
  SDFFX1 \mem1_reg[135][10]  ( .D(n15590), .SI(\mem1[135][9] ), .SE(test_se), 
        .CLK(n1490), .Q(\mem1[135][10] ), .QN(n26566) );
  SDFFX1 \mem1_reg[135][9]  ( .D(n15589), .SI(\mem1[135][8] ), .SE(test_se), 
        .CLK(n1491), .Q(\mem1[135][9] ), .QN(n26567) );
  SDFFX1 \mem1_reg[135][8]  ( .D(n15588), .SI(\mem1[134][15] ), .SE(test_se), 
        .CLK(n1491), .Q(\mem1[135][8] ), .QN(n26568) );
  SDFFX1 \mem1_reg[134][15]  ( .D(n15587), .SI(\mem1[134][14] ), .SE(test_se), 
        .CLK(n1491), .Q(\mem1[134][15] ), .QN(n26569) );
  SDFFX1 \mem1_reg[134][14]  ( .D(n15586), .SI(\mem1[134][13] ), .SE(test_se), 
        .CLK(n1491), .Q(\mem1[134][14] ), .QN(n26570) );
  SDFFX1 \mem1_reg[134][13]  ( .D(n15585), .SI(\mem1[134][12] ), .SE(test_se), 
        .CLK(n1491), .Q(\mem1[134][13] ), .QN(n26571) );
  SDFFX1 \mem1_reg[134][12]  ( .D(n15584), .SI(\mem1[134][11] ), .SE(test_se), 
        .CLK(n1491), .Q(\mem1[134][12] ), .QN(n26572) );
  SDFFX1 \mem1_reg[134][11]  ( .D(n15583), .SI(\mem1[134][10] ), .SE(test_se), 
        .CLK(n1491), .Q(\mem1[134][11] ), .QN(n26573) );
  SDFFX1 \mem1_reg[134][10]  ( .D(n15582), .SI(\mem1[134][9] ), .SE(test_se), 
        .CLK(n1491), .Q(\mem1[134][10] ), .QN(n26574) );
  SDFFX1 \mem1_reg[134][9]  ( .D(n15581), .SI(\mem1[134][8] ), .SE(test_se), 
        .CLK(n1491), .Q(\mem1[134][9] ), .QN(n26575) );
  SDFFX1 \mem1_reg[134][8]  ( .D(n15580), .SI(\mem1[133][15] ), .SE(test_se), 
        .CLK(n1491), .Q(\mem1[134][8] ), .QN(n26576) );
  SDFFX1 \mem1_reg[133][15]  ( .D(n15579), .SI(\mem1[133][14] ), .SE(test_se), 
        .CLK(n1491), .Q(\mem1[133][15] ), .QN(n26577) );
  SDFFX1 \mem1_reg[133][14]  ( .D(n15578), .SI(\mem1[133][13] ), .SE(test_se), 
        .CLK(n1491), .Q(\mem1[133][14] ), .QN(n26578) );
  SDFFX1 \mem1_reg[133][13]  ( .D(n15577), .SI(\mem1[133][12] ), .SE(test_se), 
        .CLK(n1492), .Q(\mem1[133][13] ), .QN(n26579) );
  SDFFX1 \mem1_reg[133][12]  ( .D(n15576), .SI(\mem1[133][11] ), .SE(test_se), 
        .CLK(n1492), .Q(\mem1[133][12] ), .QN(n26580) );
  SDFFX1 \mem1_reg[133][11]  ( .D(n15575), .SI(\mem1[133][10] ), .SE(test_se), 
        .CLK(n1492), .Q(\mem1[133][11] ), .QN(n26581) );
  SDFFX1 \mem1_reg[133][10]  ( .D(n15574), .SI(\mem1[133][9] ), .SE(test_se), 
        .CLK(n1492), .Q(\mem1[133][10] ), .QN(n26582) );
  SDFFX1 \mem1_reg[133][9]  ( .D(n15573), .SI(\mem1[133][8] ), .SE(test_se), 
        .CLK(n1492), .Q(\mem1[133][9] ), .QN(n26583) );
  SDFFX1 \mem1_reg[133][8]  ( .D(n15572), .SI(\mem1[132][15] ), .SE(test_se), 
        .CLK(n1492), .Q(\mem1[133][8] ), .QN(n26584) );
  SDFFX1 \mem1_reg[132][15]  ( .D(n15571), .SI(\mem1[132][14] ), .SE(test_se), 
        .CLK(n1492), .Q(\mem1[132][15] ), .QN(n26585) );
  SDFFX1 \mem1_reg[132][14]  ( .D(n15570), .SI(\mem1[132][13] ), .SE(test_se), 
        .CLK(n1492), .Q(\mem1[132][14] ), .QN(n26586) );
  SDFFX1 \mem1_reg[132][13]  ( .D(n15569), .SI(\mem1[132][12] ), .SE(test_se), 
        .CLK(n1492), .Q(\mem1[132][13] ), .QN(n26587) );
  SDFFX1 \mem1_reg[132][12]  ( .D(n15568), .SI(\mem1[132][11] ), .SE(test_se), 
        .CLK(n1492), .Q(\mem1[132][12] ), .QN(n26588) );
  SDFFX1 \mem1_reg[132][11]  ( .D(n15567), .SI(\mem1[132][10] ), .SE(test_se), 
        .CLK(n1492), .Q(\mem1[132][11] ), .QN(n26589) );
  SDFFX1 \mem1_reg[132][10]  ( .D(n15566), .SI(\mem1[132][9] ), .SE(test_se), 
        .CLK(n1492), .Q(\mem1[132][10] ), .QN(n26590) );
  SDFFX1 \mem1_reg[132][9]  ( .D(n15565), .SI(\mem1[132][8] ), .SE(test_se), 
        .CLK(n1493), .Q(\mem1[132][9] ), .QN(n26591) );
  SDFFX1 \mem1_reg[132][8]  ( .D(n15564), .SI(\mem1[131][15] ), .SE(test_se), 
        .CLK(n1493), .Q(\mem1[132][8] ), .QN(n26592) );
  SDFFX1 \mem1_reg[131][15]  ( .D(n15563), .SI(\mem1[131][14] ), .SE(test_se), 
        .CLK(n1493), .Q(\mem1[131][15] ), .QN(n26593) );
  SDFFX1 \mem1_reg[131][14]  ( .D(n15562), .SI(\mem1[131][13] ), .SE(test_se), 
        .CLK(n1493), .Q(\mem1[131][14] ), .QN(n26594) );
  SDFFX1 \mem1_reg[131][13]  ( .D(n15561), .SI(\mem1[131][12] ), .SE(test_se), 
        .CLK(n1493), .Q(\mem1[131][13] ), .QN(n26595) );
  SDFFX1 \mem1_reg[131][12]  ( .D(n15560), .SI(\mem1[131][11] ), .SE(test_se), 
        .CLK(n1493), .Q(\mem1[131][12] ), .QN(n26596) );
  SDFFX1 \mem1_reg[131][11]  ( .D(n15559), .SI(\mem1[131][10] ), .SE(test_se), 
        .CLK(n1493), .Q(\mem1[131][11] ), .QN(n26597) );
  SDFFX1 \mem1_reg[131][10]  ( .D(n15558), .SI(\mem1[131][9] ), .SE(test_se), 
        .CLK(n1493), .Q(\mem1[131][10] ), .QN(n26598) );
  SDFFX1 \mem1_reg[131][9]  ( .D(n15557), .SI(\mem1[131][8] ), .SE(test_se), 
        .CLK(n1493), .Q(\mem1[131][9] ), .QN(n26599) );
  SDFFX1 \mem1_reg[131][8]  ( .D(n15556), .SI(\mem1[130][15] ), .SE(test_se), 
        .CLK(n1493), .Q(\mem1[131][8] ), .QN(n26600) );
  SDFFX1 \mem1_reg[130][15]  ( .D(n15555), .SI(\mem1[130][14] ), .SE(test_se), 
        .CLK(n1493), .Q(\mem1[130][15] ), .QN(n26601) );
  SDFFX1 \mem1_reg[130][14]  ( .D(n15554), .SI(\mem1[130][13] ), .SE(test_se), 
        .CLK(n1493), .Q(\mem1[130][14] ), .QN(n26602) );
  SDFFX1 \mem1_reg[130][13]  ( .D(n15553), .SI(\mem1[130][12] ), .SE(test_se), 
        .CLK(n1494), .Q(\mem1[130][13] ), .QN(n26603) );
  SDFFX1 \mem1_reg[130][12]  ( .D(n15552), .SI(\mem1[130][11] ), .SE(test_se), 
        .CLK(n1494), .Q(\mem1[130][12] ), .QN(n26604) );
  SDFFX1 \mem1_reg[130][11]  ( .D(n15551), .SI(\mem1[130][10] ), .SE(test_se), 
        .CLK(n1494), .Q(\mem1[130][11] ), .QN(n26605) );
  SDFFX1 \mem1_reg[130][10]  ( .D(n15550), .SI(\mem1[130][9] ), .SE(test_se), 
        .CLK(n1494), .Q(\mem1[130][10] ), .QN(n26606) );
  SDFFX1 \mem1_reg[130][9]  ( .D(n15549), .SI(\mem1[130][8] ), .SE(test_se), 
        .CLK(n1494), .Q(\mem1[130][9] ), .QN(n26607) );
  SDFFX1 \mem1_reg[130][8]  ( .D(n15548), .SI(\mem1[129][15] ), .SE(test_se), 
        .CLK(n1494), .Q(\mem1[130][8] ), .QN(n26608) );
  SDFFX1 \mem1_reg[129][15]  ( .D(n15547), .SI(\mem1[129][14] ), .SE(test_se), 
        .CLK(n1494), .Q(\mem1[129][15] ), .QN(n26609) );
  SDFFX1 \mem1_reg[129][14]  ( .D(n15546), .SI(\mem1[129][13] ), .SE(test_se), 
        .CLK(n1494), .Q(\mem1[129][14] ), .QN(n26610) );
  SDFFX1 \mem1_reg[129][13]  ( .D(n15545), .SI(\mem1[129][12] ), .SE(test_se), 
        .CLK(n1494), .Q(\mem1[129][13] ), .QN(n26611) );
  SDFFX1 \mem1_reg[129][12]  ( .D(n15544), .SI(\mem1[129][11] ), .SE(test_se), 
        .CLK(n1494), .Q(\mem1[129][12] ), .QN(n26612) );
  SDFFX1 \mem1_reg[129][11]  ( .D(n15543), .SI(\mem1[129][10] ), .SE(test_se), 
        .CLK(n1494), .Q(\mem1[129][11] ), .QN(n26613) );
  SDFFX1 \mem1_reg[129][10]  ( .D(n15542), .SI(\mem1[129][9] ), .SE(test_se), 
        .CLK(n1494), .Q(\mem1[129][10] ), .QN(n26614) );
  SDFFX1 \mem1_reg[129][9]  ( .D(n15541), .SI(\mem1[129][8] ), .SE(test_se), 
        .CLK(n1495), .Q(\mem1[129][9] ), .QN(n26615) );
  SDFFX1 \mem1_reg[129][8]  ( .D(n15540), .SI(\mem1[128][15] ), .SE(test_se), 
        .CLK(n1495), .Q(\mem1[129][8] ), .QN(n26616) );
  SDFFX1 \mem1_reg[128][15]  ( .D(n15539), .SI(\mem1[128][14] ), .SE(test_se), 
        .CLK(n1495), .Q(\mem1[128][15] ), .QN(n26617) );
  SDFFX1 \mem1_reg[128][14]  ( .D(n15538), .SI(\mem1[128][13] ), .SE(test_se), 
        .CLK(n1495), .Q(\mem1[128][14] ), .QN(n26618) );
  SDFFX1 \mem1_reg[128][13]  ( .D(n15537), .SI(\mem1[128][12] ), .SE(test_se), 
        .CLK(n1495), .Q(\mem1[128][13] ), .QN(n26619) );
  SDFFX1 \mem1_reg[128][12]  ( .D(n15536), .SI(\mem1[128][11] ), .SE(test_se), 
        .CLK(n1495), .Q(\mem1[128][12] ), .QN(n26620) );
  SDFFX1 \mem1_reg[128][11]  ( .D(n15535), .SI(\mem1[128][10] ), .SE(test_se), 
        .CLK(n1495), .Q(\mem1[128][11] ), .QN(n26621) );
  SDFFX1 \mem1_reg[128][10]  ( .D(n15534), .SI(\mem1[128][9] ), .SE(test_se), 
        .CLK(n1495), .Q(\mem1[128][10] ), .QN(n26622) );
  SDFFX1 \mem1_reg[128][9]  ( .D(n15533), .SI(\mem1[128][8] ), .SE(test_se), 
        .CLK(n1495), .Q(\mem1[128][9] ), .QN(n26623) );
  SDFFX1 \mem1_reg[128][8]  ( .D(n15532), .SI(\mem1[127][15] ), .SE(test_se), 
        .CLK(n1495), .Q(\mem1[128][8] ), .QN(n26624) );
  SDFFX1 \mem1_reg[127][15]  ( .D(n15531), .SI(\mem1[127][14] ), .SE(test_se), 
        .CLK(n1495), .Q(\mem1[127][15] ), .QN(n26625) );
  SDFFX1 \mem1_reg[127][14]  ( .D(n15530), .SI(\mem1[127][13] ), .SE(test_se), 
        .CLK(n1495), .Q(\mem1[127][14] ), .QN(n26626) );
  SDFFX1 \mem1_reg[127][13]  ( .D(n15529), .SI(\mem1[127][12] ), .SE(test_se), 
        .CLK(n1496), .Q(\mem1[127][13] ), .QN(n26627) );
  SDFFX1 \mem1_reg[127][12]  ( .D(n15528), .SI(\mem1[127][11] ), .SE(test_se), 
        .CLK(n1496), .Q(\mem1[127][12] ), .QN(n26628) );
  SDFFX1 \mem1_reg[127][11]  ( .D(n15527), .SI(\mem1[127][10] ), .SE(test_se), 
        .CLK(n1496), .Q(\mem1[127][11] ), .QN(n26629) );
  SDFFX1 \mem1_reg[127][10]  ( .D(n15526), .SI(\mem1[127][9] ), .SE(test_se), 
        .CLK(n1496), .Q(\mem1[127][10] ), .QN(n26630) );
  SDFFX1 \mem1_reg[127][9]  ( .D(n15525), .SI(\mem1[127][8] ), .SE(test_se), 
        .CLK(n1496), .Q(\mem1[127][9] ), .QN(n26631) );
  SDFFX1 \mem1_reg[127][8]  ( .D(n15524), .SI(\mem1[126][15] ), .SE(test_se), 
        .CLK(n1496), .Q(\mem1[127][8] ), .QN(n26632) );
  SDFFX1 \mem1_reg[126][15]  ( .D(n15523), .SI(\mem1[126][14] ), .SE(test_se), 
        .CLK(n1496), .Q(\mem1[126][15] ), .QN(n26633) );
  SDFFX1 \mem1_reg[126][14]  ( .D(n15522), .SI(\mem1[126][13] ), .SE(test_se), 
        .CLK(n1496), .Q(\mem1[126][14] ), .QN(n26634) );
  SDFFX1 \mem1_reg[126][13]  ( .D(n15521), .SI(\mem1[126][12] ), .SE(test_se), 
        .CLK(n1496), .Q(\mem1[126][13] ), .QN(n26635) );
  SDFFX1 \mem1_reg[126][12]  ( .D(n15520), .SI(\mem1[126][11] ), .SE(test_se), 
        .CLK(n1496), .Q(\mem1[126][12] ), .QN(n26636) );
  SDFFX1 \mem1_reg[126][11]  ( .D(n15519), .SI(\mem1[126][10] ), .SE(test_se), 
        .CLK(n1496), .Q(\mem1[126][11] ), .QN(n26637) );
  SDFFX1 \mem1_reg[126][10]  ( .D(n15518), .SI(\mem1[126][9] ), .SE(test_se), 
        .CLK(n1496), .Q(\mem1[126][10] ), .QN(n26638) );
  SDFFX1 \mem1_reg[126][9]  ( .D(n15517), .SI(\mem1[126][8] ), .SE(test_se), 
        .CLK(n1497), .Q(\mem1[126][9] ), .QN(n26639) );
  SDFFX1 \mem1_reg[126][8]  ( .D(n15516), .SI(\mem1[125][15] ), .SE(test_se), 
        .CLK(n1497), .Q(\mem1[126][8] ), .QN(n26640) );
  SDFFX1 \mem1_reg[125][15]  ( .D(n15515), .SI(\mem1[125][14] ), .SE(test_se), 
        .CLK(n1497), .Q(\mem1[125][15] ), .QN(n26641) );
  SDFFX1 \mem1_reg[125][14]  ( .D(n15514), .SI(\mem1[125][13] ), .SE(test_se), 
        .CLK(n1497), .Q(\mem1[125][14] ), .QN(n26642) );
  SDFFX1 \mem1_reg[125][13]  ( .D(n15513), .SI(\mem1[125][12] ), .SE(test_se), 
        .CLK(n1497), .Q(\mem1[125][13] ), .QN(n26643) );
  SDFFX1 \mem1_reg[125][12]  ( .D(n15512), .SI(\mem1[125][11] ), .SE(test_se), 
        .CLK(n1497), .Q(\mem1[125][12] ), .QN(n26644) );
  SDFFX1 \mem1_reg[125][11]  ( .D(n15511), .SI(\mem1[125][10] ), .SE(test_se), 
        .CLK(n1497), .Q(\mem1[125][11] ), .QN(n26645) );
  SDFFX1 \mem1_reg[125][10]  ( .D(n15510), .SI(\mem1[125][9] ), .SE(test_se), 
        .CLK(n1497), .Q(\mem1[125][10] ), .QN(n26646) );
  SDFFX1 \mem1_reg[125][9]  ( .D(n15509), .SI(\mem1[125][8] ), .SE(test_se), 
        .CLK(n1497), .Q(\mem1[125][9] ), .QN(n26647) );
  SDFFX1 \mem1_reg[125][8]  ( .D(n15508), .SI(\mem1[124][15] ), .SE(test_se), 
        .CLK(n1497), .Q(\mem1[125][8] ), .QN(n26648) );
  SDFFX1 \mem1_reg[124][15]  ( .D(n15507), .SI(\mem1[124][14] ), .SE(test_se), 
        .CLK(n1497), .Q(\mem1[124][15] ), .QN(n26649) );
  SDFFX1 \mem1_reg[124][14]  ( .D(n15506), .SI(\mem1[124][13] ), .SE(test_se), 
        .CLK(n1497), .Q(\mem1[124][14] ), .QN(n26650) );
  SDFFX1 \mem1_reg[124][13]  ( .D(n15505), .SI(\mem1[124][12] ), .SE(test_se), 
        .CLK(n1498), .Q(\mem1[124][13] ), .QN(n26651) );
  SDFFX1 \mem1_reg[124][12]  ( .D(n15504), .SI(\mem1[124][11] ), .SE(test_se), 
        .CLK(n1498), .Q(\mem1[124][12] ), .QN(n26652) );
  SDFFX1 \mem1_reg[124][11]  ( .D(n15503), .SI(\mem1[124][10] ), .SE(test_se), 
        .CLK(n1498), .Q(\mem1[124][11] ), .QN(n26653) );
  SDFFX1 \mem1_reg[124][10]  ( .D(n15502), .SI(\mem1[124][9] ), .SE(test_se), 
        .CLK(n1498), .Q(\mem1[124][10] ), .QN(n26654) );
  SDFFX1 \mem1_reg[124][9]  ( .D(n15501), .SI(\mem1[124][8] ), .SE(test_se), 
        .CLK(n1498), .Q(\mem1[124][9] ), .QN(n26655) );
  SDFFX1 \mem1_reg[124][8]  ( .D(n15500), .SI(\mem1[123][15] ), .SE(test_se), 
        .CLK(n1498), .Q(\mem1[124][8] ), .QN(n26656) );
  SDFFX1 \mem1_reg[123][15]  ( .D(n15499), .SI(\mem1[123][14] ), .SE(test_se), 
        .CLK(n1498), .Q(\mem1[123][15] ), .QN(n26657) );
  SDFFX1 \mem1_reg[123][14]  ( .D(n15498), .SI(\mem1[123][13] ), .SE(test_se), 
        .CLK(n1498), .Q(\mem1[123][14] ), .QN(n26658) );
  SDFFX1 \mem1_reg[123][13]  ( .D(n15497), .SI(\mem1[123][12] ), .SE(test_se), 
        .CLK(n1498), .Q(\mem1[123][13] ), .QN(n26659) );
  SDFFX1 \mem1_reg[123][12]  ( .D(n15496), .SI(\mem1[123][11] ), .SE(test_se), 
        .CLK(n1498), .Q(\mem1[123][12] ), .QN(n26660) );
  SDFFX1 \mem1_reg[123][11]  ( .D(n15495), .SI(\mem1[123][10] ), .SE(test_se), 
        .CLK(n1498), .Q(\mem1[123][11] ), .QN(n26661) );
  SDFFX1 \mem1_reg[123][10]  ( .D(n15494), .SI(\mem1[123][9] ), .SE(test_se), 
        .CLK(n1498), .Q(\mem1[123][10] ), .QN(n26662) );
  SDFFX1 \mem1_reg[123][9]  ( .D(n15493), .SI(\mem1[123][8] ), .SE(test_se), 
        .CLK(n1499), .Q(\mem1[123][9] ), .QN(n26663) );
  SDFFX1 \mem1_reg[123][8]  ( .D(n15492), .SI(\mem1[122][15] ), .SE(test_se), 
        .CLK(n1499), .Q(\mem1[123][8] ), .QN(n26664) );
  SDFFX1 \mem1_reg[122][15]  ( .D(n15491), .SI(\mem1[122][14] ), .SE(test_se), 
        .CLK(n1499), .Q(\mem1[122][15] ), .QN(n26665) );
  SDFFX1 \mem1_reg[122][14]  ( .D(n15490), .SI(\mem1[122][13] ), .SE(test_se), 
        .CLK(n1499), .Q(\mem1[122][14] ), .QN(n26666) );
  SDFFX1 \mem1_reg[122][13]  ( .D(n15489), .SI(\mem1[122][12] ), .SE(test_se), 
        .CLK(n1499), .Q(\mem1[122][13] ), .QN(n26667) );
  SDFFX1 \mem1_reg[122][12]  ( .D(n15488), .SI(\mem1[122][11] ), .SE(test_se), 
        .CLK(n1499), .Q(\mem1[122][12] ), .QN(n26668) );
  SDFFX1 \mem1_reg[122][11]  ( .D(n15487), .SI(\mem1[122][10] ), .SE(test_se), 
        .CLK(n1499), .Q(\mem1[122][11] ), .QN(n26669) );
  SDFFX1 \mem1_reg[122][10]  ( .D(n15486), .SI(\mem1[122][9] ), .SE(test_se), 
        .CLK(n1499), .Q(\mem1[122][10] ), .QN(n26670) );
  SDFFX1 \mem1_reg[122][9]  ( .D(n15485), .SI(\mem1[122][8] ), .SE(test_se), 
        .CLK(n1499), .Q(\mem1[122][9] ), .QN(n26671) );
  SDFFX1 \mem1_reg[122][8]  ( .D(n15484), .SI(\mem1[121][15] ), .SE(test_se), 
        .CLK(n1499), .Q(\mem1[122][8] ), .QN(n26672) );
  SDFFX1 \mem1_reg[121][15]  ( .D(n15483), .SI(\mem1[121][14] ), .SE(test_se), 
        .CLK(n1499), .Q(\mem1[121][15] ), .QN(n26673) );
  SDFFX1 \mem1_reg[121][14]  ( .D(n15482), .SI(\mem1[121][13] ), .SE(test_se), 
        .CLK(n1499), .Q(\mem1[121][14] ), .QN(n26674) );
  SDFFX1 \mem1_reg[121][13]  ( .D(n15481), .SI(\mem1[121][12] ), .SE(test_se), 
        .CLK(n1500), .Q(\mem1[121][13] ), .QN(n26675) );
  SDFFX1 \mem1_reg[121][12]  ( .D(n15480), .SI(\mem1[121][11] ), .SE(test_se), 
        .CLK(n1500), .Q(\mem1[121][12] ), .QN(n26676) );
  SDFFX1 \mem1_reg[121][11]  ( .D(n15479), .SI(\mem1[121][10] ), .SE(test_se), 
        .CLK(n1500), .Q(\mem1[121][11] ), .QN(n26677) );
  SDFFX1 \mem1_reg[121][10]  ( .D(n15478), .SI(\mem1[121][9] ), .SE(test_se), 
        .CLK(n1500), .Q(\mem1[121][10] ), .QN(n26678) );
  SDFFX1 \mem1_reg[121][9]  ( .D(n15477), .SI(\mem1[121][8] ), .SE(test_se), 
        .CLK(n1500), .Q(\mem1[121][9] ), .QN(n26679) );
  SDFFX1 \mem1_reg[121][8]  ( .D(n15476), .SI(\mem1[120][15] ), .SE(test_se), 
        .CLK(n1500), .Q(\mem1[121][8] ), .QN(n26680) );
  SDFFX1 \mem1_reg[120][15]  ( .D(n15475), .SI(\mem1[120][14] ), .SE(test_se), 
        .CLK(n1500), .Q(\mem1[120][15] ), .QN(n26681) );
  SDFFX1 \mem1_reg[120][14]  ( .D(n15474), .SI(\mem1[120][13] ), .SE(test_se), 
        .CLK(n1500), .Q(\mem1[120][14] ), .QN(n26682) );
  SDFFX1 \mem1_reg[120][13]  ( .D(n15473), .SI(\mem1[120][12] ), .SE(test_se), 
        .CLK(n1500), .Q(\mem1[120][13] ), .QN(n26683) );
  SDFFX1 \mem1_reg[120][12]  ( .D(n15472), .SI(\mem1[120][11] ), .SE(test_se), 
        .CLK(n1500), .Q(\mem1[120][12] ), .QN(n26684) );
  SDFFX1 \mem1_reg[120][11]  ( .D(n15471), .SI(\mem1[120][10] ), .SE(test_se), 
        .CLK(n1500), .Q(\mem1[120][11] ), .QN(n26685) );
  SDFFX1 \mem1_reg[120][10]  ( .D(n15470), .SI(\mem1[120][9] ), .SE(test_se), 
        .CLK(n1500), .Q(\mem1[120][10] ), .QN(n26686) );
  SDFFX1 \mem1_reg[120][9]  ( .D(n15469), .SI(\mem1[120][8] ), .SE(test_se), 
        .CLK(n1501), .Q(\mem1[120][9] ), .QN(n26687) );
  SDFFX1 \mem1_reg[120][8]  ( .D(n15468), .SI(\mem1[119][15] ), .SE(test_se), 
        .CLK(n1501), .Q(\mem1[120][8] ), .QN(n26688) );
  SDFFX1 \mem1_reg[119][15]  ( .D(n15467), .SI(\mem1[119][14] ), .SE(test_se), 
        .CLK(n1501), .Q(\mem1[119][15] ), .QN(n26689) );
  SDFFX1 \mem1_reg[119][14]  ( .D(n15466), .SI(\mem1[119][13] ), .SE(test_se), 
        .CLK(n1501), .Q(\mem1[119][14] ), .QN(n26690) );
  SDFFX1 \mem1_reg[119][13]  ( .D(n15465), .SI(\mem1[119][12] ), .SE(test_se), 
        .CLK(n1501), .Q(\mem1[119][13] ), .QN(n26691) );
  SDFFX1 \mem1_reg[119][12]  ( .D(n15464), .SI(\mem1[119][11] ), .SE(test_se), 
        .CLK(n1501), .Q(\mem1[119][12] ), .QN(n26692) );
  SDFFX1 \mem1_reg[119][11]  ( .D(n15463), .SI(\mem1[119][10] ), .SE(test_se), 
        .CLK(n1501), .Q(\mem1[119][11] ), .QN(n26693) );
  SDFFX1 \mem1_reg[119][10]  ( .D(n15462), .SI(\mem1[119][9] ), .SE(test_se), 
        .CLK(n1501), .Q(\mem1[119][10] ), .QN(n26694) );
  SDFFX1 \mem1_reg[119][9]  ( .D(n15461), .SI(\mem1[119][8] ), .SE(test_se), 
        .CLK(n1501), .Q(\mem1[119][9] ), .QN(n26695) );
  SDFFX1 \mem1_reg[119][8]  ( .D(n15460), .SI(\mem1[118][15] ), .SE(test_se), 
        .CLK(n1501), .Q(\mem1[119][8] ), .QN(n26696) );
  SDFFX1 \mem1_reg[118][15]  ( .D(n15459), .SI(\mem1[118][14] ), .SE(test_se), 
        .CLK(n1501), .Q(\mem1[118][15] ), .QN(n26697) );
  SDFFX1 \mem1_reg[118][14]  ( .D(n15458), .SI(\mem1[118][13] ), .SE(test_se), 
        .CLK(n1501), .Q(\mem1[118][14] ), .QN(n26698) );
  SDFFX1 \mem1_reg[118][13]  ( .D(n15457), .SI(\mem1[118][12] ), .SE(test_se), 
        .CLK(n1502), .Q(\mem1[118][13] ), .QN(n26699) );
  SDFFX1 \mem1_reg[118][12]  ( .D(n15456), .SI(\mem1[118][11] ), .SE(test_se), 
        .CLK(n1502), .Q(\mem1[118][12] ), .QN(n26700) );
  SDFFX1 \mem1_reg[118][11]  ( .D(n15455), .SI(\mem1[118][10] ), .SE(test_se), 
        .CLK(n1502), .Q(\mem1[118][11] ), .QN(n26701) );
  SDFFX1 \mem1_reg[118][10]  ( .D(n15454), .SI(\mem1[118][9] ), .SE(test_se), 
        .CLK(n1502), .Q(\mem1[118][10] ), .QN(n26702) );
  SDFFX1 \mem1_reg[118][9]  ( .D(n15453), .SI(\mem1[118][8] ), .SE(test_se), 
        .CLK(n1502), .Q(\mem1[118][9] ), .QN(n26703) );
  SDFFX1 \mem1_reg[118][8]  ( .D(n15452), .SI(\mem1[117][15] ), .SE(test_se), 
        .CLK(n1502), .Q(\mem1[118][8] ), .QN(n26704) );
  SDFFX1 \mem1_reg[117][15]  ( .D(n15451), .SI(\mem1[117][14] ), .SE(test_se), 
        .CLK(n1502), .Q(\mem1[117][15] ), .QN(n26705) );
  SDFFX1 \mem1_reg[117][14]  ( .D(n15450), .SI(\mem1[117][13] ), .SE(test_se), 
        .CLK(n1502), .Q(\mem1[117][14] ), .QN(n26706) );
  SDFFX1 \mem1_reg[117][13]  ( .D(n15449), .SI(\mem1[117][12] ), .SE(test_se), 
        .CLK(n1502), .Q(\mem1[117][13] ), .QN(n26707) );
  SDFFX1 \mem1_reg[117][12]  ( .D(n15448), .SI(\mem1[117][11] ), .SE(test_se), 
        .CLK(n1502), .Q(\mem1[117][12] ), .QN(n26708) );
  SDFFX1 \mem1_reg[117][11]  ( .D(n15447), .SI(\mem1[117][10] ), .SE(test_se), 
        .CLK(n1502), .Q(\mem1[117][11] ), .QN(n26709) );
  SDFFX1 \mem1_reg[117][10]  ( .D(n15446), .SI(\mem1[117][9] ), .SE(test_se), 
        .CLK(n1502), .Q(\mem1[117][10] ), .QN(n26710) );
  SDFFX1 \mem1_reg[117][9]  ( .D(n15445), .SI(\mem1[117][8] ), .SE(test_se), 
        .CLK(n1503), .Q(\mem1[117][9] ), .QN(n26711) );
  SDFFX1 \mem1_reg[117][8]  ( .D(n15444), .SI(\mem1[116][15] ), .SE(test_se), 
        .CLK(n1503), .Q(\mem1[117][8] ), .QN(n26712) );
  SDFFX1 \mem1_reg[116][15]  ( .D(n15443), .SI(\mem1[116][14] ), .SE(test_se), 
        .CLK(n1503), .Q(\mem1[116][15] ), .QN(n26713) );
  SDFFX1 \mem1_reg[116][14]  ( .D(n15442), .SI(\mem1[116][13] ), .SE(test_se), 
        .CLK(n1503), .Q(\mem1[116][14] ), .QN(n26714) );
  SDFFX1 \mem1_reg[116][13]  ( .D(n15441), .SI(\mem1[116][12] ), .SE(test_se), 
        .CLK(n1503), .Q(\mem1[116][13] ), .QN(n26715) );
  SDFFX1 \mem1_reg[116][12]  ( .D(n15440), .SI(\mem1[116][11] ), .SE(test_se), 
        .CLK(n1503), .Q(\mem1[116][12] ), .QN(n26716) );
  SDFFX1 \mem1_reg[116][11]  ( .D(n15439), .SI(\mem1[116][10] ), .SE(test_se), 
        .CLK(n1503), .Q(\mem1[116][11] ), .QN(n26717) );
  SDFFX1 \mem1_reg[116][10]  ( .D(n15438), .SI(\mem1[116][9] ), .SE(test_se), 
        .CLK(n1503), .Q(\mem1[116][10] ), .QN(n26718) );
  SDFFX1 \mem1_reg[116][9]  ( .D(n15437), .SI(\mem1[116][8] ), .SE(test_se), 
        .CLK(n1503), .Q(\mem1[116][9] ), .QN(n26719) );
  SDFFX1 \mem1_reg[116][8]  ( .D(n15436), .SI(\mem1[115][15] ), .SE(test_se), 
        .CLK(n1503), .Q(\mem1[116][8] ), .QN(n26720) );
  SDFFX1 \mem1_reg[115][15]  ( .D(n15435), .SI(\mem1[115][14] ), .SE(test_se), 
        .CLK(n1503), .Q(\mem1[115][15] ), .QN(n26721) );
  SDFFX1 \mem1_reg[115][14]  ( .D(n15434), .SI(\mem1[115][13] ), .SE(test_se), 
        .CLK(n1503), .Q(\mem1[115][14] ), .QN(n26722) );
  SDFFX1 \mem1_reg[115][13]  ( .D(n15433), .SI(\mem1[115][12] ), .SE(test_se), 
        .CLK(n1504), .Q(\mem1[115][13] ), .QN(n26723) );
  SDFFX1 \mem1_reg[115][12]  ( .D(n15432), .SI(\mem1[115][11] ), .SE(test_se), 
        .CLK(n1504), .Q(\mem1[115][12] ), .QN(n26724) );
  SDFFX1 \mem1_reg[115][11]  ( .D(n15431), .SI(\mem1[115][10] ), .SE(test_se), 
        .CLK(n1504), .Q(\mem1[115][11] ), .QN(n26725) );
  SDFFX1 \mem1_reg[115][10]  ( .D(n15430), .SI(\mem1[115][9] ), .SE(test_se), 
        .CLK(n1504), .Q(\mem1[115][10] ), .QN(n26726) );
  SDFFX1 \mem1_reg[115][9]  ( .D(n15429), .SI(\mem1[115][8] ), .SE(test_se), 
        .CLK(n1504), .Q(\mem1[115][9] ), .QN(n26727) );
  SDFFX1 \mem1_reg[115][8]  ( .D(n15428), .SI(\mem1[114][15] ), .SE(test_se), 
        .CLK(n1504), .Q(\mem1[115][8] ), .QN(n26728) );
  SDFFX1 \mem1_reg[114][15]  ( .D(n15427), .SI(\mem1[114][14] ), .SE(test_se), 
        .CLK(n1504), .Q(\mem1[114][15] ), .QN(n26729) );
  SDFFX1 \mem1_reg[114][14]  ( .D(n15426), .SI(\mem1[114][13] ), .SE(test_se), 
        .CLK(n1504), .Q(\mem1[114][14] ), .QN(n26730) );
  SDFFX1 \mem1_reg[114][13]  ( .D(n15425), .SI(\mem1[114][12] ), .SE(test_se), 
        .CLK(n1504), .Q(\mem1[114][13] ), .QN(n26731) );
  SDFFX1 \mem1_reg[114][12]  ( .D(n15424), .SI(\mem1[114][11] ), .SE(test_se), 
        .CLK(n1504), .Q(\mem1[114][12] ), .QN(n26732) );
  SDFFX1 \mem1_reg[114][11]  ( .D(n15423), .SI(\mem1[114][10] ), .SE(test_se), 
        .CLK(n1504), .Q(\mem1[114][11] ), .QN(n26733) );
  SDFFX1 \mem1_reg[114][10]  ( .D(n15422), .SI(\mem1[114][9] ), .SE(test_se), 
        .CLK(n1504), .Q(\mem1[114][10] ), .QN(n26734) );
  SDFFX1 \mem1_reg[114][9]  ( .D(n15421), .SI(\mem1[114][8] ), .SE(test_se), 
        .CLK(n1505), .Q(\mem1[114][9] ), .QN(n26735) );
  SDFFX1 \mem1_reg[114][8]  ( .D(n15420), .SI(\mem1[113][15] ), .SE(test_se), 
        .CLK(n1505), .Q(\mem1[114][8] ), .QN(n26736) );
  SDFFX1 \mem1_reg[113][15]  ( .D(n15419), .SI(\mem1[113][14] ), .SE(test_se), 
        .CLK(n1505), .Q(\mem1[113][15] ), .QN(n26737) );
  SDFFX1 \mem1_reg[113][14]  ( .D(n15418), .SI(\mem1[113][13] ), .SE(test_se), 
        .CLK(n1505), .Q(\mem1[113][14] ), .QN(n26738) );
  SDFFX1 \mem1_reg[113][13]  ( .D(n15417), .SI(\mem1[113][12] ), .SE(test_se), 
        .CLK(n1505), .Q(\mem1[113][13] ), .QN(n26739) );
  SDFFX1 \mem1_reg[113][12]  ( .D(n15416), .SI(\mem1[113][11] ), .SE(test_se), 
        .CLK(n1505), .Q(\mem1[113][12] ), .QN(n26740) );
  SDFFX1 \mem1_reg[113][11]  ( .D(n15415), .SI(\mem1[113][10] ), .SE(test_se), 
        .CLK(n1505), .Q(\mem1[113][11] ), .QN(n26741) );
  SDFFX1 \mem1_reg[113][10]  ( .D(n15414), .SI(\mem1[113][9] ), .SE(test_se), 
        .CLK(n1505), .Q(\mem1[113][10] ), .QN(n26742) );
  SDFFX1 \mem1_reg[113][9]  ( .D(n15413), .SI(\mem1[113][8] ), .SE(test_se), 
        .CLK(n1505), .Q(\mem1[113][9] ), .QN(n26743) );
  SDFFX1 \mem1_reg[113][8]  ( .D(n15412), .SI(\mem1[112][15] ), .SE(test_se), 
        .CLK(n1505), .Q(\mem1[113][8] ), .QN(n26744) );
  SDFFX1 \mem1_reg[112][15]  ( .D(n15411), .SI(\mem1[112][14] ), .SE(test_se), 
        .CLK(n1505), .Q(\mem1[112][15] ), .QN(n26745) );
  SDFFX1 \mem1_reg[112][14]  ( .D(n15410), .SI(\mem1[112][13] ), .SE(test_se), 
        .CLK(n1505), .Q(\mem1[112][14] ), .QN(n26746) );
  SDFFX1 \mem1_reg[112][13]  ( .D(n15409), .SI(\mem1[112][12] ), .SE(test_se), 
        .CLK(n1506), .Q(\mem1[112][13] ), .QN(n26747) );
  SDFFX1 \mem1_reg[112][12]  ( .D(n15408), .SI(\mem1[112][11] ), .SE(test_se), 
        .CLK(n1506), .Q(\mem1[112][12] ), .QN(n26748) );
  SDFFX1 \mem1_reg[112][11]  ( .D(n15407), .SI(\mem1[112][10] ), .SE(test_se), 
        .CLK(n1506), .Q(\mem1[112][11] ), .QN(n26749) );
  SDFFX1 \mem1_reg[112][10]  ( .D(n15406), .SI(\mem1[112][9] ), .SE(test_se), 
        .CLK(n1506), .Q(\mem1[112][10] ), .QN(n26750) );
  SDFFX1 \mem1_reg[112][9]  ( .D(n15405), .SI(\mem1[112][8] ), .SE(test_se), 
        .CLK(n1506), .Q(\mem1[112][9] ), .QN(n26751) );
  SDFFX1 \mem1_reg[112][8]  ( .D(n15404), .SI(\mem1[111][15] ), .SE(test_se), 
        .CLK(n1506), .Q(\mem1[112][8] ), .QN(n26752) );
  SDFFX1 \mem1_reg[111][15]  ( .D(n15403), .SI(\mem1[111][14] ), .SE(test_se), 
        .CLK(n1506), .Q(\mem1[111][15] ), .QN(n26753) );
  SDFFX1 \mem1_reg[111][14]  ( .D(n15402), .SI(\mem1[111][13] ), .SE(test_se), 
        .CLK(n1506), .Q(\mem1[111][14] ), .QN(n26754) );
  SDFFX1 \mem1_reg[111][13]  ( .D(n15401), .SI(\mem1[111][12] ), .SE(test_se), 
        .CLK(n1506), .Q(\mem1[111][13] ), .QN(n26755) );
  SDFFX1 \mem1_reg[111][12]  ( .D(n15400), .SI(\mem1[111][11] ), .SE(test_se), 
        .CLK(n1506), .Q(\mem1[111][12] ), .QN(n26756) );
  SDFFX1 \mem1_reg[111][11]  ( .D(n15399), .SI(\mem1[111][10] ), .SE(test_se), 
        .CLK(n1506), .Q(\mem1[111][11] ), .QN(n26757) );
  SDFFX1 \mem1_reg[111][10]  ( .D(n15398), .SI(\mem1[111][9] ), .SE(test_se), 
        .CLK(n1506), .Q(\mem1[111][10] ), .QN(n26758) );
  SDFFX1 \mem1_reg[111][9]  ( .D(n15397), .SI(\mem1[111][8] ), .SE(test_se), 
        .CLK(n1507), .Q(\mem1[111][9] ), .QN(n26759) );
  SDFFX1 \mem1_reg[111][8]  ( .D(n15396), .SI(\mem1[110][15] ), .SE(test_se), 
        .CLK(n1507), .Q(\mem1[111][8] ), .QN(n26760) );
  SDFFX1 \mem1_reg[110][15]  ( .D(n15395), .SI(\mem1[110][14] ), .SE(test_se), 
        .CLK(n1507), .Q(\mem1[110][15] ), .QN(n26761) );
  SDFFX1 \mem1_reg[110][14]  ( .D(n15394), .SI(\mem1[110][13] ), .SE(test_se), 
        .CLK(n1507), .Q(\mem1[110][14] ), .QN(n26762) );
  SDFFX1 \mem1_reg[110][13]  ( .D(n15393), .SI(\mem1[110][12] ), .SE(test_se), 
        .CLK(n1507), .Q(\mem1[110][13] ), .QN(n26763) );
  SDFFX1 \mem1_reg[110][12]  ( .D(n15392), .SI(\mem1[110][11] ), .SE(test_se), 
        .CLK(n1507), .Q(\mem1[110][12] ), .QN(n26764) );
  SDFFX1 \mem1_reg[110][11]  ( .D(n15391), .SI(\mem1[110][10] ), .SE(test_se), 
        .CLK(n1507), .Q(\mem1[110][11] ), .QN(n26765) );
  SDFFX1 \mem1_reg[110][10]  ( .D(n15390), .SI(\mem1[110][9] ), .SE(test_se), 
        .CLK(n1507), .Q(\mem1[110][10] ), .QN(n26766) );
  SDFFX1 \mem1_reg[110][9]  ( .D(n15389), .SI(\mem1[110][8] ), .SE(test_se), 
        .CLK(n1507), .Q(\mem1[110][9] ), .QN(n26767) );
  SDFFX1 \mem1_reg[110][8]  ( .D(n15388), .SI(\mem1[109][15] ), .SE(test_se), 
        .CLK(n1507), .Q(\mem1[110][8] ), .QN(n26768) );
  SDFFX1 \mem1_reg[109][15]  ( .D(n15387), .SI(\mem1[109][14] ), .SE(test_se), 
        .CLK(n1507), .Q(\mem1[109][15] ), .QN(n26769) );
  SDFFX1 \mem1_reg[109][14]  ( .D(n15386), .SI(\mem1[109][13] ), .SE(test_se), 
        .CLK(n1507), .Q(\mem1[109][14] ), .QN(n26770) );
  SDFFX1 \mem1_reg[109][13]  ( .D(n15385), .SI(\mem1[109][12] ), .SE(test_se), 
        .CLK(n1508), .Q(\mem1[109][13] ), .QN(n26771) );
  SDFFX1 \mem1_reg[109][12]  ( .D(n15384), .SI(\mem1[109][11] ), .SE(test_se), 
        .CLK(n1508), .Q(\mem1[109][12] ), .QN(n26772) );
  SDFFX1 \mem1_reg[109][11]  ( .D(n15383), .SI(\mem1[109][10] ), .SE(test_se), 
        .CLK(n1508), .Q(\mem1[109][11] ), .QN(n26773) );
  SDFFX1 \mem1_reg[109][10]  ( .D(n15382), .SI(\mem1[109][9] ), .SE(test_se), 
        .CLK(n1508), .Q(\mem1[109][10] ), .QN(n26774) );
  SDFFX1 \mem1_reg[109][9]  ( .D(n15381), .SI(\mem1[109][8] ), .SE(test_se), 
        .CLK(n1508), .Q(\mem1[109][9] ), .QN(n26775) );
  SDFFX1 \mem1_reg[109][8]  ( .D(n15380), .SI(\mem1[108][15] ), .SE(test_se), 
        .CLK(n1508), .Q(\mem1[109][8] ), .QN(n26776) );
  SDFFX1 \mem1_reg[108][15]  ( .D(n15379), .SI(\mem1[108][14] ), .SE(test_se), 
        .CLK(n1508), .Q(\mem1[108][15] ), .QN(n26777) );
  SDFFX1 \mem1_reg[108][14]  ( .D(n15378), .SI(\mem1[108][13] ), .SE(test_se), 
        .CLK(n1508), .Q(\mem1[108][14] ), .QN(n26778) );
  SDFFX1 \mem1_reg[108][13]  ( .D(n15377), .SI(\mem1[108][12] ), .SE(test_se), 
        .CLK(n1508), .Q(\mem1[108][13] ), .QN(n26779) );
  SDFFX1 \mem1_reg[108][12]  ( .D(n15376), .SI(\mem1[108][11] ), .SE(test_se), 
        .CLK(n1508), .Q(\mem1[108][12] ), .QN(n26780) );
  SDFFX1 \mem1_reg[108][11]  ( .D(n15375), .SI(\mem1[108][10] ), .SE(test_se), 
        .CLK(n1508), .Q(\mem1[108][11] ), .QN(n26781) );
  SDFFX1 \mem1_reg[108][10]  ( .D(n15374), .SI(\mem1[108][9] ), .SE(test_se), 
        .CLK(n1508), .Q(\mem1[108][10] ), .QN(n26782) );
  SDFFX1 \mem1_reg[108][9]  ( .D(n15373), .SI(\mem1[108][8] ), .SE(test_se), 
        .CLK(n1509), .Q(\mem1[108][9] ), .QN(n26783) );
  SDFFX1 \mem1_reg[108][8]  ( .D(n15372), .SI(\mem1[107][15] ), .SE(test_se), 
        .CLK(n1509), .Q(\mem1[108][8] ), .QN(n26784) );
  SDFFX1 \mem1_reg[107][15]  ( .D(n15371), .SI(\mem1[107][14] ), .SE(test_se), 
        .CLK(n1509), .Q(\mem1[107][15] ), .QN(n26785) );
  SDFFX1 \mem1_reg[107][14]  ( .D(n15370), .SI(\mem1[107][13] ), .SE(test_se), 
        .CLK(n1509), .Q(\mem1[107][14] ), .QN(n26786) );
  SDFFX1 \mem1_reg[107][13]  ( .D(n15369), .SI(\mem1[107][12] ), .SE(test_se), 
        .CLK(n1509), .Q(\mem1[107][13] ), .QN(n26787) );
  SDFFX1 \mem1_reg[107][12]  ( .D(n15368), .SI(\mem1[107][11] ), .SE(test_se), 
        .CLK(n1509), .Q(\mem1[107][12] ), .QN(n26788) );
  SDFFX1 \mem1_reg[107][11]  ( .D(n15367), .SI(\mem1[107][10] ), .SE(test_se), 
        .CLK(n1509), .Q(\mem1[107][11] ), .QN(n26789) );
  SDFFX1 \mem1_reg[107][10]  ( .D(n15366), .SI(\mem1[107][9] ), .SE(test_se), 
        .CLK(n1509), .Q(\mem1[107][10] ), .QN(n26790) );
  SDFFX1 \mem1_reg[107][9]  ( .D(n15365), .SI(\mem1[107][8] ), .SE(test_se), 
        .CLK(n1509), .Q(\mem1[107][9] ), .QN(n26791) );
  SDFFX1 \mem1_reg[107][8]  ( .D(n15364), .SI(\mem1[106][15] ), .SE(test_se), 
        .CLK(n1509), .Q(\mem1[107][8] ), .QN(n26792) );
  SDFFX1 \mem1_reg[106][15]  ( .D(n15363), .SI(\mem1[106][14] ), .SE(test_se), 
        .CLK(n1509), .Q(\mem1[106][15] ), .QN(n26793) );
  SDFFX1 \mem1_reg[106][14]  ( .D(n15362), .SI(\mem1[106][13] ), .SE(test_se), 
        .CLK(n1509), .Q(\mem1[106][14] ), .QN(n26794) );
  SDFFX1 \mem1_reg[106][13]  ( .D(n15361), .SI(\mem1[106][12] ), .SE(test_se), 
        .CLK(n1510), .Q(\mem1[106][13] ), .QN(n26795) );
  SDFFX1 \mem1_reg[106][12]  ( .D(n15360), .SI(\mem1[106][11] ), .SE(test_se), 
        .CLK(n1510), .Q(\mem1[106][12] ), .QN(n26796) );
  SDFFX1 \mem1_reg[106][11]  ( .D(n15359), .SI(\mem1[106][10] ), .SE(test_se), 
        .CLK(n1510), .Q(\mem1[106][11] ), .QN(n26797) );
  SDFFX1 \mem1_reg[106][10]  ( .D(n15358), .SI(\mem1[106][9] ), .SE(test_se), 
        .CLK(n1510), .Q(\mem1[106][10] ), .QN(n26798) );
  SDFFX1 \mem1_reg[106][9]  ( .D(n15357), .SI(\mem1[106][8] ), .SE(test_se), 
        .CLK(n1510), .Q(\mem1[106][9] ), .QN(n26799) );
  SDFFX1 \mem1_reg[106][8]  ( .D(n15356), .SI(\mem1[105][15] ), .SE(test_se), 
        .CLK(n1510), .Q(\mem1[106][8] ), .QN(n26800) );
  SDFFX1 \mem1_reg[105][15]  ( .D(n15355), .SI(\mem1[105][14] ), .SE(test_se), 
        .CLK(n1510), .Q(\mem1[105][15] ), .QN(n26801) );
  SDFFX1 \mem1_reg[105][14]  ( .D(n15354), .SI(\mem1[105][13] ), .SE(test_se), 
        .CLK(n1510), .Q(\mem1[105][14] ), .QN(n26802) );
  SDFFX1 \mem1_reg[105][13]  ( .D(n15353), .SI(\mem1[105][12] ), .SE(test_se), 
        .CLK(n1510), .Q(\mem1[105][13] ), .QN(n26803) );
  SDFFX1 \mem1_reg[105][12]  ( .D(n15352), .SI(\mem1[105][11] ), .SE(test_se), 
        .CLK(n1510), .Q(\mem1[105][12] ), .QN(n26804) );
  SDFFX1 \mem1_reg[105][11]  ( .D(n15351), .SI(\mem1[105][10] ), .SE(test_se), 
        .CLK(n1510), .Q(\mem1[105][11] ), .QN(n26805) );
  SDFFX1 \mem1_reg[105][10]  ( .D(n15350), .SI(\mem1[105][9] ), .SE(test_se), 
        .CLK(n1510), .Q(\mem1[105][10] ), .QN(n26806) );
  SDFFX1 \mem1_reg[105][9]  ( .D(n15349), .SI(\mem1[105][8] ), .SE(test_se), 
        .CLK(n1511), .Q(\mem1[105][9] ), .QN(n26807) );
  SDFFX1 \mem1_reg[105][8]  ( .D(n15348), .SI(\mem1[104][15] ), .SE(test_se), 
        .CLK(n1511), .Q(\mem1[105][8] ), .QN(n26808) );
  SDFFX1 \mem1_reg[104][15]  ( .D(n15347), .SI(\mem1[104][14] ), .SE(test_se), 
        .CLK(n1511), .Q(\mem1[104][15] ), .QN(n26809) );
  SDFFX1 \mem1_reg[104][14]  ( .D(n15346), .SI(\mem1[104][13] ), .SE(test_se), 
        .CLK(n1511), .Q(\mem1[104][14] ), .QN(n26810) );
  SDFFX1 \mem1_reg[104][13]  ( .D(n15345), .SI(\mem1[104][12] ), .SE(test_se), 
        .CLK(n1511), .Q(\mem1[104][13] ), .QN(n26811) );
  SDFFX1 \mem1_reg[104][12]  ( .D(n15344), .SI(\mem1[104][11] ), .SE(test_se), 
        .CLK(n1511), .Q(\mem1[104][12] ), .QN(n26812) );
  SDFFX1 \mem1_reg[104][11]  ( .D(n15343), .SI(\mem1[104][10] ), .SE(test_se), 
        .CLK(n1511), .Q(\mem1[104][11] ), .QN(n26813) );
  SDFFX1 \mem1_reg[104][10]  ( .D(n15342), .SI(\mem1[104][9] ), .SE(test_se), 
        .CLK(n1511), .Q(\mem1[104][10] ), .QN(n26814) );
  SDFFX1 \mem1_reg[104][9]  ( .D(n15341), .SI(\mem1[104][8] ), .SE(test_se), 
        .CLK(n1511), .Q(\mem1[104][9] ), .QN(n26815) );
  SDFFX1 \mem1_reg[104][8]  ( .D(n15340), .SI(\mem1[103][15] ), .SE(test_se), 
        .CLK(n1511), .Q(\mem1[104][8] ), .QN(n26816) );
  SDFFX1 \mem1_reg[103][15]  ( .D(n15339), .SI(\mem1[103][14] ), .SE(test_se), 
        .CLK(n1511), .Q(\mem1[103][15] ), .QN(n26817) );
  SDFFX1 \mem1_reg[103][14]  ( .D(n15338), .SI(\mem1[103][13] ), .SE(test_se), 
        .CLK(n1511), .Q(\mem1[103][14] ), .QN(n26818) );
  SDFFX1 \mem1_reg[103][13]  ( .D(n15337), .SI(\mem1[103][12] ), .SE(test_se), 
        .CLK(n1512), .Q(\mem1[103][13] ), .QN(n26819) );
  SDFFX1 \mem1_reg[103][12]  ( .D(n15336), .SI(\mem1[103][11] ), .SE(test_se), 
        .CLK(n1512), .Q(\mem1[103][12] ), .QN(n26820) );
  SDFFX1 \mem1_reg[103][11]  ( .D(n15335), .SI(\mem1[103][10] ), .SE(test_se), 
        .CLK(n1512), .Q(\mem1[103][11] ), .QN(n26821) );
  SDFFX1 \mem1_reg[103][10]  ( .D(n15334), .SI(\mem1[103][9] ), .SE(test_se), 
        .CLK(n1512), .Q(\mem1[103][10] ), .QN(n26822) );
  SDFFX1 \mem1_reg[103][9]  ( .D(n15333), .SI(\mem1[103][8] ), .SE(test_se), 
        .CLK(n1512), .Q(\mem1[103][9] ), .QN(n26823) );
  SDFFX1 \mem1_reg[103][8]  ( .D(n15332), .SI(\mem1[102][15] ), .SE(test_se), 
        .CLK(n1512), .Q(\mem1[103][8] ), .QN(n26824) );
  SDFFX1 \mem1_reg[102][15]  ( .D(n15331), .SI(\mem1[102][14] ), .SE(test_se), 
        .CLK(n1512), .Q(\mem1[102][15] ), .QN(n26825) );
  SDFFX1 \mem1_reg[102][14]  ( .D(n15330), .SI(\mem1[102][13] ), .SE(test_se), 
        .CLK(n1512), .Q(\mem1[102][14] ), .QN(n26826) );
  SDFFX1 \mem1_reg[102][13]  ( .D(n15329), .SI(\mem1[102][12] ), .SE(test_se), 
        .CLK(n1512), .Q(\mem1[102][13] ), .QN(n26827) );
  SDFFX1 \mem1_reg[102][12]  ( .D(n15328), .SI(\mem1[102][11] ), .SE(test_se), 
        .CLK(n1512), .Q(\mem1[102][12] ), .QN(n26828) );
  SDFFX1 \mem1_reg[102][11]  ( .D(n15327), .SI(\mem1[102][10] ), .SE(test_se), 
        .CLK(n1512), .Q(\mem1[102][11] ), .QN(n26829) );
  SDFFX1 \mem1_reg[102][10]  ( .D(n15326), .SI(\mem1[102][9] ), .SE(test_se), 
        .CLK(n1512), .Q(\mem1[102][10] ), .QN(n26830) );
  SDFFX1 \mem1_reg[102][9]  ( .D(n15325), .SI(\mem1[102][8] ), .SE(test_se), 
        .CLK(n1513), .Q(\mem1[102][9] ), .QN(n26831) );
  SDFFX1 \mem1_reg[102][8]  ( .D(n15324), .SI(\mem1[101][15] ), .SE(test_se), 
        .CLK(n1513), .Q(\mem1[102][8] ), .QN(n26832) );
  SDFFX1 \mem1_reg[101][15]  ( .D(n15323), .SI(\mem1[101][14] ), .SE(test_se), 
        .CLK(n1513), .Q(\mem1[101][15] ), .QN(n26833) );
  SDFFX1 \mem1_reg[101][14]  ( .D(n15322), .SI(\mem1[101][13] ), .SE(test_se), 
        .CLK(n1513), .Q(\mem1[101][14] ), .QN(n26834) );
  SDFFX1 \mem1_reg[101][13]  ( .D(n15321), .SI(\mem1[101][12] ), .SE(test_se), 
        .CLK(n1513), .Q(\mem1[101][13] ), .QN(n26835) );
  SDFFX1 \mem1_reg[101][12]  ( .D(n15320), .SI(\mem1[101][11] ), .SE(test_se), 
        .CLK(n1513), .Q(\mem1[101][12] ), .QN(n26836) );
  SDFFX1 \mem1_reg[101][11]  ( .D(n15319), .SI(\mem1[101][10] ), .SE(test_se), 
        .CLK(n1513), .Q(\mem1[101][11] ), .QN(n26837) );
  SDFFX1 \mem1_reg[101][10]  ( .D(n15318), .SI(\mem1[101][9] ), .SE(test_se), 
        .CLK(n1513), .Q(\mem1[101][10] ), .QN(n26838) );
  SDFFX1 \mem1_reg[101][9]  ( .D(n15317), .SI(\mem1[101][8] ), .SE(test_se), 
        .CLK(n1513), .Q(\mem1[101][9] ), .QN(n26839) );
  SDFFX1 \mem1_reg[101][8]  ( .D(n15316), .SI(\mem1[100][15] ), .SE(test_se), 
        .CLK(n1513), .Q(\mem1[101][8] ), .QN(n26840) );
  SDFFX1 \mem1_reg[100][15]  ( .D(n15315), .SI(\mem1[100][14] ), .SE(test_se), 
        .CLK(n1513), .Q(\mem1[100][15] ), .QN(n26841) );
  SDFFX1 \mem1_reg[100][14]  ( .D(n15314), .SI(\mem1[100][13] ), .SE(test_se), 
        .CLK(n1513), .Q(\mem1[100][14] ), .QN(n26842) );
  SDFFX1 \mem1_reg[100][13]  ( .D(n15313), .SI(\mem1[100][12] ), .SE(test_se), 
        .CLK(n1514), .Q(\mem1[100][13] ), .QN(n26843) );
  SDFFX1 \mem1_reg[100][12]  ( .D(n15312), .SI(\mem1[100][11] ), .SE(test_se), 
        .CLK(n1514), .Q(\mem1[100][12] ), .QN(n26844) );
  SDFFX1 \mem1_reg[100][11]  ( .D(n15311), .SI(\mem1[100][10] ), .SE(test_se), 
        .CLK(n1514), .Q(\mem1[100][11] ), .QN(n26845) );
  SDFFX1 \mem1_reg[100][10]  ( .D(n15310), .SI(\mem1[100][9] ), .SE(test_se), 
        .CLK(n1514), .Q(\mem1[100][10] ), .QN(n26846) );
  SDFFX1 \mem1_reg[100][9]  ( .D(n15309), .SI(\mem1[100][8] ), .SE(test_se), 
        .CLK(n1514), .Q(\mem1[100][9] ), .QN(n26847) );
  SDFFX1 \mem1_reg[100][8]  ( .D(n15308), .SI(\mem1[99][15] ), .SE(test_se), 
        .CLK(n1514), .Q(\mem1[100][8] ), .QN(n26848) );
  SDFFX1 \mem1_reg[99][15]  ( .D(n15307), .SI(\mem1[99][14] ), .SE(test_se), 
        .CLK(n1514), .Q(\mem1[99][15] ), .QN(n26849) );
  SDFFX1 \mem1_reg[99][14]  ( .D(n15306), .SI(\mem1[99][13] ), .SE(test_se), 
        .CLK(n1514), .Q(\mem1[99][14] ), .QN(n26850) );
  SDFFX1 \mem1_reg[99][13]  ( .D(n15305), .SI(\mem1[99][12] ), .SE(test_se), 
        .CLK(n1514), .Q(\mem1[99][13] ), .QN(n26851) );
  SDFFX1 \mem1_reg[99][12]  ( .D(n15304), .SI(\mem1[99][11] ), .SE(test_se), 
        .CLK(n1514), .Q(\mem1[99][12] ), .QN(n26852) );
  SDFFX1 \mem1_reg[99][11]  ( .D(n15303), .SI(\mem1[99][10] ), .SE(test_se), 
        .CLK(n1514), .Q(\mem1[99][11] ), .QN(n26853) );
  SDFFX1 \mem1_reg[99][10]  ( .D(n15302), .SI(\mem1[99][9] ), .SE(test_se), 
        .CLK(n1514), .Q(\mem1[99][10] ), .QN(n26854) );
  SDFFX1 \mem1_reg[99][9]  ( .D(n15301), .SI(\mem1[99][8] ), .SE(test_se), 
        .CLK(n1515), .Q(\mem1[99][9] ), .QN(n26855) );
  SDFFX1 \mem1_reg[99][8]  ( .D(n15300), .SI(\mem1[98][15] ), .SE(test_se), 
        .CLK(n1515), .Q(\mem1[99][8] ), .QN(n26856) );
  SDFFX1 \mem1_reg[98][15]  ( .D(n15299), .SI(\mem1[98][14] ), .SE(test_se), 
        .CLK(n1515), .Q(\mem1[98][15] ), .QN(n26857) );
  SDFFX1 \mem1_reg[98][14]  ( .D(n15298), .SI(\mem1[98][13] ), .SE(test_se), 
        .CLK(n1515), .Q(\mem1[98][14] ), .QN(n26858) );
  SDFFX1 \mem1_reg[98][13]  ( .D(n15297), .SI(\mem1[98][12] ), .SE(test_se), 
        .CLK(n1515), .Q(\mem1[98][13] ), .QN(n26859) );
  SDFFX1 \mem1_reg[98][12]  ( .D(n15296), .SI(\mem1[98][11] ), .SE(test_se), 
        .CLK(n1515), .Q(\mem1[98][12] ), .QN(n26860) );
  SDFFX1 \mem1_reg[98][11]  ( .D(n15295), .SI(\mem1[98][10] ), .SE(test_se), 
        .CLK(n1515), .Q(\mem1[98][11] ), .QN(n26861) );
  SDFFX1 \mem1_reg[98][10]  ( .D(n15294), .SI(\mem1[98][9] ), .SE(test_se), 
        .CLK(n1515), .Q(\mem1[98][10] ), .QN(n26862) );
  SDFFX1 \mem1_reg[98][9]  ( .D(n15293), .SI(\mem1[98][8] ), .SE(test_se), 
        .CLK(n1515), .Q(\mem1[98][9] ), .QN(n26863) );
  SDFFX1 \mem1_reg[98][8]  ( .D(n15292), .SI(\mem1[97][15] ), .SE(test_se), 
        .CLK(n1515), .Q(\mem1[98][8] ), .QN(n26864) );
  SDFFX1 \mem1_reg[97][15]  ( .D(n15291), .SI(\mem1[97][14] ), .SE(test_se), 
        .CLK(n1515), .Q(\mem1[97][15] ), .QN(n26865) );
  SDFFX1 \mem1_reg[97][14]  ( .D(n15290), .SI(\mem1[97][13] ), .SE(test_se), 
        .CLK(n1515), .Q(\mem1[97][14] ), .QN(n26866) );
  SDFFX1 \mem1_reg[97][13]  ( .D(n15289), .SI(\mem1[97][12] ), .SE(test_se), 
        .CLK(n1516), .Q(\mem1[97][13] ), .QN(n26867) );
  SDFFX1 \mem1_reg[97][12]  ( .D(n15288), .SI(\mem1[97][11] ), .SE(test_se), 
        .CLK(n1516), .Q(\mem1[97][12] ), .QN(n26868) );
  SDFFX1 \mem1_reg[97][11]  ( .D(n15287), .SI(\mem1[97][10] ), .SE(test_se), 
        .CLK(n1516), .Q(\mem1[97][11] ), .QN(n26869) );
  SDFFX1 \mem1_reg[97][10]  ( .D(n15286), .SI(\mem1[97][9] ), .SE(test_se), 
        .CLK(n1516), .Q(\mem1[97][10] ), .QN(n26870) );
  SDFFX1 \mem1_reg[97][9]  ( .D(n15285), .SI(\mem1[97][8] ), .SE(test_se), 
        .CLK(n1516), .Q(\mem1[97][9] ), .QN(n26871) );
  SDFFX1 \mem1_reg[97][8]  ( .D(n15284), .SI(\mem1[96][15] ), .SE(test_se), 
        .CLK(n1516), .Q(\mem1[97][8] ), .QN(n26872) );
  SDFFX1 \mem1_reg[96][15]  ( .D(n15283), .SI(\mem1[96][14] ), .SE(test_se), 
        .CLK(n1516), .Q(\mem1[96][15] ), .QN(n26873) );
  SDFFX1 \mem1_reg[96][14]  ( .D(n15282), .SI(\mem1[96][13] ), .SE(test_se), 
        .CLK(n1516), .Q(\mem1[96][14] ), .QN(n26874) );
  SDFFX1 \mem1_reg[96][13]  ( .D(n15281), .SI(\mem1[96][12] ), .SE(test_se), 
        .CLK(n1516), .Q(\mem1[96][13] ), .QN(n26875) );
  SDFFX1 \mem1_reg[96][12]  ( .D(n15280), .SI(\mem1[96][11] ), .SE(test_se), 
        .CLK(n1516), .Q(\mem1[96][12] ), .QN(n26876) );
  SDFFX1 \mem1_reg[96][11]  ( .D(n15279), .SI(\mem1[96][10] ), .SE(test_se), 
        .CLK(n1516), .Q(\mem1[96][11] ), .QN(n26877) );
  SDFFX1 \mem1_reg[96][10]  ( .D(n15278), .SI(\mem1[96][9] ), .SE(test_se), 
        .CLK(n1516), .Q(\mem1[96][10] ), .QN(n26878) );
  SDFFX1 \mem1_reg[96][9]  ( .D(n15277), .SI(\mem1[96][8] ), .SE(test_se), 
        .CLK(n1517), .Q(\mem1[96][9] ), .QN(n26879) );
  SDFFX1 \mem1_reg[96][8]  ( .D(n15276), .SI(\mem1[95][15] ), .SE(test_se), 
        .CLK(n1517), .Q(\mem1[96][8] ), .QN(n26880) );
  SDFFX1 \mem1_reg[95][15]  ( .D(n15275), .SI(\mem1[95][14] ), .SE(test_se), 
        .CLK(n1517), .Q(\mem1[95][15] ), .QN(n26881) );
  SDFFX1 \mem1_reg[95][14]  ( .D(n15274), .SI(\mem1[95][13] ), .SE(test_se), 
        .CLK(n1517), .Q(\mem1[95][14] ), .QN(n26882) );
  SDFFX1 \mem1_reg[95][13]  ( .D(n15273), .SI(\mem1[95][12] ), .SE(test_se), 
        .CLK(n1517), .Q(\mem1[95][13] ), .QN(n26883) );
  SDFFX1 \mem1_reg[95][12]  ( .D(n15272), .SI(test_si4), .SE(test_se), .CLK(
        n1517), .Q(\mem1[95][12] ), .QN(n26884) );
  SDFFX1 \mem1_reg[95][11]  ( .D(n15271), .SI(\mem1[95][10] ), .SE(test_se), 
        .CLK(n1517), .Q(\mem1[95][11] ), .QN(n26885) );
  SDFFX1 \mem1_reg[95][10]  ( .D(n15270), .SI(\mem1[95][9] ), .SE(test_se), 
        .CLK(n1517), .Q(\mem1[95][10] ), .QN(n26886) );
  SDFFX1 \mem1_reg[95][9]  ( .D(n15269), .SI(\mem1[95][8] ), .SE(test_se), 
        .CLK(n1517), .Q(\mem1[95][9] ), .QN(n26887) );
  SDFFX1 \mem1_reg[95][8]  ( .D(n15268), .SI(\mem1[94][15] ), .SE(test_se), 
        .CLK(n1517), .Q(\mem1[95][8] ), .QN(n26888) );
  SDFFX1 \mem1_reg[94][15]  ( .D(n15267), .SI(\mem1[94][14] ), .SE(test_se), 
        .CLK(n1517), .Q(\mem1[94][15] ), .QN(n26889) );
  SDFFX1 \mem1_reg[94][14]  ( .D(n15266), .SI(\mem1[94][13] ), .SE(test_se), 
        .CLK(n1517), .Q(\mem1[94][14] ), .QN(n26890) );
  SDFFX1 \mem1_reg[94][13]  ( .D(n15265), .SI(\mem1[94][12] ), .SE(test_se), 
        .CLK(n1518), .Q(\mem1[94][13] ), .QN(n26891) );
  SDFFX1 \mem1_reg[94][12]  ( .D(n15264), .SI(\mem1[94][11] ), .SE(test_se), 
        .CLK(n1518), .Q(\mem1[94][12] ), .QN(n26892) );
  SDFFX1 \mem1_reg[94][11]  ( .D(n15263), .SI(\mem1[94][10] ), .SE(test_se), 
        .CLK(n1518), .Q(\mem1[94][11] ), .QN(n26893) );
  SDFFX1 \mem1_reg[94][10]  ( .D(n15262), .SI(\mem1[94][9] ), .SE(test_se), 
        .CLK(n1518), .Q(\mem1[94][10] ), .QN(n26894) );
  SDFFX1 \mem1_reg[94][9]  ( .D(n15261), .SI(\mem1[94][8] ), .SE(test_se), 
        .CLK(n1518), .Q(\mem1[94][9] ), .QN(n26895) );
  SDFFX1 \mem1_reg[94][8]  ( .D(n15260), .SI(\mem1[93][15] ), .SE(test_se), 
        .CLK(n1518), .Q(\mem1[94][8] ), .QN(n26896) );
  SDFFX1 \mem1_reg[93][15]  ( .D(n15259), .SI(\mem1[93][14] ), .SE(test_se), 
        .CLK(n1518), .Q(\mem1[93][15] ), .QN(n26897) );
  SDFFX1 \mem1_reg[93][14]  ( .D(n15258), .SI(\mem1[93][13] ), .SE(test_se), 
        .CLK(n1518), .Q(\mem1[93][14] ), .QN(n26898) );
  SDFFX1 \mem1_reg[93][13]  ( .D(n15257), .SI(\mem1[93][12] ), .SE(test_se), 
        .CLK(n1518), .Q(\mem1[93][13] ), .QN(n26899) );
  SDFFX1 \mem1_reg[93][12]  ( .D(n15256), .SI(\mem1[93][11] ), .SE(test_se), 
        .CLK(n1518), .Q(\mem1[93][12] ), .QN(n26900) );
  SDFFX1 \mem1_reg[93][11]  ( .D(n15255), .SI(\mem1[93][10] ), .SE(test_se), 
        .CLK(n1518), .Q(\mem1[93][11] ), .QN(n26901) );
  SDFFX1 \mem1_reg[93][10]  ( .D(n15254), .SI(\mem1[93][9] ), .SE(test_se), 
        .CLK(n1518), .Q(\mem1[93][10] ), .QN(n26902) );
  SDFFX1 \mem1_reg[93][9]  ( .D(n15253), .SI(\mem1[93][8] ), .SE(test_se), 
        .CLK(n1519), .Q(\mem1[93][9] ), .QN(n26903) );
  SDFFX1 \mem1_reg[93][8]  ( .D(n15252), .SI(\mem1[92][15] ), .SE(test_se), 
        .CLK(n1519), .Q(\mem1[93][8] ), .QN(n26904) );
  SDFFX1 \mem1_reg[92][15]  ( .D(n15251), .SI(\mem1[92][14] ), .SE(test_se), 
        .CLK(n1519), .Q(\mem1[92][15] ), .QN(n26905) );
  SDFFX1 \mem1_reg[92][14]  ( .D(n15250), .SI(\mem1[92][13] ), .SE(test_se), 
        .CLK(n1519), .Q(\mem1[92][14] ), .QN(n26906) );
  SDFFX1 \mem1_reg[92][13]  ( .D(n15249), .SI(\mem1[92][12] ), .SE(test_se), 
        .CLK(n1519), .Q(\mem1[92][13] ), .QN(n26907) );
  SDFFX1 \mem1_reg[92][12]  ( .D(n15248), .SI(\mem1[92][11] ), .SE(test_se), 
        .CLK(n1519), .Q(\mem1[92][12] ), .QN(n26908) );
  SDFFX1 \mem1_reg[92][11]  ( .D(n15247), .SI(\mem1[92][10] ), .SE(test_se), 
        .CLK(n1519), .Q(\mem1[92][11] ), .QN(n26909) );
  SDFFX1 \mem1_reg[92][10]  ( .D(n15246), .SI(\mem1[92][9] ), .SE(test_se), 
        .CLK(n1519), .Q(\mem1[92][10] ), .QN(n26910) );
  SDFFX1 \mem1_reg[92][9]  ( .D(n15245), .SI(\mem1[92][8] ), .SE(test_se), 
        .CLK(n1519), .Q(\mem1[92][9] ), .QN(n26911) );
  SDFFX1 \mem1_reg[92][8]  ( .D(n15244), .SI(\mem1[91][15] ), .SE(test_se), 
        .CLK(n1519), .Q(\mem1[92][8] ), .QN(n26912) );
  SDFFX1 \mem1_reg[91][15]  ( .D(n15243), .SI(\mem1[91][14] ), .SE(test_se), 
        .CLK(n1519), .Q(\mem1[91][15] ), .QN(n26913) );
  SDFFX1 \mem1_reg[91][14]  ( .D(n15242), .SI(\mem1[91][13] ), .SE(test_se), 
        .CLK(n1519), .Q(\mem1[91][14] ), .QN(n26914) );
  SDFFX1 \mem1_reg[91][13]  ( .D(n15241), .SI(\mem1[91][12] ), .SE(test_se), 
        .CLK(n1520), .Q(\mem1[91][13] ), .QN(n26915) );
  SDFFX1 \mem1_reg[91][12]  ( .D(n15240), .SI(\mem1[91][11] ), .SE(test_se), 
        .CLK(n1520), .Q(\mem1[91][12] ), .QN(n26916) );
  SDFFX1 \mem1_reg[91][11]  ( .D(n15239), .SI(\mem1[91][10] ), .SE(test_se), 
        .CLK(n1520), .Q(\mem1[91][11] ), .QN(n26917) );
  SDFFX1 \mem1_reg[91][10]  ( .D(n15238), .SI(\mem1[91][9] ), .SE(test_se), 
        .CLK(n1520), .Q(\mem1[91][10] ), .QN(n26918) );
  SDFFX1 \mem1_reg[91][9]  ( .D(n15237), .SI(\mem1[91][8] ), .SE(test_se), 
        .CLK(n1520), .Q(\mem1[91][9] ), .QN(n26919) );
  SDFFX1 \mem1_reg[91][8]  ( .D(n15236), .SI(\mem1[90][15] ), .SE(test_se), 
        .CLK(n1520), .Q(\mem1[91][8] ), .QN(n26920) );
  SDFFX1 \mem1_reg[90][15]  ( .D(n15235), .SI(\mem1[90][14] ), .SE(test_se), 
        .CLK(n1520), .Q(\mem1[90][15] ), .QN(n26921) );
  SDFFX1 \mem1_reg[90][14]  ( .D(n15234), .SI(\mem1[90][13] ), .SE(test_se), 
        .CLK(n1520), .Q(\mem1[90][14] ), .QN(n26922) );
  SDFFX1 \mem1_reg[90][13]  ( .D(n15233), .SI(\mem1[90][12] ), .SE(test_se), 
        .CLK(n1520), .Q(\mem1[90][13] ), .QN(n26923) );
  SDFFX1 \mem1_reg[90][12]  ( .D(n15232), .SI(\mem1[90][11] ), .SE(test_se), 
        .CLK(n1520), .Q(\mem1[90][12] ), .QN(n26924) );
  SDFFX1 \mem1_reg[90][11]  ( .D(n15231), .SI(\mem1[90][10] ), .SE(test_se), 
        .CLK(n1520), .Q(\mem1[90][11] ), .QN(n26925) );
  SDFFX1 \mem1_reg[90][10]  ( .D(n15230), .SI(\mem1[90][9] ), .SE(test_se), 
        .CLK(n1520), .Q(\mem1[90][10] ), .QN(n26926) );
  SDFFX1 \mem1_reg[90][9]  ( .D(n15229), .SI(\mem1[90][8] ), .SE(test_se), 
        .CLK(n1521), .Q(\mem1[90][9] ), .QN(n26927) );
  SDFFX1 \mem1_reg[90][8]  ( .D(n15228), .SI(\mem1[89][15] ), .SE(test_se), 
        .CLK(n1521), .Q(\mem1[90][8] ), .QN(n26928) );
  SDFFX1 \mem1_reg[89][15]  ( .D(n15227), .SI(\mem1[89][14] ), .SE(test_se), 
        .CLK(n1521), .Q(\mem1[89][15] ), .QN(n26929) );
  SDFFX1 \mem1_reg[89][14]  ( .D(n15226), .SI(\mem1[89][13] ), .SE(test_se), 
        .CLK(n1521), .Q(\mem1[89][14] ), .QN(n26930) );
  SDFFX1 \mem1_reg[89][13]  ( .D(n15225), .SI(\mem1[89][12] ), .SE(test_se), 
        .CLK(n1521), .Q(\mem1[89][13] ), .QN(n26931) );
  SDFFX1 \mem1_reg[89][12]  ( .D(n15224), .SI(\mem1[89][11] ), .SE(test_se), 
        .CLK(n1521), .Q(\mem1[89][12] ), .QN(n26932) );
  SDFFX1 \mem1_reg[89][11]  ( .D(n15223), .SI(\mem1[89][10] ), .SE(test_se), 
        .CLK(n1521), .Q(\mem1[89][11] ), .QN(n26933) );
  SDFFX1 \mem1_reg[89][10]  ( .D(n15222), .SI(\mem1[89][9] ), .SE(test_se), 
        .CLK(n1521), .Q(\mem1[89][10] ), .QN(n26934) );
  SDFFX1 \mem1_reg[89][9]  ( .D(n15221), .SI(\mem1[89][8] ), .SE(test_se), 
        .CLK(n1521), .Q(\mem1[89][9] ), .QN(n26935) );
  SDFFX1 \mem1_reg[89][8]  ( .D(n15220), .SI(\mem1[88][15] ), .SE(test_se), 
        .CLK(n1521), .Q(\mem1[89][8] ), .QN(n26936) );
  SDFFX1 \mem1_reg[88][15]  ( .D(n15219), .SI(\mem1[88][14] ), .SE(test_se), 
        .CLK(n1521), .Q(\mem1[88][15] ), .QN(n26937) );
  SDFFX1 \mem1_reg[88][14]  ( .D(n15218), .SI(\mem1[88][13] ), .SE(test_se), 
        .CLK(n1521), .Q(\mem1[88][14] ), .QN(n26938) );
  SDFFX1 \mem1_reg[88][13]  ( .D(n15217), .SI(\mem1[88][12] ), .SE(test_se), 
        .CLK(n1522), .Q(\mem1[88][13] ), .QN(n26939) );
  SDFFX1 \mem1_reg[88][12]  ( .D(n15216), .SI(\mem1[88][11] ), .SE(test_se), 
        .CLK(n1522), .Q(\mem1[88][12] ), .QN(n26940) );
  SDFFX1 \mem1_reg[88][11]  ( .D(n15215), .SI(\mem1[88][10] ), .SE(test_se), 
        .CLK(n1522), .Q(\mem1[88][11] ), .QN(n26941) );
  SDFFX1 \mem1_reg[88][10]  ( .D(n15214), .SI(\mem1[88][9] ), .SE(test_se), 
        .CLK(n1522), .Q(\mem1[88][10] ), .QN(n26942) );
  SDFFX1 \mem1_reg[88][9]  ( .D(n15213), .SI(\mem1[88][8] ), .SE(test_se), 
        .CLK(n1522), .Q(\mem1[88][9] ), .QN(n26943) );
  SDFFX1 \mem1_reg[88][8]  ( .D(n15212), .SI(\mem1[87][15] ), .SE(test_se), 
        .CLK(n1522), .Q(\mem1[88][8] ), .QN(n26944) );
  SDFFX1 \mem1_reg[87][15]  ( .D(n15211), .SI(\mem1[87][14] ), .SE(test_se), 
        .CLK(n1522), .Q(\mem1[87][15] ), .QN(n26945) );
  SDFFX1 \mem1_reg[87][14]  ( .D(n15210), .SI(\mem1[87][13] ), .SE(test_se), 
        .CLK(n1522), .Q(\mem1[87][14] ), .QN(n26946) );
  SDFFX1 \mem1_reg[87][13]  ( .D(n15209), .SI(\mem1[87][12] ), .SE(test_se), 
        .CLK(n1522), .Q(\mem1[87][13] ), .QN(n26947) );
  SDFFX1 \mem1_reg[87][12]  ( .D(n15208), .SI(\mem1[87][11] ), .SE(test_se), 
        .CLK(n1522), .Q(\mem1[87][12] ), .QN(n26948) );
  SDFFX1 \mem1_reg[87][11]  ( .D(n15207), .SI(\mem1[87][10] ), .SE(test_se), 
        .CLK(n1522), .Q(\mem1[87][11] ), .QN(n26949) );
  SDFFX1 \mem1_reg[87][10]  ( .D(n15206), .SI(\mem1[87][9] ), .SE(test_se), 
        .CLK(n1522), .Q(\mem1[87][10] ), .QN(n26950) );
  SDFFX1 \mem1_reg[87][9]  ( .D(n15205), .SI(\mem1[87][8] ), .SE(test_se), 
        .CLK(n1523), .Q(\mem1[87][9] ), .QN(n26951) );
  SDFFX1 \mem1_reg[87][8]  ( .D(n15204), .SI(\mem1[86][15] ), .SE(test_se), 
        .CLK(n1523), .Q(\mem1[87][8] ), .QN(n26952) );
  SDFFX1 \mem1_reg[86][15]  ( .D(n15203), .SI(\mem1[86][14] ), .SE(test_se), 
        .CLK(n1523), .Q(\mem1[86][15] ), .QN(n26953) );
  SDFFX1 \mem1_reg[86][14]  ( .D(n15202), .SI(\mem1[86][13] ), .SE(test_se), 
        .CLK(n1523), .Q(\mem1[86][14] ), .QN(n26954) );
  SDFFX1 \mem1_reg[86][13]  ( .D(n15201), .SI(\mem1[86][12] ), .SE(test_se), 
        .CLK(n1523), .Q(\mem1[86][13] ), .QN(n26955) );
  SDFFX1 \mem1_reg[86][12]  ( .D(n15200), .SI(\mem1[86][11] ), .SE(test_se), 
        .CLK(n1523), .Q(\mem1[86][12] ), .QN(n26956) );
  SDFFX1 \mem1_reg[86][11]  ( .D(n15199), .SI(\mem1[86][10] ), .SE(test_se), 
        .CLK(n1523), .Q(\mem1[86][11] ), .QN(n26957) );
  SDFFX1 \mem1_reg[86][10]  ( .D(n15198), .SI(\mem1[86][9] ), .SE(test_se), 
        .CLK(n1523), .Q(\mem1[86][10] ), .QN(n26958) );
  SDFFX1 \mem1_reg[86][9]  ( .D(n15197), .SI(\mem1[86][8] ), .SE(test_se), 
        .CLK(n1523), .Q(\mem1[86][9] ), .QN(n26959) );
  SDFFX1 \mem1_reg[86][8]  ( .D(n15196), .SI(\mem1[85][15] ), .SE(test_se), 
        .CLK(n1523), .Q(\mem1[86][8] ), .QN(n26960) );
  SDFFX1 \mem1_reg[85][15]  ( .D(n15195), .SI(\mem1[85][14] ), .SE(test_se), 
        .CLK(n1523), .Q(\mem1[85][15] ), .QN(n26961) );
  SDFFX1 \mem1_reg[85][14]  ( .D(n15194), .SI(\mem1[85][13] ), .SE(test_se), 
        .CLK(n1523), .Q(\mem1[85][14] ), .QN(n26962) );
  SDFFX1 \mem1_reg[85][13]  ( .D(n15193), .SI(\mem1[85][12] ), .SE(test_se), 
        .CLK(n1524), .Q(\mem1[85][13] ), .QN(n26963) );
  SDFFX1 \mem1_reg[85][12]  ( .D(n15192), .SI(\mem1[85][11] ), .SE(test_se), 
        .CLK(n1524), .Q(\mem1[85][12] ), .QN(n26964) );
  SDFFX1 \mem1_reg[85][11]  ( .D(n15191), .SI(\mem1[85][10] ), .SE(test_se), 
        .CLK(n1524), .Q(\mem1[85][11] ), .QN(n26965) );
  SDFFX1 \mem1_reg[85][10]  ( .D(n15190), .SI(\mem1[85][9] ), .SE(test_se), 
        .CLK(n1524), .Q(\mem1[85][10] ), .QN(n26966) );
  SDFFX1 \mem1_reg[85][9]  ( .D(n15189), .SI(\mem1[85][8] ), .SE(test_se), 
        .CLK(n1524), .Q(\mem1[85][9] ), .QN(n26967) );
  SDFFX1 \mem1_reg[85][8]  ( .D(n15188), .SI(\mem1[84][15] ), .SE(test_se), 
        .CLK(n1524), .Q(\mem1[85][8] ), .QN(n26968) );
  SDFFX1 \mem1_reg[84][15]  ( .D(n15187), .SI(\mem1[84][14] ), .SE(test_se), 
        .CLK(n1524), .Q(\mem1[84][15] ), .QN(n26969) );
  SDFFX1 \mem1_reg[84][14]  ( .D(n15186), .SI(\mem1[84][13] ), .SE(test_se), 
        .CLK(n1524), .Q(\mem1[84][14] ), .QN(n26970) );
  SDFFX1 \mem1_reg[84][13]  ( .D(n15185), .SI(\mem1[84][12] ), .SE(test_se), 
        .CLK(n1524), .Q(\mem1[84][13] ), .QN(n26971) );
  SDFFX1 \mem1_reg[84][12]  ( .D(n15184), .SI(\mem1[84][11] ), .SE(test_se), 
        .CLK(n1524), .Q(\mem1[84][12] ), .QN(n26972) );
  SDFFX1 \mem1_reg[84][11]  ( .D(n15183), .SI(\mem1[84][10] ), .SE(test_se), 
        .CLK(n1524), .Q(\mem1[84][11] ), .QN(n26973) );
  SDFFX1 \mem1_reg[84][10]  ( .D(n15182), .SI(\mem1[84][9] ), .SE(test_se), 
        .CLK(n1524), .Q(\mem1[84][10] ), .QN(n26974) );
  SDFFX1 \mem1_reg[84][9]  ( .D(n15181), .SI(\mem1[84][8] ), .SE(test_se), 
        .CLK(n1525), .Q(\mem1[84][9] ), .QN(n26975) );
  SDFFX1 \mem1_reg[84][8]  ( .D(n15180), .SI(\mem1[83][15] ), .SE(test_se), 
        .CLK(n1525), .Q(\mem1[84][8] ), .QN(n26976) );
  SDFFX1 \mem1_reg[83][15]  ( .D(n15179), .SI(\mem1[83][14] ), .SE(test_se), 
        .CLK(n1525), .Q(\mem1[83][15] ), .QN(n26977) );
  SDFFX1 \mem1_reg[83][14]  ( .D(n15178), .SI(\mem1[83][13] ), .SE(test_se), 
        .CLK(n1525), .Q(\mem1[83][14] ), .QN(n26978) );
  SDFFX1 \mem1_reg[83][13]  ( .D(n15177), .SI(\mem1[83][12] ), .SE(test_se), 
        .CLK(n1525), .Q(\mem1[83][13] ), .QN(n26979) );
  SDFFX1 \mem1_reg[83][12]  ( .D(n15176), .SI(\mem1[83][11] ), .SE(test_se), 
        .CLK(n1525), .Q(\mem1[83][12] ), .QN(n26980) );
  SDFFX1 \mem1_reg[83][11]  ( .D(n15175), .SI(\mem1[83][10] ), .SE(test_se), 
        .CLK(n1525), .Q(\mem1[83][11] ), .QN(n26981) );
  SDFFX1 \mem1_reg[83][10]  ( .D(n15174), .SI(\mem1[83][9] ), .SE(test_se), 
        .CLK(n1525), .Q(\mem1[83][10] ), .QN(n26982) );
  SDFFX1 \mem1_reg[83][9]  ( .D(n15173), .SI(\mem1[83][8] ), .SE(test_se), 
        .CLK(n1525), .Q(\mem1[83][9] ), .QN(n26983) );
  SDFFX1 \mem1_reg[83][8]  ( .D(n15172), .SI(\mem1[82][15] ), .SE(test_se), 
        .CLK(n1525), .Q(\mem1[83][8] ), .QN(n26984) );
  SDFFX1 \mem1_reg[82][15]  ( .D(n15171), .SI(\mem1[82][14] ), .SE(test_se), 
        .CLK(n1525), .Q(\mem1[82][15] ), .QN(n26985) );
  SDFFX1 \mem1_reg[82][14]  ( .D(n15170), .SI(\mem1[82][13] ), .SE(test_se), 
        .CLK(n1525), .Q(\mem1[82][14] ), .QN(n26986) );
  SDFFX1 \mem1_reg[82][13]  ( .D(n15169), .SI(\mem1[82][12] ), .SE(test_se), 
        .CLK(n1526), .Q(\mem1[82][13] ), .QN(n26987) );
  SDFFX1 \mem1_reg[82][12]  ( .D(n15168), .SI(\mem1[82][11] ), .SE(test_se), 
        .CLK(n1526), .Q(\mem1[82][12] ), .QN(n26988) );
  SDFFX1 \mem1_reg[82][11]  ( .D(n15167), .SI(\mem1[82][10] ), .SE(test_se), 
        .CLK(n1526), .Q(\mem1[82][11] ), .QN(n26989) );
  SDFFX1 \mem1_reg[82][10]  ( .D(n15166), .SI(\mem1[82][9] ), .SE(test_se), 
        .CLK(n1526), .Q(\mem1[82][10] ), .QN(n26990) );
  SDFFX1 \mem1_reg[82][9]  ( .D(n15165), .SI(\mem1[82][8] ), .SE(test_se), 
        .CLK(n1526), .Q(\mem1[82][9] ), .QN(n26991) );
  SDFFX1 \mem1_reg[82][8]  ( .D(n15164), .SI(\mem1[81][15] ), .SE(test_se), 
        .CLK(n1526), .Q(\mem1[82][8] ), .QN(n26992) );
  SDFFX1 \mem1_reg[81][15]  ( .D(n15163), .SI(\mem1[81][14] ), .SE(test_se), 
        .CLK(n1526), .Q(\mem1[81][15] ), .QN(n26993) );
  SDFFX1 \mem1_reg[81][14]  ( .D(n15162), .SI(\mem1[81][13] ), .SE(test_se), 
        .CLK(n1526), .Q(\mem1[81][14] ), .QN(n26994) );
  SDFFX1 \mem1_reg[81][13]  ( .D(n15161), .SI(\mem1[81][12] ), .SE(test_se), 
        .CLK(n1526), .Q(\mem1[81][13] ), .QN(n26995) );
  SDFFX1 \mem1_reg[81][12]  ( .D(n15160), .SI(\mem1[81][11] ), .SE(test_se), 
        .CLK(n1526), .Q(\mem1[81][12] ), .QN(n26996) );
  SDFFX1 \mem1_reg[81][11]  ( .D(n15159), .SI(\mem1[81][10] ), .SE(test_se), 
        .CLK(n1526), .Q(\mem1[81][11] ), .QN(n26997) );
  SDFFX1 \mem1_reg[81][10]  ( .D(n15158), .SI(\mem1[81][9] ), .SE(test_se), 
        .CLK(n1526), .Q(\mem1[81][10] ), .QN(n26998) );
  SDFFX1 \mem1_reg[81][9]  ( .D(n15157), .SI(\mem1[81][8] ), .SE(test_se), 
        .CLK(n1527), .Q(\mem1[81][9] ), .QN(n26999) );
  SDFFX1 \mem1_reg[81][8]  ( .D(n15156), .SI(\mem1[80][15] ), .SE(test_se), 
        .CLK(n1527), .Q(\mem1[81][8] ), .QN(n27000) );
  SDFFX1 \mem1_reg[80][15]  ( .D(n15155), .SI(\mem1[80][14] ), .SE(test_se), 
        .CLK(n1527), .Q(\mem1[80][15] ), .QN(n27001) );
  SDFFX1 \mem1_reg[80][14]  ( .D(n15154), .SI(\mem1[80][13] ), .SE(test_se), 
        .CLK(n1527), .Q(\mem1[80][14] ), .QN(n27002) );
  SDFFX1 \mem1_reg[80][13]  ( .D(n15153), .SI(\mem1[80][12] ), .SE(test_se), 
        .CLK(n1527), .Q(\mem1[80][13] ), .QN(n27003) );
  SDFFX1 \mem1_reg[80][12]  ( .D(n15152), .SI(\mem1[80][11] ), .SE(test_se), 
        .CLK(n1527), .Q(\mem1[80][12] ), .QN(n27004) );
  SDFFX1 \mem1_reg[80][11]  ( .D(n15151), .SI(\mem1[80][10] ), .SE(test_se), 
        .CLK(n1527), .Q(\mem1[80][11] ), .QN(n27005) );
  SDFFX1 \mem1_reg[80][10]  ( .D(n15150), .SI(\mem1[80][9] ), .SE(test_se), 
        .CLK(n1527), .Q(\mem1[80][10] ), .QN(n27006) );
  SDFFX1 \mem1_reg[80][9]  ( .D(n15149), .SI(\mem1[80][8] ), .SE(test_se), 
        .CLK(n1527), .Q(\mem1[80][9] ), .QN(n27007) );
  SDFFX1 \mem1_reg[80][8]  ( .D(n15148), .SI(\mem1[79][15] ), .SE(test_se), 
        .CLK(n1527), .Q(\mem1[80][8] ), .QN(n27008) );
  SDFFX1 \mem1_reg[79][15]  ( .D(n15147), .SI(\mem1[79][14] ), .SE(test_se), 
        .CLK(n1527), .Q(\mem1[79][15] ), .QN(n27009) );
  SDFFX1 \mem1_reg[79][14]  ( .D(n15146), .SI(\mem1[79][13] ), .SE(test_se), 
        .CLK(n1527), .Q(\mem1[79][14] ), .QN(n27010) );
  SDFFX1 \mem1_reg[79][13]  ( .D(n15145), .SI(\mem1[79][12] ), .SE(test_se), 
        .CLK(n1528), .Q(\mem1[79][13] ), .QN(n27011) );
  SDFFX1 \mem1_reg[79][12]  ( .D(n15144), .SI(\mem1[79][11] ), .SE(test_se), 
        .CLK(n1528), .Q(\mem1[79][12] ), .QN(n27012) );
  SDFFX1 \mem1_reg[79][11]  ( .D(n15143), .SI(\mem1[79][10] ), .SE(test_se), 
        .CLK(n1528), .Q(\mem1[79][11] ), .QN(n27013) );
  SDFFX1 \mem1_reg[79][10]  ( .D(n15142), .SI(\mem1[79][9] ), .SE(test_se), 
        .CLK(n1528), .Q(\mem1[79][10] ), .QN(n27014) );
  SDFFX1 \mem1_reg[79][9]  ( .D(n15141), .SI(\mem1[79][8] ), .SE(test_se), 
        .CLK(n1528), .Q(\mem1[79][9] ), .QN(n27015) );
  SDFFX1 \mem1_reg[79][8]  ( .D(n15140), .SI(\mem1[78][15] ), .SE(test_se), 
        .CLK(n1528), .Q(\mem1[79][8] ), .QN(n27016) );
  SDFFX1 \mem1_reg[78][15]  ( .D(n15139), .SI(\mem1[78][14] ), .SE(test_se), 
        .CLK(n1528), .Q(\mem1[78][15] ), .QN(n27017) );
  SDFFX1 \mem1_reg[78][14]  ( .D(n15138), .SI(\mem1[78][13] ), .SE(test_se), 
        .CLK(n1528), .Q(\mem1[78][14] ), .QN(n27018) );
  SDFFX1 \mem1_reg[78][13]  ( .D(n15137), .SI(\mem1[78][12] ), .SE(test_se), 
        .CLK(n1528), .Q(\mem1[78][13] ), .QN(n27019) );
  SDFFX1 \mem1_reg[78][12]  ( .D(n15136), .SI(\mem1[78][11] ), .SE(test_se), 
        .CLK(n1528), .Q(\mem1[78][12] ), .QN(n27020) );
  SDFFX1 \mem1_reg[78][11]  ( .D(n15135), .SI(\mem1[78][10] ), .SE(test_se), 
        .CLK(n1528), .Q(\mem1[78][11] ), .QN(n27021) );
  SDFFX1 \mem1_reg[78][10]  ( .D(n15134), .SI(\mem1[78][9] ), .SE(test_se), 
        .CLK(n1528), .Q(\mem1[78][10] ), .QN(n27022) );
  SDFFX1 \mem1_reg[78][9]  ( .D(n15133), .SI(\mem1[78][8] ), .SE(test_se), 
        .CLK(n1529), .Q(\mem1[78][9] ), .QN(n27023) );
  SDFFX1 \mem1_reg[78][8]  ( .D(n15132), .SI(\mem1[77][15] ), .SE(test_se), 
        .CLK(n1529), .Q(\mem1[78][8] ), .QN(n27024) );
  SDFFX1 \mem1_reg[77][15]  ( .D(n15131), .SI(\mem1[77][14] ), .SE(test_se), 
        .CLK(n1529), .Q(\mem1[77][15] ), .QN(n27025) );
  SDFFX1 \mem1_reg[77][14]  ( .D(n15130), .SI(\mem1[77][13] ), .SE(test_se), 
        .CLK(n1529), .Q(\mem1[77][14] ), .QN(n27026) );
  SDFFX1 \mem1_reg[77][13]  ( .D(n15129), .SI(\mem1[77][12] ), .SE(test_se), 
        .CLK(n1529), .Q(\mem1[77][13] ), .QN(n27027) );
  SDFFX1 \mem1_reg[77][12]  ( .D(n15128), .SI(\mem1[77][11] ), .SE(test_se), 
        .CLK(n1529), .Q(\mem1[77][12] ), .QN(n27028) );
  SDFFX1 \mem1_reg[77][11]  ( .D(n15127), .SI(\mem1[77][10] ), .SE(test_se), 
        .CLK(n1529), .Q(\mem1[77][11] ), .QN(n27029) );
  SDFFX1 \mem1_reg[77][10]  ( .D(n15126), .SI(\mem1[77][9] ), .SE(test_se), 
        .CLK(n1529), .Q(\mem1[77][10] ), .QN(n27030) );
  SDFFX1 \mem1_reg[77][9]  ( .D(n15125), .SI(\mem1[77][8] ), .SE(test_se), 
        .CLK(n1529), .Q(\mem1[77][9] ), .QN(n27031) );
  SDFFX1 \mem1_reg[77][8]  ( .D(n15124), .SI(\mem1[76][15] ), .SE(test_se), 
        .CLK(n1529), .Q(\mem1[77][8] ), .QN(n27032) );
  SDFFX1 \mem1_reg[76][15]  ( .D(n15123), .SI(\mem1[76][14] ), .SE(test_se), 
        .CLK(n1529), .Q(\mem1[76][15] ), .QN(n27033) );
  SDFFX1 \mem1_reg[76][14]  ( .D(n15122), .SI(\mem1[76][13] ), .SE(test_se), 
        .CLK(n1529), .Q(\mem1[76][14] ), .QN(n27034) );
  SDFFX1 \mem1_reg[76][13]  ( .D(n15121), .SI(\mem1[76][12] ), .SE(test_se), 
        .CLK(n1530), .Q(\mem1[76][13] ), .QN(n27035) );
  SDFFX1 \mem1_reg[76][12]  ( .D(n15120), .SI(\mem1[76][11] ), .SE(test_se), 
        .CLK(n1530), .Q(\mem1[76][12] ), .QN(n27036) );
  SDFFX1 \mem1_reg[76][11]  ( .D(n15119), .SI(\mem1[76][10] ), .SE(test_se), 
        .CLK(n1530), .Q(\mem1[76][11] ), .QN(n27037) );
  SDFFX1 \mem1_reg[76][10]  ( .D(n15118), .SI(\mem1[76][9] ), .SE(test_se), 
        .CLK(n1530), .Q(\mem1[76][10] ), .QN(n27038) );
  SDFFX1 \mem1_reg[76][9]  ( .D(n15117), .SI(\mem1[76][8] ), .SE(test_se), 
        .CLK(n1530), .Q(\mem1[76][9] ), .QN(n27039) );
  SDFFX1 \mem1_reg[76][8]  ( .D(n15116), .SI(\mem1[75][15] ), .SE(test_se), 
        .CLK(n1530), .Q(\mem1[76][8] ), .QN(n27040) );
  SDFFX1 \mem1_reg[75][15]  ( .D(n15115), .SI(\mem1[75][14] ), .SE(test_se), 
        .CLK(n1530), .Q(\mem1[75][15] ), .QN(n27041) );
  SDFFX1 \mem1_reg[75][14]  ( .D(n15114), .SI(\mem1[75][13] ), .SE(test_se), 
        .CLK(n1530), .Q(\mem1[75][14] ), .QN(n27042) );
  SDFFX1 \mem1_reg[75][13]  ( .D(n15113), .SI(\mem1[75][12] ), .SE(test_se), 
        .CLK(n1530), .Q(\mem1[75][13] ), .QN(n27043) );
  SDFFX1 \mem1_reg[75][12]  ( .D(n15112), .SI(\mem1[75][11] ), .SE(test_se), 
        .CLK(n1530), .Q(\mem1[75][12] ), .QN(n27044) );
  SDFFX1 \mem1_reg[75][11]  ( .D(n15111), .SI(\mem1[75][10] ), .SE(test_se), 
        .CLK(n1530), .Q(\mem1[75][11] ), .QN(n27045) );
  SDFFX1 \mem1_reg[75][10]  ( .D(n15110), .SI(\mem1[75][9] ), .SE(test_se), 
        .CLK(n1530), .Q(\mem1[75][10] ), .QN(n27046) );
  SDFFX1 \mem1_reg[75][9]  ( .D(n15109), .SI(\mem1[75][8] ), .SE(test_se), 
        .CLK(n1531), .Q(\mem1[75][9] ), .QN(n27047) );
  SDFFX1 \mem1_reg[75][8]  ( .D(n15108), .SI(\mem1[74][15] ), .SE(test_se), 
        .CLK(n1531), .Q(\mem1[75][8] ), .QN(n27048) );
  SDFFX1 \mem1_reg[74][15]  ( .D(n15107), .SI(\mem1[74][14] ), .SE(test_se), 
        .CLK(n1531), .Q(\mem1[74][15] ), .QN(n27049) );
  SDFFX1 \mem1_reg[74][14]  ( .D(n15106), .SI(\mem1[74][13] ), .SE(test_se), 
        .CLK(n1531), .Q(\mem1[74][14] ), .QN(n27050) );
  SDFFX1 \mem1_reg[74][13]  ( .D(n15105), .SI(\mem1[74][12] ), .SE(test_se), 
        .CLK(n1531), .Q(\mem1[74][13] ), .QN(n27051) );
  SDFFX1 \mem1_reg[74][12]  ( .D(n15104), .SI(\mem1[74][11] ), .SE(test_se), 
        .CLK(n1531), .Q(\mem1[74][12] ), .QN(n27052) );
  SDFFX1 \mem1_reg[74][11]  ( .D(n15103), .SI(\mem1[74][10] ), .SE(test_se), 
        .CLK(n1531), .Q(\mem1[74][11] ), .QN(n27053) );
  SDFFX1 \mem1_reg[74][10]  ( .D(n15102), .SI(\mem1[74][9] ), .SE(test_se), 
        .CLK(n1531), .Q(\mem1[74][10] ), .QN(n27054) );
  SDFFX1 \mem1_reg[74][9]  ( .D(n15101), .SI(\mem1[74][8] ), .SE(test_se), 
        .CLK(n1531), .Q(\mem1[74][9] ), .QN(n27055) );
  SDFFX1 \mem1_reg[74][8]  ( .D(n15100), .SI(\mem1[73][15] ), .SE(test_se), 
        .CLK(n1531), .Q(\mem1[74][8] ), .QN(n27056) );
  SDFFX1 \mem1_reg[73][15]  ( .D(n15099), .SI(\mem1[73][14] ), .SE(test_se), 
        .CLK(n1531), .Q(\mem1[73][15] ), .QN(n27057) );
  SDFFX1 \mem1_reg[73][14]  ( .D(n15098), .SI(\mem1[73][13] ), .SE(test_se), 
        .CLK(n1531), .Q(\mem1[73][14] ), .QN(n27058) );
  SDFFX1 \mem1_reg[73][13]  ( .D(n15097), .SI(\mem1[73][12] ), .SE(test_se), 
        .CLK(n1532), .Q(\mem1[73][13] ), .QN(n27059) );
  SDFFX1 \mem1_reg[73][12]  ( .D(n15096), .SI(\mem1[73][11] ), .SE(test_se), 
        .CLK(n1532), .Q(\mem1[73][12] ), .QN(n27060) );
  SDFFX1 \mem1_reg[73][11]  ( .D(n15095), .SI(\mem1[73][10] ), .SE(test_se), 
        .CLK(n1532), .Q(\mem1[73][11] ), .QN(n27061) );
  SDFFX1 \mem1_reg[73][10]  ( .D(n15094), .SI(\mem1[73][9] ), .SE(test_se), 
        .CLK(n1532), .Q(\mem1[73][10] ), .QN(n27062) );
  SDFFX1 \mem1_reg[73][9]  ( .D(n15093), .SI(\mem1[73][8] ), .SE(test_se), 
        .CLK(n1532), .Q(\mem1[73][9] ), .QN(n27063) );
  SDFFX1 \mem1_reg[73][8]  ( .D(n15092), .SI(\mem1[72][15] ), .SE(test_se), 
        .CLK(n1532), .Q(\mem1[73][8] ), .QN(n27064) );
  SDFFX1 \mem1_reg[72][15]  ( .D(n15091), .SI(\mem1[72][14] ), .SE(test_se), 
        .CLK(n1532), .Q(\mem1[72][15] ), .QN(n27065) );
  SDFFX1 \mem1_reg[72][14]  ( .D(n15090), .SI(\mem1[72][13] ), .SE(test_se), 
        .CLK(n1532), .Q(\mem1[72][14] ), .QN(n27066) );
  SDFFX1 \mem1_reg[72][13]  ( .D(n15089), .SI(\mem1[72][12] ), .SE(test_se), 
        .CLK(n1532), .Q(\mem1[72][13] ), .QN(n27067) );
  SDFFX1 \mem1_reg[72][12]  ( .D(n15088), .SI(\mem1[72][11] ), .SE(test_se), 
        .CLK(n1532), .Q(\mem1[72][12] ), .QN(n27068) );
  SDFFX1 \mem1_reg[72][11]  ( .D(n15087), .SI(\mem1[72][10] ), .SE(test_se), 
        .CLK(n1532), .Q(\mem1[72][11] ), .QN(n27069) );
  SDFFX1 \mem1_reg[72][10]  ( .D(n15086), .SI(\mem1[72][9] ), .SE(test_se), 
        .CLK(n1532), .Q(\mem1[72][10] ), .QN(n27070) );
  SDFFX1 \mem1_reg[72][9]  ( .D(n15085), .SI(\mem1[72][8] ), .SE(test_se), 
        .CLK(n1533), .Q(\mem1[72][9] ), .QN(n27071) );
  SDFFX1 \mem1_reg[72][8]  ( .D(n15084), .SI(\mem1[71][15] ), .SE(test_se), 
        .CLK(n1533), .Q(\mem1[72][8] ), .QN(n27072) );
  SDFFX1 \mem1_reg[71][15]  ( .D(n15083), .SI(\mem1[71][14] ), .SE(test_se), 
        .CLK(n1533), .Q(\mem1[71][15] ), .QN(n27073) );
  SDFFX1 \mem1_reg[71][14]  ( .D(n15082), .SI(\mem1[71][13] ), .SE(test_se), 
        .CLK(n1533), .Q(\mem1[71][14] ), .QN(n27074) );
  SDFFX1 \mem1_reg[71][13]  ( .D(n15081), .SI(\mem1[71][12] ), .SE(test_se), 
        .CLK(n1533), .Q(\mem1[71][13] ), .QN(n27075) );
  SDFFX1 \mem1_reg[71][12]  ( .D(n15080), .SI(\mem1[71][11] ), .SE(test_se), 
        .CLK(n1533), .Q(\mem1[71][12] ), .QN(n27076) );
  SDFFX1 \mem1_reg[71][11]  ( .D(n15079), .SI(\mem1[71][10] ), .SE(test_se), 
        .CLK(n1533), .Q(\mem1[71][11] ), .QN(n27077) );
  SDFFX1 \mem1_reg[71][10]  ( .D(n15078), .SI(\mem1[71][9] ), .SE(test_se), 
        .CLK(n1533), .Q(\mem1[71][10] ), .QN(n27078) );
  SDFFX1 \mem1_reg[71][9]  ( .D(n15077), .SI(\mem1[71][8] ), .SE(test_se), 
        .CLK(n1533), .Q(\mem1[71][9] ), .QN(n27079) );
  SDFFX1 \mem1_reg[71][8]  ( .D(n15076), .SI(\mem1[70][15] ), .SE(test_se), 
        .CLK(n1533), .Q(\mem1[71][8] ), .QN(n27080) );
  SDFFX1 \mem1_reg[70][15]  ( .D(n15075), .SI(\mem1[70][14] ), .SE(test_se), 
        .CLK(n1533), .Q(\mem1[70][15] ), .QN(n27081) );
  SDFFX1 \mem1_reg[70][14]  ( .D(n15074), .SI(\mem1[70][13] ), .SE(test_se), 
        .CLK(n1533), .Q(\mem1[70][14] ), .QN(n27082) );
  SDFFX1 \mem1_reg[70][13]  ( .D(n15073), .SI(\mem1[70][12] ), .SE(test_se), 
        .CLK(n1534), .Q(\mem1[70][13] ), .QN(n27083) );
  SDFFX1 \mem1_reg[70][12]  ( .D(n15072), .SI(\mem1[70][11] ), .SE(test_se), 
        .CLK(n1534), .Q(\mem1[70][12] ), .QN(n27084) );
  SDFFX1 \mem1_reg[70][11]  ( .D(n15071), .SI(\mem1[70][10] ), .SE(test_se), 
        .CLK(n1534), .Q(\mem1[70][11] ), .QN(n27085) );
  SDFFX1 \mem1_reg[70][10]  ( .D(n15070), .SI(\mem1[70][9] ), .SE(test_se), 
        .CLK(n1534), .Q(\mem1[70][10] ), .QN(n27086) );
  SDFFX1 \mem1_reg[70][9]  ( .D(n15069), .SI(\mem1[70][8] ), .SE(test_se), 
        .CLK(n1534), .Q(\mem1[70][9] ), .QN(n27087) );
  SDFFX1 \mem1_reg[70][8]  ( .D(n15068), .SI(\mem1[69][15] ), .SE(test_se), 
        .CLK(n1534), .Q(\mem1[70][8] ), .QN(n27088) );
  SDFFX1 \mem1_reg[69][15]  ( .D(n15067), .SI(\mem1[69][14] ), .SE(test_se), 
        .CLK(n1534), .Q(\mem1[69][15] ), .QN(n27089) );
  SDFFX1 \mem1_reg[69][14]  ( .D(n15066), .SI(\mem1[69][13] ), .SE(test_se), 
        .CLK(n1534), .Q(\mem1[69][14] ), .QN(n27090) );
  SDFFX1 \mem1_reg[69][13]  ( .D(n15065), .SI(\mem1[69][12] ), .SE(test_se), 
        .CLK(n1534), .Q(\mem1[69][13] ), .QN(n27091) );
  SDFFX1 \mem1_reg[69][12]  ( .D(n15064), .SI(\mem1[69][11] ), .SE(test_se), 
        .CLK(n1534), .Q(\mem1[69][12] ), .QN(n27092) );
  SDFFX1 \mem1_reg[69][11]  ( .D(n15063), .SI(\mem1[69][10] ), .SE(test_se), 
        .CLK(n1534), .Q(\mem1[69][11] ), .QN(n27093) );
  SDFFX1 \mem1_reg[69][10]  ( .D(n15062), .SI(\mem1[69][9] ), .SE(test_se), 
        .CLK(n1534), .Q(\mem1[69][10] ), .QN(n27094) );
  SDFFX1 \mem1_reg[69][9]  ( .D(n15061), .SI(\mem1[69][8] ), .SE(test_se), 
        .CLK(n1535), .Q(\mem1[69][9] ), .QN(n27095) );
  SDFFX1 \mem1_reg[69][8]  ( .D(n15060), .SI(\mem1[68][15] ), .SE(test_se), 
        .CLK(n1535), .Q(\mem1[69][8] ), .QN(n27096) );
  SDFFX1 \mem1_reg[68][15]  ( .D(n15059), .SI(\mem1[68][14] ), .SE(test_se), 
        .CLK(n1535), .Q(\mem1[68][15] ), .QN(n27097) );
  SDFFX1 \mem1_reg[68][14]  ( .D(n15058), .SI(\mem1[68][13] ), .SE(test_se), 
        .CLK(n1535), .Q(\mem1[68][14] ), .QN(n27098) );
  SDFFX1 \mem1_reg[68][13]  ( .D(n15057), .SI(\mem1[68][12] ), .SE(test_se), 
        .CLK(n1535), .Q(\mem1[68][13] ), .QN(n27099) );
  SDFFX1 \mem1_reg[68][12]  ( .D(n15056), .SI(\mem1[68][11] ), .SE(test_se), 
        .CLK(n1535), .Q(\mem1[68][12] ), .QN(n27100) );
  SDFFX1 \mem1_reg[68][11]  ( .D(n15055), .SI(\mem1[68][10] ), .SE(test_se), 
        .CLK(n1535), .Q(\mem1[68][11] ), .QN(n27101) );
  SDFFX1 \mem1_reg[68][10]  ( .D(n15054), .SI(\mem1[68][9] ), .SE(test_se), 
        .CLK(n1535), .Q(\mem1[68][10] ), .QN(n27102) );
  SDFFX1 \mem1_reg[68][9]  ( .D(n15053), .SI(\mem1[68][8] ), .SE(test_se), 
        .CLK(n1535), .Q(\mem1[68][9] ), .QN(n27103) );
  SDFFX1 \mem1_reg[68][8]  ( .D(n15052), .SI(\mem1[67][15] ), .SE(test_se), 
        .CLK(n1535), .Q(\mem1[68][8] ), .QN(n27104) );
  SDFFX1 \mem1_reg[67][15]  ( .D(n15051), .SI(\mem1[67][14] ), .SE(test_se), 
        .CLK(n1535), .Q(\mem1[67][15] ), .QN(n27105) );
  SDFFX1 \mem1_reg[67][14]  ( .D(n15050), .SI(\mem1[67][13] ), .SE(test_se), 
        .CLK(n1535), .Q(\mem1[67][14] ), .QN(n27106) );
  SDFFX1 \mem1_reg[67][13]  ( .D(n15049), .SI(\mem1[67][12] ), .SE(test_se), 
        .CLK(n1536), .Q(\mem1[67][13] ), .QN(n27107) );
  SDFFX1 \mem1_reg[67][12]  ( .D(n15048), .SI(\mem1[67][11] ), .SE(test_se), 
        .CLK(n1536), .Q(\mem1[67][12] ), .QN(n27108) );
  SDFFX1 \mem1_reg[67][11]  ( .D(n15047), .SI(\mem1[67][10] ), .SE(test_se), 
        .CLK(n1536), .Q(\mem1[67][11] ), .QN(n27109) );
  SDFFX1 \mem1_reg[67][10]  ( .D(n15046), .SI(\mem1[67][9] ), .SE(test_se), 
        .CLK(n1536), .Q(\mem1[67][10] ), .QN(n27110) );
  SDFFX1 \mem1_reg[67][9]  ( .D(n15045), .SI(\mem1[67][8] ), .SE(test_se), 
        .CLK(n1536), .Q(\mem1[67][9] ), .QN(n27111) );
  SDFFX1 \mem1_reg[67][8]  ( .D(n15044), .SI(\mem1[66][15] ), .SE(test_se), 
        .CLK(n1536), .Q(\mem1[67][8] ), .QN(n27112) );
  SDFFX1 \mem1_reg[66][15]  ( .D(n15043), .SI(\mem1[66][14] ), .SE(test_se), 
        .CLK(n1536), .Q(\mem1[66][15] ), .QN(n27113) );
  SDFFX1 \mem1_reg[66][14]  ( .D(n15042), .SI(\mem1[66][13] ), .SE(test_se), 
        .CLK(n1536), .Q(\mem1[66][14] ), .QN(n27114) );
  SDFFX1 \mem1_reg[66][13]  ( .D(n15041), .SI(\mem1[66][12] ), .SE(test_se), 
        .CLK(n1536), .Q(\mem1[66][13] ), .QN(n27115) );
  SDFFX1 \mem1_reg[66][12]  ( .D(n15040), .SI(\mem1[66][11] ), .SE(test_se), 
        .CLK(n1536), .Q(\mem1[66][12] ), .QN(n27116) );
  SDFFX1 \mem1_reg[66][11]  ( .D(n15039), .SI(\mem1[66][10] ), .SE(test_se), 
        .CLK(n1536), .Q(\mem1[66][11] ), .QN(n27117) );
  SDFFX1 \mem1_reg[66][10]  ( .D(n15038), .SI(\mem1[66][9] ), .SE(test_se), 
        .CLK(n1536), .Q(\mem1[66][10] ), .QN(n27118) );
  SDFFX1 \mem1_reg[66][9]  ( .D(n15037), .SI(\mem1[66][8] ), .SE(test_se), 
        .CLK(n1537), .Q(\mem1[66][9] ), .QN(n27119) );
  SDFFX1 \mem1_reg[66][8]  ( .D(n15036), .SI(\mem1[65][15] ), .SE(test_se), 
        .CLK(n1537), .Q(\mem1[66][8] ), .QN(n27120) );
  SDFFX1 \mem1_reg[65][15]  ( .D(n15035), .SI(\mem1[65][14] ), .SE(test_se), 
        .CLK(n1537), .Q(\mem1[65][15] ), .QN(n27121) );
  SDFFX1 \mem1_reg[65][14]  ( .D(n15034), .SI(\mem1[65][13] ), .SE(test_se), 
        .CLK(n1537), .Q(\mem1[65][14] ), .QN(n27122) );
  SDFFX1 \mem1_reg[65][13]  ( .D(n15033), .SI(\mem1[65][12] ), .SE(test_se), 
        .CLK(n1537), .Q(\mem1[65][13] ), .QN(n27123) );
  SDFFX1 \mem1_reg[65][12]  ( .D(n15032), .SI(\mem1[65][11] ), .SE(test_se), 
        .CLK(n1537), .Q(\mem1[65][12] ), .QN(n27124) );
  SDFFX1 \mem1_reg[65][11]  ( .D(n15031), .SI(\mem1[65][10] ), .SE(test_se), 
        .CLK(n1537), .Q(\mem1[65][11] ), .QN(n27125) );
  SDFFX1 \mem1_reg[65][10]  ( .D(n15030), .SI(\mem1[65][9] ), .SE(test_se), 
        .CLK(n1537), .Q(\mem1[65][10] ), .QN(n27126) );
  SDFFX1 \mem1_reg[65][9]  ( .D(n15029), .SI(\mem1[65][8] ), .SE(test_se), 
        .CLK(n1537), .Q(\mem1[65][9] ), .QN(n27127) );
  SDFFX1 \mem1_reg[65][8]  ( .D(n15028), .SI(\mem1[64][15] ), .SE(test_se), 
        .CLK(n1537), .Q(\mem1[65][8] ), .QN(n27128) );
  SDFFX1 \mem1_reg[64][15]  ( .D(n15027), .SI(\mem1[64][14] ), .SE(test_se), 
        .CLK(n1537), .Q(\mem1[64][15] ), .QN(n27129) );
  SDFFX1 \mem1_reg[64][14]  ( .D(n15026), .SI(\mem1[64][13] ), .SE(test_se), 
        .CLK(n1537), .Q(\mem1[64][14] ), .QN(n27130) );
  SDFFX1 \mem1_reg[64][13]  ( .D(n15025), .SI(\mem1[64][12] ), .SE(test_se), 
        .CLK(n1538), .Q(\mem1[64][13] ), .QN(n27131) );
  SDFFX1 \mem1_reg[64][12]  ( .D(n15024), .SI(\mem1[64][11] ), .SE(test_se), 
        .CLK(n1538), .Q(\mem1[64][12] ), .QN(n27132) );
  SDFFX1 \mem1_reg[64][11]  ( .D(n15023), .SI(\mem1[64][10] ), .SE(test_se), 
        .CLK(n1538), .Q(\mem1[64][11] ), .QN(n27133) );
  SDFFX1 \mem1_reg[64][10]  ( .D(n15022), .SI(\mem1[64][9] ), .SE(test_se), 
        .CLK(n1538), .Q(\mem1[64][10] ), .QN(n27134) );
  SDFFX1 \mem1_reg[64][9]  ( .D(n15021), .SI(\mem1[64][8] ), .SE(test_se), 
        .CLK(n1538), .Q(\mem1[64][9] ), .QN(n27135) );
  SDFFX1 \mem1_reg[64][8]  ( .D(n15020), .SI(\mem1[63][15] ), .SE(test_se), 
        .CLK(n1538), .Q(\mem1[64][8] ), .QN(n27136) );
  SDFFX1 \mem1_reg[63][15]  ( .D(n15019), .SI(\mem1[63][14] ), .SE(test_se), 
        .CLK(n1538), .Q(\mem1[63][15] ), .QN(n27137) );
  SDFFX1 \mem1_reg[63][14]  ( .D(n15018), .SI(\mem1[63][13] ), .SE(test_se), 
        .CLK(n1538), .Q(\mem1[63][14] ), .QN(n27138) );
  SDFFX1 \mem1_reg[63][13]  ( .D(n15017), .SI(\mem1[63][12] ), .SE(test_se), 
        .CLK(n1538), .Q(\mem1[63][13] ), .QN(n27139) );
  SDFFX1 \mem1_reg[63][12]  ( .D(n15016), .SI(\mem1[63][11] ), .SE(test_se), 
        .CLK(n1538), .Q(\mem1[63][12] ), .QN(n27140) );
  SDFFX1 \mem1_reg[63][11]  ( .D(n15015), .SI(\mem1[63][10] ), .SE(test_se), 
        .CLK(n1538), .Q(\mem1[63][11] ), .QN(n27141) );
  SDFFX1 \mem1_reg[63][10]  ( .D(n15014), .SI(\mem1[63][9] ), .SE(test_se), 
        .CLK(n1538), .Q(\mem1[63][10] ), .QN(n27142) );
  SDFFX1 \mem1_reg[63][9]  ( .D(n15013), .SI(\mem1[63][8] ), .SE(test_se), 
        .CLK(n1539), .Q(\mem1[63][9] ), .QN(n27143) );
  SDFFX1 \mem1_reg[63][8]  ( .D(n15012), .SI(\mem1[62][15] ), .SE(test_se), 
        .CLK(n1539), .Q(\mem1[63][8] ), .QN(n27144) );
  SDFFX1 \mem1_reg[62][15]  ( .D(n15011), .SI(\mem1[62][14] ), .SE(test_se), 
        .CLK(n1539), .Q(\mem1[62][15] ), .QN(n27145) );
  SDFFX1 \mem1_reg[62][14]  ( .D(n15010), .SI(\mem1[62][13] ), .SE(test_se), 
        .CLK(n1539), .Q(\mem1[62][14] ), .QN(n27146) );
  SDFFX1 \mem1_reg[62][13]  ( .D(n15009), .SI(\mem1[62][12] ), .SE(test_se), 
        .CLK(n1539), .Q(\mem1[62][13] ), .QN(n27147) );
  SDFFX1 \mem1_reg[62][12]  ( .D(n15008), .SI(\mem1[62][11] ), .SE(test_se), 
        .CLK(n1539), .Q(\mem1[62][12] ), .QN(n27148) );
  SDFFX1 \mem1_reg[62][11]  ( .D(n15007), .SI(\mem1[62][10] ), .SE(test_se), 
        .CLK(n1539), .Q(\mem1[62][11] ), .QN(n27149) );
  SDFFX1 \mem1_reg[62][10]  ( .D(n15006), .SI(\mem1[62][9] ), .SE(test_se), 
        .CLK(n1539), .Q(\mem1[62][10] ), .QN(n27150) );
  SDFFX1 \mem1_reg[62][9]  ( .D(n15005), .SI(\mem1[62][8] ), .SE(test_se), 
        .CLK(n1539), .Q(\mem1[62][9] ), .QN(n27151) );
  SDFFX1 \mem1_reg[62][8]  ( .D(n15004), .SI(\mem1[61][15] ), .SE(test_se), 
        .CLK(n1539), .Q(\mem1[62][8] ), .QN(n27152) );
  SDFFX1 \mem1_reg[61][15]  ( .D(n15003), .SI(\mem1[61][14] ), .SE(test_se), 
        .CLK(n1539), .Q(\mem1[61][15] ), .QN(n27153) );
  SDFFX1 \mem1_reg[61][14]  ( .D(n15002), .SI(\mem1[61][13] ), .SE(test_se), 
        .CLK(n1539), .Q(\mem1[61][14] ), .QN(n27154) );
  SDFFX1 \mem1_reg[61][13]  ( .D(n15001), .SI(\mem1[61][12] ), .SE(test_se), 
        .CLK(n1540), .Q(\mem1[61][13] ), .QN(n27155) );
  SDFFX1 \mem1_reg[61][12]  ( .D(n15000), .SI(\mem1[61][11] ), .SE(test_se), 
        .CLK(n1540), .Q(\mem1[61][12] ), .QN(n27156) );
  SDFFX1 \mem1_reg[61][11]  ( .D(n14999), .SI(\mem1[61][10] ), .SE(test_se), 
        .CLK(n1540), .Q(\mem1[61][11] ), .QN(n27157) );
  SDFFX1 \mem1_reg[61][10]  ( .D(n14998), .SI(\mem1[61][9] ), .SE(test_se), 
        .CLK(n1540), .Q(\mem1[61][10] ), .QN(n27158) );
  SDFFX1 \mem1_reg[61][9]  ( .D(n14997), .SI(\mem1[61][8] ), .SE(test_se), 
        .CLK(n1540), .Q(\mem1[61][9] ), .QN(n27159) );
  SDFFX1 \mem1_reg[61][8]  ( .D(n14996), .SI(\mem1[60][15] ), .SE(test_se), 
        .CLK(n1540), .Q(\mem1[61][8] ), .QN(n27160) );
  SDFFX1 \mem1_reg[60][15]  ( .D(n14995), .SI(\mem1[60][14] ), .SE(test_se), 
        .CLK(n1540), .Q(\mem1[60][15] ), .QN(n27161) );
  SDFFX1 \mem1_reg[60][14]  ( .D(n14994), .SI(\mem1[60][13] ), .SE(test_se), 
        .CLK(n1540), .Q(\mem1[60][14] ), .QN(n27162) );
  SDFFX1 \mem1_reg[60][13]  ( .D(n14993), .SI(\mem1[60][12] ), .SE(test_se), 
        .CLK(n1540), .Q(\mem1[60][13] ), .QN(n27163) );
  SDFFX1 \mem1_reg[60][12]  ( .D(n14992), .SI(\mem1[60][11] ), .SE(test_se), 
        .CLK(n1540), .Q(\mem1[60][12] ), .QN(n27164) );
  SDFFX1 \mem1_reg[60][11]  ( .D(n14991), .SI(\mem1[60][10] ), .SE(test_se), 
        .CLK(n1540), .Q(\mem1[60][11] ), .QN(n27165) );
  SDFFX1 \mem1_reg[60][10]  ( .D(n14990), .SI(\mem1[60][9] ), .SE(test_se), 
        .CLK(n1540), .Q(\mem1[60][10] ), .QN(n27166) );
  SDFFX1 \mem1_reg[60][9]  ( .D(n14989), .SI(\mem1[60][8] ), .SE(test_se), 
        .CLK(n1541), .Q(\mem1[60][9] ), .QN(n27167) );
  SDFFX1 \mem1_reg[60][8]  ( .D(n14988), .SI(\mem1[59][15] ), .SE(test_se), 
        .CLK(n1541), .Q(\mem1[60][8] ), .QN(n27168) );
  SDFFX1 \mem1_reg[59][15]  ( .D(n14987), .SI(\mem1[59][14] ), .SE(test_se), 
        .CLK(n1541), .Q(\mem1[59][15] ), .QN(n27169) );
  SDFFX1 \mem1_reg[59][14]  ( .D(n14986), .SI(\mem1[59][13] ), .SE(test_se), 
        .CLK(n1541), .Q(\mem1[59][14] ), .QN(n27170) );
  SDFFX1 \mem1_reg[59][13]  ( .D(n14985), .SI(\mem1[59][12] ), .SE(test_se), 
        .CLK(n1541), .Q(\mem1[59][13] ), .QN(n27171) );
  SDFFX1 \mem1_reg[59][12]  ( .D(n14984), .SI(\mem1[59][11] ), .SE(test_se), 
        .CLK(n1541), .Q(\mem1[59][12] ), .QN(n27172) );
  SDFFX1 \mem1_reg[59][11]  ( .D(n14983), .SI(\mem1[59][10] ), .SE(test_se), 
        .CLK(n1541), .Q(\mem1[59][11] ), .QN(n27173) );
  SDFFX1 \mem1_reg[59][10]  ( .D(n14982), .SI(\mem1[59][9] ), .SE(test_se), 
        .CLK(n1541), .Q(\mem1[59][10] ), .QN(n27174) );
  SDFFX1 \mem1_reg[59][9]  ( .D(n14981), .SI(\mem1[59][8] ), .SE(test_se), 
        .CLK(n1541), .Q(\mem1[59][9] ), .QN(n27175) );
  SDFFX1 \mem1_reg[59][8]  ( .D(n14980), .SI(\mem1[58][15] ), .SE(test_se), 
        .CLK(n1541), .Q(\mem1[59][8] ), .QN(n27176) );
  SDFFX1 \mem1_reg[58][15]  ( .D(n14979), .SI(\mem1[58][14] ), .SE(test_se), 
        .CLK(n1541), .Q(\mem1[58][15] ), .QN(n27177) );
  SDFFX1 \mem1_reg[58][14]  ( .D(n14978), .SI(\mem1[58][13] ), .SE(test_se), 
        .CLK(n1541), .Q(\mem1[58][14] ), .QN(n27178) );
  SDFFX1 \mem1_reg[58][13]  ( .D(n14977), .SI(\mem1[58][12] ), .SE(test_se), 
        .CLK(n1542), .Q(\mem1[58][13] ), .QN(n27179) );
  SDFFX1 \mem1_reg[58][12]  ( .D(n14976), .SI(\mem1[58][11] ), .SE(test_se), 
        .CLK(n1542), .Q(\mem1[58][12] ), .QN(n27180) );
  SDFFX1 \mem1_reg[58][11]  ( .D(n14975), .SI(\mem1[58][10] ), .SE(test_se), 
        .CLK(n1542), .Q(\mem1[58][11] ), .QN(n27181) );
  SDFFX1 \mem1_reg[58][10]  ( .D(n14974), .SI(\mem1[58][9] ), .SE(test_se), 
        .CLK(n1542), .Q(\mem1[58][10] ), .QN(n27182) );
  SDFFX1 \mem1_reg[58][9]  ( .D(n14973), .SI(\mem1[58][8] ), .SE(test_se), 
        .CLK(n1542), .Q(\mem1[58][9] ), .QN(n27183) );
  SDFFX1 \mem1_reg[58][8]  ( .D(n14972), .SI(\mem1[57][15] ), .SE(test_se), 
        .CLK(n1542), .Q(\mem1[58][8] ), .QN(n27184) );
  SDFFX1 \mem1_reg[57][15]  ( .D(n14971), .SI(\mem1[57][14] ), .SE(test_se), 
        .CLK(n1542), .Q(\mem1[57][15] ), .QN(n27185) );
  SDFFX1 \mem1_reg[57][14]  ( .D(n14970), .SI(\mem1[57][13] ), .SE(test_se), 
        .CLK(n1542), .Q(\mem1[57][14] ), .QN(n27186) );
  SDFFX1 \mem1_reg[57][13]  ( .D(n14969), .SI(\mem1[57][12] ), .SE(test_se), 
        .CLK(n1542), .Q(\mem1[57][13] ), .QN(n27187) );
  SDFFX1 \mem1_reg[57][12]  ( .D(n14968), .SI(\mem1[57][11] ), .SE(test_se), 
        .CLK(n1542), .Q(\mem1[57][12] ), .QN(n27188) );
  SDFFX1 \mem1_reg[57][11]  ( .D(n14967), .SI(\mem1[57][10] ), .SE(test_se), 
        .CLK(n1542), .Q(\mem1[57][11] ), .QN(n27189) );
  SDFFX1 \mem1_reg[57][10]  ( .D(n14966), .SI(\mem1[57][9] ), .SE(test_se), 
        .CLK(n1542), .Q(\mem1[57][10] ), .QN(n27190) );
  SDFFX1 \mem1_reg[57][9]  ( .D(n14965), .SI(\mem1[57][8] ), .SE(test_se), 
        .CLK(n1543), .Q(\mem1[57][9] ), .QN(n27191) );
  SDFFX1 \mem1_reg[57][8]  ( .D(n14964), .SI(\mem1[56][15] ), .SE(test_se), 
        .CLK(n1543), .Q(\mem1[57][8] ), .QN(n27192) );
  SDFFX1 \mem1_reg[56][15]  ( .D(n14963), .SI(\mem1[56][14] ), .SE(test_se), 
        .CLK(n1543), .Q(\mem1[56][15] ), .QN(n27193) );
  SDFFX1 \mem1_reg[56][14]  ( .D(n14962), .SI(\mem1[56][13] ), .SE(test_se), 
        .CLK(n1543), .Q(\mem1[56][14] ), .QN(n27194) );
  SDFFX1 \mem1_reg[56][13]  ( .D(n14961), .SI(\mem1[56][12] ), .SE(test_se), 
        .CLK(n1543), .Q(\mem1[56][13] ), .QN(n27195) );
  SDFFX1 \mem1_reg[56][12]  ( .D(n14960), .SI(\mem1[56][11] ), .SE(test_se), 
        .CLK(n1543), .Q(\mem1[56][12] ), .QN(n27196) );
  SDFFX1 \mem1_reg[56][11]  ( .D(n14959), .SI(\mem1[56][10] ), .SE(test_se), 
        .CLK(n1543), .Q(\mem1[56][11] ), .QN(n27197) );
  SDFFX1 \mem1_reg[56][10]  ( .D(n14958), .SI(\mem1[56][9] ), .SE(test_se), 
        .CLK(n1543), .Q(\mem1[56][10] ), .QN(n27198) );
  SDFFX1 \mem1_reg[56][9]  ( .D(n14957), .SI(\mem1[56][8] ), .SE(test_se), 
        .CLK(n1543), .Q(\mem1[56][9] ), .QN(n27199) );
  SDFFX1 \mem1_reg[56][8]  ( .D(n14956), .SI(\mem1[55][15] ), .SE(test_se), 
        .CLK(n1543), .Q(\mem1[56][8] ), .QN(n27200) );
  SDFFX1 \mem1_reg[55][15]  ( .D(n14955), .SI(\mem1[55][14] ), .SE(test_se), 
        .CLK(n1543), .Q(\mem1[55][15] ), .QN(n27201) );
  SDFFX1 \mem1_reg[55][14]  ( .D(n14954), .SI(\mem1[55][13] ), .SE(test_se), 
        .CLK(n1543), .Q(\mem1[55][14] ), .QN(n27202) );
  SDFFX1 \mem1_reg[55][13]  ( .D(n14953), .SI(\mem1[55][12] ), .SE(test_se), 
        .CLK(n1544), .Q(\mem1[55][13] ), .QN(n27203) );
  SDFFX1 \mem1_reg[55][12]  ( .D(n14952), .SI(\mem1[55][11] ), .SE(test_se), 
        .CLK(n1544), .Q(\mem1[55][12] ), .QN(n27204) );
  SDFFX1 \mem1_reg[55][11]  ( .D(n14951), .SI(\mem1[55][10] ), .SE(test_se), 
        .CLK(n1544), .Q(\mem1[55][11] ), .QN(n27205) );
  SDFFX1 \mem1_reg[55][10]  ( .D(n14950), .SI(\mem1[55][9] ), .SE(test_se), 
        .CLK(n1544), .Q(\mem1[55][10] ), .QN(n27206) );
  SDFFX1 \mem1_reg[55][9]  ( .D(n14949), .SI(\mem1[55][8] ), .SE(test_se), 
        .CLK(n1544), .Q(\mem1[55][9] ), .QN(n27207) );
  SDFFX1 \mem1_reg[55][8]  ( .D(n14948), .SI(\mem1[54][15] ), .SE(test_se), 
        .CLK(n1544), .Q(\mem1[55][8] ), .QN(n27208) );
  SDFFX1 \mem1_reg[54][15]  ( .D(n14947), .SI(\mem1[54][14] ), .SE(test_se), 
        .CLK(n1544), .Q(\mem1[54][15] ), .QN(n27209) );
  SDFFX1 \mem1_reg[54][14]  ( .D(n14946), .SI(\mem1[54][13] ), .SE(test_se), 
        .CLK(n1544), .Q(\mem1[54][14] ), .QN(n27210) );
  SDFFX1 \mem1_reg[54][13]  ( .D(n14945), .SI(\mem1[54][12] ), .SE(test_se), 
        .CLK(n1544), .Q(\mem1[54][13] ), .QN(n27211) );
  SDFFX1 \mem1_reg[54][12]  ( .D(n14944), .SI(\mem1[54][11] ), .SE(test_se), 
        .CLK(n1544), .Q(\mem1[54][12] ), .QN(n27212) );
  SDFFX1 \mem1_reg[54][11]  ( .D(n14943), .SI(\mem1[54][10] ), .SE(test_se), 
        .CLK(n1544), .Q(\mem1[54][11] ), .QN(n27213) );
  SDFFX1 \mem1_reg[54][10]  ( .D(n14942), .SI(\mem1[54][9] ), .SE(test_se), 
        .CLK(n1544), .Q(\mem1[54][10] ), .QN(n27214) );
  SDFFX1 \mem1_reg[54][9]  ( .D(n14941), .SI(\mem1[54][8] ), .SE(test_se), 
        .CLK(n1545), .Q(\mem1[54][9] ), .QN(n27215) );
  SDFFX1 \mem1_reg[54][8]  ( .D(n14940), .SI(\mem1[53][15] ), .SE(test_se), 
        .CLK(n1545), .Q(\mem1[54][8] ), .QN(n27216) );
  SDFFX1 \mem1_reg[53][15]  ( .D(n14939), .SI(\mem1[53][14] ), .SE(test_se), 
        .CLK(n1545), .Q(\mem1[53][15] ), .QN(n27217) );
  SDFFX1 \mem1_reg[53][14]  ( .D(n14938), .SI(\mem1[53][13] ), .SE(test_se), 
        .CLK(n1545), .Q(\mem1[53][14] ), .QN(n27218) );
  SDFFX1 \mem1_reg[53][13]  ( .D(n14937), .SI(\mem1[53][12] ), .SE(test_se), 
        .CLK(n1545), .Q(\mem1[53][13] ), .QN(n27219) );
  SDFFX1 \mem1_reg[53][12]  ( .D(n14936), .SI(\mem1[53][11] ), .SE(test_se), 
        .CLK(n1545), .Q(\mem1[53][12] ), .QN(n27220) );
  SDFFX1 \mem1_reg[53][11]  ( .D(n14935), .SI(\mem1[53][10] ), .SE(test_se), 
        .CLK(n1545), .Q(\mem1[53][11] ), .QN(n27221) );
  SDFFX1 \mem1_reg[53][10]  ( .D(n14934), .SI(\mem1[53][9] ), .SE(test_se), 
        .CLK(n1545), .Q(\mem1[53][10] ), .QN(n27222) );
  SDFFX1 \mem1_reg[53][9]  ( .D(n14933), .SI(\mem1[53][8] ), .SE(test_se), 
        .CLK(n1545), .Q(\mem1[53][9] ), .QN(n27223) );
  SDFFX1 \mem1_reg[53][8]  ( .D(n14932), .SI(\mem1[52][15] ), .SE(test_se), 
        .CLK(n1545), .Q(\mem1[53][8] ), .QN(n27224) );
  SDFFX1 \mem1_reg[52][15]  ( .D(n14931), .SI(\mem1[52][14] ), .SE(test_se), 
        .CLK(n1545), .Q(\mem1[52][15] ), .QN(n27225) );
  SDFFX1 \mem1_reg[52][14]  ( .D(n14930), .SI(\mem1[52][13] ), .SE(test_se), 
        .CLK(n1545), .Q(\mem1[52][14] ), .QN(n27226) );
  SDFFX1 \mem1_reg[52][13]  ( .D(n14929), .SI(\mem1[52][12] ), .SE(test_se), 
        .CLK(n1546), .Q(\mem1[52][13] ), .QN(n27227) );
  SDFFX1 \mem1_reg[52][12]  ( .D(n14928), .SI(\mem1[52][11] ), .SE(test_se), 
        .CLK(n1546), .Q(\mem1[52][12] ), .QN(n27228) );
  SDFFX1 \mem1_reg[52][11]  ( .D(n14927), .SI(\mem1[52][10] ), .SE(test_se), 
        .CLK(n1546), .Q(\mem1[52][11] ), .QN(n27229) );
  SDFFX1 \mem1_reg[52][10]  ( .D(n14926), .SI(\mem1[52][9] ), .SE(test_se), 
        .CLK(n1546), .Q(\mem1[52][10] ), .QN(n27230) );
  SDFFX1 \mem1_reg[52][9]  ( .D(n14925), .SI(\mem1[52][8] ), .SE(test_se), 
        .CLK(n1546), .Q(\mem1[52][9] ), .QN(n27231) );
  SDFFX1 \mem1_reg[52][8]  ( .D(n14924), .SI(\mem1[51][15] ), .SE(test_se), 
        .CLK(n1546), .Q(\mem1[52][8] ), .QN(n27232) );
  SDFFX1 \mem1_reg[51][15]  ( .D(n14923), .SI(\mem1[51][14] ), .SE(test_se), 
        .CLK(n1546), .Q(\mem1[51][15] ), .QN(n27233) );
  SDFFX1 \mem1_reg[51][14]  ( .D(n14922), .SI(\mem1[51][13] ), .SE(test_se), 
        .CLK(n1546), .Q(\mem1[51][14] ), .QN(n27234) );
  SDFFX1 \mem1_reg[51][13]  ( .D(n14921), .SI(\mem1[51][12] ), .SE(test_se), 
        .CLK(n1546), .Q(\mem1[51][13] ), .QN(n27235) );
  SDFFX1 \mem1_reg[51][12]  ( .D(n14920), .SI(\mem1[51][11] ), .SE(test_se), 
        .CLK(n1546), .Q(\mem1[51][12] ), .QN(n27236) );
  SDFFX1 \mem1_reg[51][11]  ( .D(n14919), .SI(\mem1[51][10] ), .SE(test_se), 
        .CLK(n1546), .Q(\mem1[51][11] ), .QN(n27237) );
  SDFFX1 \mem1_reg[51][10]  ( .D(n14918), .SI(\mem1[51][9] ), .SE(test_se), 
        .CLK(n1546), .Q(\mem1[51][10] ), .QN(n27238) );
  SDFFX1 \mem1_reg[51][9]  ( .D(n14917), .SI(\mem1[51][8] ), .SE(test_se), 
        .CLK(n1547), .Q(\mem1[51][9] ), .QN(n27239) );
  SDFFX1 \mem1_reg[51][8]  ( .D(n14916), .SI(\mem1[50][15] ), .SE(test_se), 
        .CLK(n1547), .Q(\mem1[51][8] ), .QN(n27240) );
  SDFFX1 \mem1_reg[50][15]  ( .D(n14915), .SI(\mem1[50][14] ), .SE(test_se), 
        .CLK(n1547), .Q(\mem1[50][15] ), .QN(n27241) );
  SDFFX1 \mem1_reg[50][14]  ( .D(n14914), .SI(\mem1[50][13] ), .SE(test_se), 
        .CLK(n1547), .Q(\mem1[50][14] ), .QN(n27242) );
  SDFFX1 \mem1_reg[50][13]  ( .D(n14913), .SI(\mem1[50][12] ), .SE(test_se), 
        .CLK(n1547), .Q(\mem1[50][13] ), .QN(n27243) );
  SDFFX1 \mem1_reg[50][12]  ( .D(n14912), .SI(\mem1[50][11] ), .SE(test_se), 
        .CLK(n1547), .Q(\mem1[50][12] ), .QN(n27244) );
  SDFFX1 \mem1_reg[50][11]  ( .D(n14911), .SI(\mem1[50][10] ), .SE(test_se), 
        .CLK(n1547), .Q(\mem1[50][11] ), .QN(n27245) );
  SDFFX1 \mem1_reg[50][10]  ( .D(n14910), .SI(\mem1[50][9] ), .SE(test_se), 
        .CLK(n1547), .Q(\mem1[50][10] ), .QN(n27246) );
  SDFFX1 \mem1_reg[50][9]  ( .D(n14909), .SI(\mem1[50][8] ), .SE(test_se), 
        .CLK(n1547), .Q(\mem1[50][9] ), .QN(n27247) );
  SDFFX1 \mem1_reg[50][8]  ( .D(n14908), .SI(\mem1[49][15] ), .SE(test_se), 
        .CLK(n1547), .Q(\mem1[50][8] ), .QN(n27248) );
  SDFFX1 \mem1_reg[49][15]  ( .D(n14907), .SI(\mem1[49][14] ), .SE(test_se), 
        .CLK(n1547), .Q(\mem1[49][15] ), .QN(n27249) );
  SDFFX1 \mem1_reg[49][14]  ( .D(n14906), .SI(\mem1[49][13] ), .SE(test_se), 
        .CLK(n1547), .Q(\mem1[49][14] ), .QN(n27250) );
  SDFFX1 \mem1_reg[49][13]  ( .D(n14905), .SI(\mem1[49][12] ), .SE(test_se), 
        .CLK(n1548), .Q(\mem1[49][13] ), .QN(n27251) );
  SDFFX1 \mem1_reg[49][12]  ( .D(n14904), .SI(\mem1[49][11] ), .SE(test_se), 
        .CLK(n1548), .Q(\mem1[49][12] ), .QN(n27252) );
  SDFFX1 \mem1_reg[49][11]  ( .D(n14903), .SI(\mem1[49][10] ), .SE(test_se), 
        .CLK(n1548), .Q(\mem1[49][11] ), .QN(n27253) );
  SDFFX1 \mem1_reg[49][10]  ( .D(n14902), .SI(\mem1[49][9] ), .SE(test_se), 
        .CLK(n1548), .Q(\mem1[49][10] ), .QN(n27254) );
  SDFFX1 \mem1_reg[49][9]  ( .D(n14901), .SI(\mem1[49][8] ), .SE(test_se), 
        .CLK(n1548), .Q(\mem1[49][9] ), .QN(n27255) );
  SDFFX1 \mem1_reg[49][8]  ( .D(n14900), .SI(\mem1[48][15] ), .SE(test_se), 
        .CLK(n1548), .Q(\mem1[49][8] ), .QN(n27256) );
  SDFFX1 \mem1_reg[48][15]  ( .D(n14899), .SI(\mem1[48][14] ), .SE(test_se), 
        .CLK(n1548), .Q(\mem1[48][15] ), .QN(n27257) );
  SDFFX1 \mem1_reg[48][14]  ( .D(n14898), .SI(\mem1[48][13] ), .SE(test_se), 
        .CLK(n1548), .Q(\mem1[48][14] ), .QN(n27258) );
  SDFFX1 \mem1_reg[48][13]  ( .D(n14897), .SI(\mem1[48][12] ), .SE(test_se), 
        .CLK(n1548), .Q(\mem1[48][13] ), .QN(n27259) );
  SDFFX1 \mem1_reg[48][12]  ( .D(n14896), .SI(\mem1[48][11] ), .SE(test_se), 
        .CLK(n1548), .Q(\mem1[48][12] ), .QN(n27260) );
  SDFFX1 \mem1_reg[48][11]  ( .D(n14895), .SI(\mem1[48][10] ), .SE(test_se), 
        .CLK(n1548), .Q(\mem1[48][11] ), .QN(n27261) );
  SDFFX1 \mem1_reg[48][10]  ( .D(n14894), .SI(\mem1[48][9] ), .SE(test_se), 
        .CLK(n1548), .Q(\mem1[48][10] ), .QN(n27262) );
  SDFFX1 \mem1_reg[48][9]  ( .D(n14893), .SI(\mem1[48][8] ), .SE(test_se), 
        .CLK(n1549), .Q(\mem1[48][9] ), .QN(n27263) );
  SDFFX1 \mem1_reg[48][8]  ( .D(n14892), .SI(\mem1[47][15] ), .SE(test_se), 
        .CLK(n1549), .Q(\mem1[48][8] ), .QN(n27264) );
  SDFFX1 \mem1_reg[47][15]  ( .D(n14891), .SI(\mem1[47][14] ), .SE(test_se), 
        .CLK(n1549), .Q(\mem1[47][15] ), .QN(n27265) );
  SDFFX1 \mem1_reg[47][14]  ( .D(n14890), .SI(\mem1[47][13] ), .SE(test_se), 
        .CLK(n1549), .Q(\mem1[47][14] ), .QN(n27266) );
  SDFFX1 \mem1_reg[47][13]  ( .D(n14889), .SI(\mem1[47][12] ), .SE(test_se), 
        .CLK(n1549), .Q(\mem1[47][13] ), .QN(n27267) );
  SDFFX1 \mem1_reg[47][12]  ( .D(n14888), .SI(\mem1[47][11] ), .SE(test_se), 
        .CLK(n1549), .Q(\mem1[47][12] ), .QN(n27268) );
  SDFFX1 \mem1_reg[47][11]  ( .D(n14887), .SI(\mem1[47][10] ), .SE(test_se), 
        .CLK(n1549), .Q(\mem1[47][11] ), .QN(n27269) );
  SDFFX1 \mem1_reg[47][10]  ( .D(n14886), .SI(\mem1[47][9] ), .SE(test_se), 
        .CLK(n1549), .Q(\mem1[47][10] ), .QN(n27270) );
  SDFFX1 \mem1_reg[47][9]  ( .D(n14885), .SI(\mem1[47][8] ), .SE(test_se), 
        .CLK(n1549), .Q(\mem1[47][9] ), .QN(n27271) );
  SDFFX1 \mem1_reg[47][8]  ( .D(n14884), .SI(\mem1[46][15] ), .SE(test_se), 
        .CLK(n1549), .Q(\mem1[47][8] ), .QN(n27272) );
  SDFFX1 \mem1_reg[46][15]  ( .D(n14883), .SI(\mem1[46][14] ), .SE(test_se), 
        .CLK(n1549), .Q(\mem1[46][15] ), .QN(n27273) );
  SDFFX1 \mem1_reg[46][14]  ( .D(n14882), .SI(\mem1[46][13] ), .SE(test_se), 
        .CLK(n1549), .Q(\mem1[46][14] ), .QN(n27274) );
  SDFFX1 \mem1_reg[46][13]  ( .D(n14881), .SI(\mem1[46][12] ), .SE(test_se), 
        .CLK(n1550), .Q(\mem1[46][13] ), .QN(n27275) );
  SDFFX1 \mem1_reg[46][12]  ( .D(n14880), .SI(\mem1[46][11] ), .SE(test_se), 
        .CLK(n1550), .Q(\mem1[46][12] ), .QN(n27276) );
  SDFFX1 \mem1_reg[46][11]  ( .D(n14879), .SI(\mem1[46][10] ), .SE(test_se), 
        .CLK(n1550), .Q(\mem1[46][11] ), .QN(n27277) );
  SDFFX1 \mem1_reg[46][10]  ( .D(n14878), .SI(\mem1[46][9] ), .SE(test_se), 
        .CLK(n1550), .Q(\mem1[46][10] ), .QN(n27278) );
  SDFFX1 \mem1_reg[46][9]  ( .D(n14877), .SI(\mem1[46][8] ), .SE(test_se), 
        .CLK(n1550), .Q(\mem1[46][9] ), .QN(n27279) );
  SDFFX1 \mem1_reg[46][8]  ( .D(n14876), .SI(\mem1[45][15] ), .SE(test_se), 
        .CLK(n1550), .Q(\mem1[46][8] ), .QN(n27280) );
  SDFFX1 \mem1_reg[45][15]  ( .D(n14875), .SI(\mem1[45][14] ), .SE(test_se), 
        .CLK(n1550), .Q(\mem1[45][15] ), .QN(n27281) );
  SDFFX1 \mem1_reg[45][14]  ( .D(n14874), .SI(\mem1[45][13] ), .SE(test_se), 
        .CLK(n1550), .Q(\mem1[45][14] ), .QN(n27282) );
  SDFFX1 \mem1_reg[45][13]  ( .D(n14873), .SI(\mem1[45][12] ), .SE(test_se), 
        .CLK(n1550), .Q(\mem1[45][13] ), .QN(n27283) );
  SDFFX1 \mem1_reg[45][12]  ( .D(n14872), .SI(\mem1[45][11] ), .SE(test_se), 
        .CLK(n1550), .Q(\mem1[45][12] ), .QN(n27284) );
  SDFFX1 \mem1_reg[45][11]  ( .D(n14871), .SI(\mem1[45][10] ), .SE(test_se), 
        .CLK(n1550), .Q(\mem1[45][11] ), .QN(n27285) );
  SDFFX1 \mem1_reg[45][10]  ( .D(n14870), .SI(\mem1[45][9] ), .SE(test_se), 
        .CLK(n1550), .Q(\mem1[45][10] ), .QN(n27286) );
  SDFFX1 \mem1_reg[45][9]  ( .D(n14869), .SI(\mem1[45][8] ), .SE(test_se), 
        .CLK(n1551), .Q(\mem1[45][9] ), .QN(n27287) );
  SDFFX1 \mem1_reg[45][8]  ( .D(n14868), .SI(\mem1[44][15] ), .SE(test_se), 
        .CLK(n1551), .Q(\mem1[45][8] ), .QN(n27288) );
  SDFFX1 \mem1_reg[44][15]  ( .D(n14867), .SI(\mem1[44][14] ), .SE(test_se), 
        .CLK(n1551), .Q(\mem1[44][15] ), .QN(n27289) );
  SDFFX1 \mem1_reg[44][14]  ( .D(n14866), .SI(\mem1[44][13] ), .SE(test_se), 
        .CLK(n1551), .Q(\mem1[44][14] ), .QN(n27290) );
  SDFFX1 \mem1_reg[44][13]  ( .D(n14865), .SI(\mem1[44][12] ), .SE(test_se), 
        .CLK(n1551), .Q(\mem1[44][13] ), .QN(n27291) );
  SDFFX1 \mem1_reg[44][12]  ( .D(n14864), .SI(\mem1[44][11] ), .SE(test_se), 
        .CLK(n1551), .Q(\mem1[44][12] ), .QN(n27292) );
  SDFFX1 \mem1_reg[44][11]  ( .D(n14863), .SI(\mem1[44][10] ), .SE(test_se), 
        .CLK(n1551), .Q(\mem1[44][11] ), .QN(n27293) );
  SDFFX1 \mem1_reg[44][10]  ( .D(n14862), .SI(\mem1[44][9] ), .SE(test_se), 
        .CLK(n1551), .Q(\mem1[44][10] ), .QN(n27294) );
  SDFFX1 \mem1_reg[44][9]  ( .D(n14861), .SI(\mem1[44][8] ), .SE(test_se), 
        .CLK(n1551), .Q(\mem1[44][9] ), .QN(n27295) );
  SDFFX1 \mem1_reg[44][8]  ( .D(n14860), .SI(\mem1[43][15] ), .SE(test_se), 
        .CLK(n1551), .Q(\mem1[44][8] ), .QN(n27296) );
  SDFFX1 \mem1_reg[43][15]  ( .D(n14859), .SI(\mem1[43][14] ), .SE(test_se), 
        .CLK(n1551), .Q(\mem1[43][15] ), .QN(n27297) );
  SDFFX1 \mem1_reg[43][14]  ( .D(n14858), .SI(\mem1[43][13] ), .SE(test_se), 
        .CLK(n1551), .Q(\mem1[43][14] ), .QN(n27298) );
  SDFFX1 \mem1_reg[43][13]  ( .D(n14857), .SI(\mem1[43][12] ), .SE(test_se), 
        .CLK(n1552), .Q(\mem1[43][13] ), .QN(n27299) );
  SDFFX1 \mem1_reg[43][12]  ( .D(n14856), .SI(\mem1[43][11] ), .SE(test_se), 
        .CLK(n1552), .Q(\mem1[43][12] ), .QN(n27300) );
  SDFFX1 \mem1_reg[43][11]  ( .D(n14855), .SI(\mem1[43][10] ), .SE(test_se), 
        .CLK(n1552), .Q(\mem1[43][11] ), .QN(n27301) );
  SDFFX1 \mem1_reg[43][10]  ( .D(n14854), .SI(\mem1[43][9] ), .SE(test_se), 
        .CLK(n1552), .Q(\mem1[43][10] ), .QN(n27302) );
  SDFFX1 \mem1_reg[43][9]  ( .D(n14853), .SI(\mem1[43][8] ), .SE(test_se), 
        .CLK(n1552), .Q(\mem1[43][9] ), .QN(n27303) );
  SDFFX1 \mem1_reg[43][8]  ( .D(n14852), .SI(\mem1[42][15] ), .SE(test_se), 
        .CLK(n1552), .Q(\mem1[43][8] ), .QN(n27304) );
  SDFFX1 \mem1_reg[42][15]  ( .D(n14851), .SI(\mem1[42][14] ), .SE(test_se), 
        .CLK(n1552), .Q(\mem1[42][15] ), .QN(n27305) );
  SDFFX1 \mem1_reg[42][14]  ( .D(n14850), .SI(\mem1[42][13] ), .SE(test_se), 
        .CLK(n1552), .Q(\mem1[42][14] ), .QN(n27306) );
  SDFFX1 \mem1_reg[42][13]  ( .D(n14849), .SI(\mem1[42][12] ), .SE(test_se), 
        .CLK(n1552), .Q(\mem1[42][13] ), .QN(n27307) );
  SDFFX1 \mem1_reg[42][12]  ( .D(n14848), .SI(\mem1[42][11] ), .SE(test_se), 
        .CLK(n1552), .Q(\mem1[42][12] ), .QN(n27308) );
  SDFFX1 \mem1_reg[42][11]  ( .D(n14847), .SI(\mem1[42][10] ), .SE(test_se), 
        .CLK(n1552), .Q(\mem1[42][11] ), .QN(n27309) );
  SDFFX1 \mem1_reg[42][10]  ( .D(n14846), .SI(\mem1[42][9] ), .SE(test_se), 
        .CLK(n1552), .Q(\mem1[42][10] ), .QN(n27310) );
  SDFFX1 \mem1_reg[42][9]  ( .D(n14845), .SI(\mem1[42][8] ), .SE(test_se), 
        .CLK(n1553), .Q(\mem1[42][9] ), .QN(n27311) );
  SDFFX1 \mem1_reg[42][8]  ( .D(n14844), .SI(\mem1[41][15] ), .SE(test_se), 
        .CLK(n1553), .Q(\mem1[42][8] ), .QN(n27312) );
  SDFFX1 \mem1_reg[41][15]  ( .D(n14843), .SI(\mem1[41][14] ), .SE(test_se), 
        .CLK(n1553), .Q(\mem1[41][15] ), .QN(n27313) );
  SDFFX1 \mem1_reg[41][14]  ( .D(n14842), .SI(\mem1[41][13] ), .SE(test_se), 
        .CLK(n1553), .Q(\mem1[41][14] ), .QN(n27314) );
  SDFFX1 \mem1_reg[41][13]  ( .D(n14841), .SI(\mem1[41][12] ), .SE(test_se), 
        .CLK(n1553), .Q(\mem1[41][13] ), .QN(n27315) );
  SDFFX1 \mem1_reg[41][12]  ( .D(n14840), .SI(\mem1[41][11] ), .SE(test_se), 
        .CLK(n1553), .Q(\mem1[41][12] ), .QN(n27316) );
  SDFFX1 \mem1_reg[41][11]  ( .D(n14839), .SI(\mem1[41][10] ), .SE(test_se), 
        .CLK(n1553), .Q(\mem1[41][11] ), .QN(n27317) );
  SDFFX1 \mem1_reg[41][10]  ( .D(n14838), .SI(\mem1[41][9] ), .SE(test_se), 
        .CLK(n1553), .Q(\mem1[41][10] ), .QN(n27318) );
  SDFFX1 \mem1_reg[41][9]  ( .D(n14837), .SI(\mem1[41][8] ), .SE(test_se), 
        .CLK(n1553), .Q(\mem1[41][9] ), .QN(n27319) );
  SDFFX1 \mem1_reg[41][8]  ( .D(n14836), .SI(\mem1[40][15] ), .SE(test_se), 
        .CLK(n1553), .Q(\mem1[41][8] ), .QN(n27320) );
  SDFFX1 \mem1_reg[40][15]  ( .D(n14835), .SI(\mem1[40][14] ), .SE(test_se), 
        .CLK(n1553), .Q(\mem1[40][15] ), .QN(n27321) );
  SDFFX1 \mem1_reg[40][14]  ( .D(n14834), .SI(\mem1[40][13] ), .SE(test_se), 
        .CLK(n1553), .Q(\mem1[40][14] ), .QN(n27322) );
  SDFFX1 \mem1_reg[40][13]  ( .D(n14833), .SI(\mem1[40][12] ), .SE(test_se), 
        .CLK(n1554), .Q(\mem1[40][13] ), .QN(n27323) );
  SDFFX1 \mem1_reg[40][12]  ( .D(n14832), .SI(\mem1[40][11] ), .SE(test_se), 
        .CLK(n1554), .Q(\mem1[40][12] ), .QN(n27324) );
  SDFFX1 \mem1_reg[40][11]  ( .D(n14831), .SI(\mem1[40][10] ), .SE(test_se), 
        .CLK(n1554), .Q(\mem1[40][11] ), .QN(n27325) );
  SDFFX1 \mem1_reg[40][10]  ( .D(n14830), .SI(\mem1[40][9] ), .SE(test_se), 
        .CLK(n1554), .Q(\mem1[40][10] ), .QN(n27326) );
  SDFFX1 \mem1_reg[40][9]  ( .D(n14829), .SI(\mem1[40][8] ), .SE(test_se), 
        .CLK(n1554), .Q(\mem1[40][9] ), .QN(n27327) );
  SDFFX1 \mem1_reg[40][8]  ( .D(n14828), .SI(\mem1[39][15] ), .SE(test_se), 
        .CLK(n1554), .Q(\mem1[40][8] ), .QN(n27328) );
  SDFFX1 \mem1_reg[39][15]  ( .D(n14827), .SI(\mem1[39][14] ), .SE(test_se), 
        .CLK(n1554), .Q(\mem1[39][15] ), .QN(n27329) );
  SDFFX1 \mem1_reg[39][14]  ( .D(n14826), .SI(\mem1[39][13] ), .SE(test_se), 
        .CLK(n1554), .Q(\mem1[39][14] ), .QN(n27330) );
  SDFFX1 \mem1_reg[39][13]  ( .D(n14825), .SI(\mem1[39][12] ), .SE(test_se), 
        .CLK(n1554), .Q(\mem1[39][13] ), .QN(n27331) );
  SDFFX1 \mem1_reg[39][12]  ( .D(n14824), .SI(\mem1[39][11] ), .SE(test_se), 
        .CLK(n1554), .Q(\mem1[39][12] ), .QN(n27332) );
  SDFFX1 \mem1_reg[39][11]  ( .D(n14823), .SI(\mem1[39][10] ), .SE(test_se), 
        .CLK(n1554), .Q(\mem1[39][11] ), .QN(n27333) );
  SDFFX1 \mem1_reg[39][10]  ( .D(n14822), .SI(\mem1[39][9] ), .SE(test_se), 
        .CLK(n1554), .Q(\mem1[39][10] ), .QN(n27334) );
  SDFFX1 \mem1_reg[39][9]  ( .D(n14821), .SI(\mem1[39][8] ), .SE(test_se), 
        .CLK(n1555), .Q(\mem1[39][9] ), .QN(n27335) );
  SDFFX1 \mem1_reg[39][8]  ( .D(n14820), .SI(\mem1[38][15] ), .SE(test_se), 
        .CLK(n1555), .Q(\mem1[39][8] ), .QN(n27336) );
  SDFFX1 \mem1_reg[38][15]  ( .D(n14819), .SI(\mem1[38][14] ), .SE(test_se), 
        .CLK(n1555), .Q(\mem1[38][15] ), .QN(n27337) );
  SDFFX1 \mem1_reg[38][14]  ( .D(n14818), .SI(\mem1[38][13] ), .SE(test_se), 
        .CLK(n1555), .Q(\mem1[38][14] ), .QN(n27338) );
  SDFFX1 \mem1_reg[38][13]  ( .D(n14817), .SI(\mem1[38][12] ), .SE(test_se), 
        .CLK(n1555), .Q(\mem1[38][13] ), .QN(n27339) );
  SDFFX1 \mem1_reg[38][12]  ( .D(n14816), .SI(\mem1[38][11] ), .SE(test_se), 
        .CLK(n1555), .Q(\mem1[38][12] ), .QN(n27340) );
  SDFFX1 \mem1_reg[38][11]  ( .D(n14815), .SI(\mem1[38][10] ), .SE(test_se), 
        .CLK(n1555), .Q(\mem1[38][11] ), .QN(n27341) );
  SDFFX1 \mem1_reg[38][10]  ( .D(n14814), .SI(\mem1[38][9] ), .SE(test_se), 
        .CLK(n1555), .Q(\mem1[38][10] ), .QN(n27342) );
  SDFFX1 \mem1_reg[38][9]  ( .D(n14813), .SI(\mem1[38][8] ), .SE(test_se), 
        .CLK(n1555), .Q(\mem1[38][9] ), .QN(n27343) );
  SDFFX1 \mem1_reg[38][8]  ( .D(n14812), .SI(\mem1[37][15] ), .SE(test_se), 
        .CLK(n1555), .Q(\mem1[38][8] ), .QN(n27344) );
  SDFFX1 \mem1_reg[37][15]  ( .D(n14811), .SI(\mem1[37][14] ), .SE(test_se), 
        .CLK(n1555), .Q(\mem1[37][15] ), .QN(n27345) );
  SDFFX1 \mem1_reg[37][14]  ( .D(n14810), .SI(\mem1[37][13] ), .SE(test_se), 
        .CLK(n1555), .Q(\mem1[37][14] ), .QN(n27346) );
  SDFFX1 \mem1_reg[37][13]  ( .D(n14809), .SI(\mem1[37][12] ), .SE(test_se), 
        .CLK(n1556), .Q(\mem1[37][13] ), .QN(n27347) );
  SDFFX1 \mem1_reg[37][12]  ( .D(n14808), .SI(\mem1[37][11] ), .SE(test_se), 
        .CLK(n1556), .Q(\mem1[37][12] ), .QN(n27348) );
  SDFFX1 \mem1_reg[37][11]  ( .D(n14807), .SI(\mem1[37][10] ), .SE(test_se), 
        .CLK(n1556), .Q(\mem1[37][11] ), .QN(n27349) );
  SDFFX1 \mem1_reg[37][10]  ( .D(n14806), .SI(\mem1[37][9] ), .SE(test_se), 
        .CLK(n1556), .Q(\mem1[37][10] ), .QN(n27350) );
  SDFFX1 \mem1_reg[37][9]  ( .D(n14805), .SI(\mem1[37][8] ), .SE(test_se), 
        .CLK(n1556), .Q(\mem1[37][9] ), .QN(n27351) );
  SDFFX1 \mem1_reg[37][8]  ( .D(n14804), .SI(\mem1[36][15] ), .SE(test_se), 
        .CLK(n1556), .Q(\mem1[37][8] ), .QN(n27352) );
  SDFFX1 \mem1_reg[36][15]  ( .D(n14803), .SI(\mem1[36][14] ), .SE(test_se), 
        .CLK(n1556), .Q(\mem1[36][15] ), .QN(n27353) );
  SDFFX1 \mem1_reg[36][14]  ( .D(n14802), .SI(\mem1[36][13] ), .SE(test_se), 
        .CLK(n1556), .Q(\mem1[36][14] ), .QN(n27354) );
  SDFFX1 \mem1_reg[36][13]  ( .D(n14801), .SI(\mem1[36][12] ), .SE(test_se), 
        .CLK(n1556), .Q(\mem1[36][13] ), .QN(n27355) );
  SDFFX1 \mem1_reg[36][12]  ( .D(n14800), .SI(\mem1[36][11] ), .SE(test_se), 
        .CLK(n1556), .Q(\mem1[36][12] ), .QN(n27356) );
  SDFFX1 \mem1_reg[36][11]  ( .D(n14799), .SI(\mem1[36][10] ), .SE(test_se), 
        .CLK(n1556), .Q(\mem1[36][11] ), .QN(n27357) );
  SDFFX1 \mem1_reg[36][10]  ( .D(n14798), .SI(\mem1[36][9] ), .SE(test_se), 
        .CLK(n1556), .Q(\mem1[36][10] ), .QN(n27358) );
  SDFFX1 \mem1_reg[36][9]  ( .D(n14797), .SI(\mem1[36][8] ), .SE(test_se), 
        .CLK(n1557), .Q(\mem1[36][9] ), .QN(n27359) );
  SDFFX1 \mem1_reg[36][8]  ( .D(n14796), .SI(\mem1[35][15] ), .SE(test_se), 
        .CLK(n1557), .Q(\mem1[36][8] ), .QN(n27360) );
  SDFFX1 \mem1_reg[35][15]  ( .D(n14795), .SI(\mem1[35][14] ), .SE(test_se), 
        .CLK(n1557), .Q(\mem1[35][15] ), .QN(n27361) );
  SDFFX1 \mem1_reg[35][14]  ( .D(n14794), .SI(\mem1[35][13] ), .SE(test_se), 
        .CLK(n1557), .Q(\mem1[35][14] ), .QN(n27362) );
  SDFFX1 \mem1_reg[35][13]  ( .D(n14793), .SI(\mem1[35][12] ), .SE(test_se), 
        .CLK(n1557), .Q(\mem1[35][13] ), .QN(n27363) );
  SDFFX1 \mem1_reg[35][12]  ( .D(n14792), .SI(\mem1[35][11] ), .SE(test_se), 
        .CLK(n1557), .Q(\mem1[35][12] ), .QN(n27364) );
  SDFFX1 \mem1_reg[35][11]  ( .D(n14791), .SI(\mem1[35][10] ), .SE(test_se), 
        .CLK(n1557), .Q(\mem1[35][11] ), .QN(n27365) );
  SDFFX1 \mem1_reg[35][10]  ( .D(n14790), .SI(\mem1[35][9] ), .SE(test_se), 
        .CLK(n1557), .Q(\mem1[35][10] ), .QN(n27366) );
  SDFFX1 \mem1_reg[35][9]  ( .D(n14789), .SI(\mem1[35][8] ), .SE(test_se), 
        .CLK(n1557), .Q(\mem1[35][9] ), .QN(n27367) );
  SDFFX1 \mem1_reg[35][8]  ( .D(n14788), .SI(\mem1[34][15] ), .SE(test_se), 
        .CLK(n1557), .Q(\mem1[35][8] ), .QN(n27368) );
  SDFFX1 \mem1_reg[34][15]  ( .D(n14787), .SI(\mem1[34][14] ), .SE(test_se), 
        .CLK(n1557), .Q(\mem1[34][15] ), .QN(n27369) );
  SDFFX1 \mem1_reg[34][14]  ( .D(n14786), .SI(\mem1[34][13] ), .SE(test_se), 
        .CLK(n1557), .Q(\mem1[34][14] ), .QN(n27370) );
  SDFFX1 \mem1_reg[34][13]  ( .D(n14785), .SI(\mem1[34][12] ), .SE(test_se), 
        .CLK(n1558), .Q(\mem1[34][13] ), .QN(n27371) );
  SDFFX1 \mem1_reg[34][12]  ( .D(n14784), .SI(\mem1[34][11] ), .SE(test_se), 
        .CLK(n1558), .Q(\mem1[34][12] ), .QN(n27372) );
  SDFFX1 \mem1_reg[34][11]  ( .D(n14783), .SI(\mem1[34][10] ), .SE(test_se), 
        .CLK(n1558), .Q(\mem1[34][11] ), .QN(n27373) );
  SDFFX1 \mem1_reg[34][10]  ( .D(n14782), .SI(\mem1[34][9] ), .SE(test_se), 
        .CLK(n1558), .Q(\mem1[34][10] ), .QN(n27374) );
  SDFFX1 \mem1_reg[34][9]  ( .D(n14781), .SI(\mem1[34][8] ), .SE(test_se), 
        .CLK(n1558), .Q(\mem1[34][9] ), .QN(n27375) );
  SDFFX1 \mem1_reg[34][8]  ( .D(n14780), .SI(\mem1[33][15] ), .SE(test_se), 
        .CLK(n1558), .Q(\mem1[34][8] ), .QN(n27376) );
  SDFFX1 \mem1_reg[33][15]  ( .D(n14779), .SI(\mem1[33][14] ), .SE(test_se), 
        .CLK(n1558), .Q(\mem1[33][15] ), .QN(n27377) );
  SDFFX1 \mem1_reg[33][14]  ( .D(n14778), .SI(\mem1[33][13] ), .SE(test_se), 
        .CLK(n1558), .Q(\mem1[33][14] ), .QN(n27378) );
  SDFFX1 \mem1_reg[33][13]  ( .D(n14777), .SI(\mem1[33][12] ), .SE(test_se), 
        .CLK(n1558), .Q(\mem1[33][13] ), .QN(n27379) );
  SDFFX1 \mem1_reg[33][12]  ( .D(n14776), .SI(\mem1[33][11] ), .SE(test_se), 
        .CLK(n1558), .Q(\mem1[33][12] ), .QN(n27380) );
  SDFFX1 \mem1_reg[33][11]  ( .D(n14775), .SI(\mem1[33][10] ), .SE(test_se), 
        .CLK(n1558), .Q(\mem1[33][11] ), .QN(n27381) );
  SDFFX1 \mem1_reg[33][10]  ( .D(n14774), .SI(\mem1[33][9] ), .SE(test_se), 
        .CLK(n1558), .Q(\mem1[33][10] ), .QN(n27382) );
  SDFFX1 \mem1_reg[33][9]  ( .D(n14773), .SI(\mem1[33][8] ), .SE(test_se), 
        .CLK(n1559), .Q(\mem1[33][9] ), .QN(n27383) );
  SDFFX1 \mem1_reg[33][8]  ( .D(n14772), .SI(\mem1[32][15] ), .SE(test_se), 
        .CLK(n1559), .Q(\mem1[33][8] ), .QN(n27384) );
  SDFFX1 \mem1_reg[32][15]  ( .D(n14771), .SI(\mem1[32][14] ), .SE(test_se), 
        .CLK(n1559), .Q(\mem1[32][15] ), .QN(n27385) );
  SDFFX1 \mem1_reg[32][14]  ( .D(n14770), .SI(\mem1[32][13] ), .SE(test_se), 
        .CLK(n1559), .Q(\mem1[32][14] ), .QN(n27386) );
  SDFFX1 \mem1_reg[32][13]  ( .D(n14769), .SI(\mem1[32][12] ), .SE(test_se), 
        .CLK(n1559), .Q(\mem1[32][13] ), .QN(n27387) );
  SDFFX1 \mem1_reg[32][12]  ( .D(n14768), .SI(\mem1[32][11] ), .SE(test_se), 
        .CLK(n1559), .Q(\mem1[32][12] ), .QN(n27388) );
  SDFFX1 \mem1_reg[32][11]  ( .D(n14767), .SI(\mem1[32][10] ), .SE(test_se), 
        .CLK(n1559), .Q(\mem1[32][11] ), .QN(n27389) );
  SDFFX1 \mem1_reg[32][10]  ( .D(n14766), .SI(\mem1[32][9] ), .SE(test_se), 
        .CLK(n1559), .Q(\mem1[32][10] ), .QN(n27390) );
  SDFFX1 \mem1_reg[32][9]  ( .D(n14765), .SI(\mem1[32][8] ), .SE(test_se), 
        .CLK(n1559), .Q(\mem1[32][9] ), .QN(n27391) );
  SDFFX1 \mem1_reg[32][8]  ( .D(n14764), .SI(\mem1[31][15] ), .SE(test_se), 
        .CLK(n1559), .Q(\mem1[32][8] ), .QN(n27392) );
  SDFFX1 \mem1_reg[31][15]  ( .D(n14763), .SI(\mem1[31][14] ), .SE(test_se), 
        .CLK(n1559), .Q(\mem1[31][15] ), .QN(n27393) );
  SDFFX1 \mem1_reg[31][14]  ( .D(n14762), .SI(\mem1[31][13] ), .SE(test_se), 
        .CLK(n1559), .Q(\mem1[31][14] ), .QN(n27394) );
  SDFFX1 \mem1_reg[31][13]  ( .D(n14761), .SI(\mem1[31][12] ), .SE(test_se), 
        .CLK(n1560), .Q(\mem1[31][13] ), .QN(n27395) );
  SDFFX1 \mem1_reg[31][12]  ( .D(n14760), .SI(\mem1[31][11] ), .SE(test_se), 
        .CLK(n1560), .Q(\mem1[31][12] ), .QN(n27396) );
  SDFFX1 \mem1_reg[31][11]  ( .D(n14759), .SI(\mem1[31][10] ), .SE(test_se), 
        .CLK(n1560), .Q(\mem1[31][11] ), .QN(n27397) );
  SDFFX1 \mem1_reg[31][10]  ( .D(n14758), .SI(\mem1[31][9] ), .SE(test_se), 
        .CLK(n1560), .Q(\mem1[31][10] ), .QN(n27398) );
  SDFFX1 \mem1_reg[31][9]  ( .D(n14757), .SI(\mem1[31][8] ), .SE(test_se), 
        .CLK(n1560), .Q(\mem1[31][9] ), .QN(n27399) );
  SDFFX1 \mem1_reg[31][8]  ( .D(n14756), .SI(\mem1[30][15] ), .SE(test_se), 
        .CLK(n1560), .Q(\mem1[31][8] ), .QN(n27400) );
  SDFFX1 \mem1_reg[30][15]  ( .D(n14755), .SI(\mem1[30][14] ), .SE(test_se), 
        .CLK(n1560), .Q(\mem1[30][15] ), .QN(n27401) );
  SDFFX1 \mem1_reg[30][14]  ( .D(n14754), .SI(\mem1[30][13] ), .SE(test_se), 
        .CLK(n1560), .Q(\mem1[30][14] ), .QN(n27402) );
  SDFFX1 \mem1_reg[30][13]  ( .D(n14753), .SI(\mem1[30][12] ), .SE(test_se), 
        .CLK(n1560), .Q(\mem1[30][13] ), .QN(n27403) );
  SDFFX1 \mem1_reg[30][12]  ( .D(n14752), .SI(\mem1[30][11] ), .SE(test_se), 
        .CLK(n1560), .Q(\mem1[30][12] ), .QN(n27404) );
  SDFFX1 \mem1_reg[30][11]  ( .D(n14751), .SI(\mem1[30][10] ), .SE(test_se), 
        .CLK(n1560), .Q(\mem1[30][11] ), .QN(n27405) );
  SDFFX1 \mem1_reg[30][10]  ( .D(n14750), .SI(\mem1[30][9] ), .SE(test_se), 
        .CLK(n1560), .Q(\mem1[30][10] ), .QN(n27406) );
  SDFFX1 \mem1_reg[30][9]  ( .D(n14749), .SI(\mem1[30][8] ), .SE(test_se), 
        .CLK(n1561), .Q(\mem1[30][9] ), .QN(n27407) );
  SDFFX1 \mem1_reg[30][8]  ( .D(n14748), .SI(\mem1[29][15] ), .SE(test_se), 
        .CLK(n1561), .Q(\mem1[30][8] ), .QN(n27408) );
  SDFFX1 \mem1_reg[29][15]  ( .D(n14747), .SI(\mem1[29][14] ), .SE(test_se), 
        .CLK(n1561), .Q(\mem1[29][15] ), .QN(n27409) );
  SDFFX1 \mem1_reg[29][14]  ( .D(n14746), .SI(\mem1[29][13] ), .SE(test_se), 
        .CLK(n1561), .Q(\mem1[29][14] ), .QN(n27410) );
  SDFFX1 \mem1_reg[29][13]  ( .D(n14745), .SI(\mem1[29][12] ), .SE(test_se), 
        .CLK(n1561), .Q(\mem1[29][13] ), .QN(n27411) );
  SDFFX1 \mem1_reg[29][12]  ( .D(n14744), .SI(\mem1[29][11] ), .SE(test_se), 
        .CLK(n1561), .Q(\mem1[29][12] ), .QN(n27412) );
  SDFFX1 \mem1_reg[29][11]  ( .D(n14743), .SI(\mem1[29][10] ), .SE(test_se), 
        .CLK(n1561), .Q(\mem1[29][11] ), .QN(n27413) );
  SDFFX1 \mem1_reg[29][10]  ( .D(n14742), .SI(\mem1[29][9] ), .SE(test_se), 
        .CLK(n1561), .Q(\mem1[29][10] ), .QN(n27414) );
  SDFFX1 \mem1_reg[29][9]  ( .D(n14741), .SI(\mem1[29][8] ), .SE(test_se), 
        .CLK(n1561), .Q(\mem1[29][9] ), .QN(n27415) );
  SDFFX1 \mem1_reg[29][8]  ( .D(n14740), .SI(\mem1[28][15] ), .SE(test_se), 
        .CLK(n1561), .Q(\mem1[29][8] ), .QN(n27416) );
  SDFFX1 \mem1_reg[28][15]  ( .D(n14739), .SI(\mem1[28][14] ), .SE(test_se), 
        .CLK(n1561), .Q(\mem1[28][15] ), .QN(n27417) );
  SDFFX1 \mem1_reg[28][14]  ( .D(n14738), .SI(\mem1[28][13] ), .SE(test_se), 
        .CLK(n1561), .Q(\mem1[28][14] ), .QN(n27418) );
  SDFFX1 \mem1_reg[28][13]  ( .D(n14737), .SI(\mem1[28][12] ), .SE(test_se), 
        .CLK(n1562), .Q(\mem1[28][13] ), .QN(n27419) );
  SDFFX1 \mem1_reg[28][12]  ( .D(n14736), .SI(\mem1[28][11] ), .SE(test_se), 
        .CLK(n1562), .Q(\mem1[28][12] ), .QN(n27420) );
  SDFFX1 \mem1_reg[28][11]  ( .D(n14735), .SI(\mem1[28][10] ), .SE(test_se), 
        .CLK(n1562), .Q(\mem1[28][11] ), .QN(n27421) );
  SDFFX1 \mem1_reg[28][10]  ( .D(n14734), .SI(\mem1[28][9] ), .SE(test_se), 
        .CLK(n1562), .Q(\mem1[28][10] ), .QN(n27422) );
  SDFFX1 \mem1_reg[28][9]  ( .D(n14733), .SI(\mem1[28][8] ), .SE(test_se), 
        .CLK(n1562), .Q(\mem1[28][9] ), .QN(n27423) );
  SDFFX1 \mem1_reg[28][8]  ( .D(n14732), .SI(\mem1[27][15] ), .SE(test_se), 
        .CLK(n1562), .Q(\mem1[28][8] ), .QN(n27424) );
  SDFFX1 \mem1_reg[27][15]  ( .D(n14731), .SI(\mem1[27][14] ), .SE(test_se), 
        .CLK(n1562), .Q(\mem1[27][15] ), .QN(n27425) );
  SDFFX1 \mem1_reg[27][14]  ( .D(n14730), .SI(\mem1[27][13] ), .SE(test_se), 
        .CLK(n1562), .Q(\mem1[27][14] ), .QN(n27426) );
  SDFFX1 \mem1_reg[27][13]  ( .D(n14729), .SI(\mem1[27][12] ), .SE(test_se), 
        .CLK(n1562), .Q(\mem1[27][13] ), .QN(n27427) );
  SDFFX1 \mem1_reg[27][12]  ( .D(n14728), .SI(\mem1[27][11] ), .SE(test_se), 
        .CLK(n1562), .Q(\mem1[27][12] ), .QN(n27428) );
  SDFFX1 \mem1_reg[27][11]  ( .D(n14727), .SI(\mem1[27][10] ), .SE(test_se), 
        .CLK(n1562), .Q(\mem1[27][11] ), .QN(n27429) );
  SDFFX1 \mem1_reg[27][10]  ( .D(n14726), .SI(\mem1[27][9] ), .SE(test_se), 
        .CLK(n1562), .Q(\mem1[27][10] ), .QN(n27430) );
  SDFFX1 \mem1_reg[27][9]  ( .D(n14725), .SI(\mem1[27][8] ), .SE(test_se), 
        .CLK(n1563), .Q(\mem1[27][9] ), .QN(n27431) );
  SDFFX1 \mem1_reg[27][8]  ( .D(n14724), .SI(\mem1[26][15] ), .SE(test_se), 
        .CLK(n1563), .Q(\mem1[27][8] ), .QN(n27432) );
  SDFFX1 \mem1_reg[26][15]  ( .D(n14723), .SI(\mem1[26][14] ), .SE(test_se), 
        .CLK(n1563), .Q(\mem1[26][15] ), .QN(n27433) );
  SDFFX1 \mem1_reg[26][14]  ( .D(n14722), .SI(\mem1[26][13] ), .SE(test_se), 
        .CLK(n1563), .Q(\mem1[26][14] ), .QN(n27434) );
  SDFFX1 \mem1_reg[26][13]  ( .D(n14721), .SI(\mem1[26][12] ), .SE(test_se), 
        .CLK(n1563), .Q(\mem1[26][13] ), .QN(n27435) );
  SDFFX1 \mem1_reg[26][12]  ( .D(n14720), .SI(\mem1[26][11] ), .SE(test_se), 
        .CLK(n1563), .Q(\mem1[26][12] ), .QN(n27436) );
  SDFFX1 \mem1_reg[26][11]  ( .D(n14719), .SI(\mem1[26][10] ), .SE(test_se), 
        .CLK(n1563), .Q(\mem1[26][11] ), .QN(n27437) );
  SDFFX1 \mem1_reg[26][10]  ( .D(n14718), .SI(\mem1[26][9] ), .SE(test_se), 
        .CLK(n1563), .Q(\mem1[26][10] ), .QN(n27438) );
  SDFFX1 \mem1_reg[26][9]  ( .D(n14717), .SI(\mem1[26][8] ), .SE(test_se), 
        .CLK(n1563), .Q(\mem1[26][9] ), .QN(n27439) );
  SDFFX1 \mem1_reg[26][8]  ( .D(n14716), .SI(\mem1[25][15] ), .SE(test_se), 
        .CLK(n1563), .Q(\mem1[26][8] ), .QN(n27440) );
  SDFFX1 \mem1_reg[25][15]  ( .D(n14715), .SI(\mem1[25][14] ), .SE(test_se), 
        .CLK(n1563), .Q(\mem1[25][15] ), .QN(n27441) );
  SDFFX1 \mem1_reg[25][14]  ( .D(n14714), .SI(\mem1[25][13] ), .SE(test_se), 
        .CLK(n1563), .Q(\mem1[25][14] ), .QN(n27442) );
  SDFFX1 \mem1_reg[25][13]  ( .D(n14713), .SI(\mem1[25][12] ), .SE(test_se), 
        .CLK(n1564), .Q(\mem1[25][13] ), .QN(n27443) );
  SDFFX1 \mem1_reg[25][12]  ( .D(n14712), .SI(\mem1[25][11] ), .SE(test_se), 
        .CLK(n1564), .Q(\mem1[25][12] ), .QN(n27444) );
  SDFFX1 \mem1_reg[25][11]  ( .D(n14711), .SI(\mem1[25][10] ), .SE(test_se), 
        .CLK(n1564), .Q(\mem1[25][11] ), .QN(n27445) );
  SDFFX1 \mem1_reg[25][10]  ( .D(n14710), .SI(\mem1[25][9] ), .SE(test_se), 
        .CLK(n1564), .Q(\mem1[25][10] ), .QN(n27446) );
  SDFFX1 \mem1_reg[25][9]  ( .D(n14709), .SI(\mem1[25][8] ), .SE(test_se), 
        .CLK(n1564), .Q(\mem1[25][9] ), .QN(n27447) );
  SDFFX1 \mem1_reg[25][8]  ( .D(n14708), .SI(\mem1[24][15] ), .SE(test_se), 
        .CLK(n1564), .Q(\mem1[25][8] ), .QN(n27448) );
  SDFFX1 \mem1_reg[24][15]  ( .D(n14707), .SI(\mem1[24][14] ), .SE(test_se), 
        .CLK(n1564), .Q(\mem1[24][15] ), .QN(n27449) );
  SDFFX1 \mem1_reg[24][14]  ( .D(n14706), .SI(\mem1[24][13] ), .SE(test_se), 
        .CLK(n1564), .Q(\mem1[24][14] ), .QN(n27450) );
  SDFFX1 \mem1_reg[24][13]  ( .D(n14705), .SI(\mem1[24][12] ), .SE(test_se), 
        .CLK(n1564), .Q(\mem1[24][13] ), .QN(n27451) );
  SDFFX1 \mem1_reg[24][12]  ( .D(n14704), .SI(\mem1[24][11] ), .SE(test_se), 
        .CLK(n1564), .Q(\mem1[24][12] ), .QN(n27452) );
  SDFFX1 \mem1_reg[24][11]  ( .D(n14703), .SI(\mem1[24][10] ), .SE(test_se), 
        .CLK(n1564), .Q(\mem1[24][11] ), .QN(n27453) );
  SDFFX1 \mem1_reg[24][10]  ( .D(n14702), .SI(\mem1[24][9] ), .SE(test_se), 
        .CLK(n1564), .Q(\mem1[24][10] ), .QN(n27454) );
  SDFFX1 \mem1_reg[24][9]  ( .D(n14701), .SI(\mem1[24][8] ), .SE(test_se), 
        .CLK(n1565), .Q(\mem1[24][9] ), .QN(n27455) );
  SDFFX1 \mem1_reg[24][8]  ( .D(n14700), .SI(\mem1[23][15] ), .SE(test_se), 
        .CLK(n1565), .Q(\mem1[24][8] ), .QN(n27456) );
  SDFFX1 \mem1_reg[23][15]  ( .D(n14699), .SI(\mem1[23][14] ), .SE(test_se), 
        .CLK(n1565), .Q(\mem1[23][15] ), .QN(n27457) );
  SDFFX1 \mem1_reg[23][14]  ( .D(n14698), .SI(\mem1[23][13] ), .SE(test_se), 
        .CLK(n1565), .Q(\mem1[23][14] ), .QN(n27458) );
  SDFFX1 \mem1_reg[23][13]  ( .D(n14697), .SI(\mem1[23][12] ), .SE(test_se), 
        .CLK(n1565), .Q(\mem1[23][13] ), .QN(n27459) );
  SDFFX1 \mem1_reg[23][12]  ( .D(n14696), .SI(\mem1[23][11] ), .SE(test_se), 
        .CLK(n1565), .Q(\mem1[23][12] ), .QN(n27460) );
  SDFFX1 \mem1_reg[23][11]  ( .D(n14695), .SI(\mem1[23][10] ), .SE(test_se), 
        .CLK(n1565), .Q(\mem1[23][11] ), .QN(n27461) );
  SDFFX1 \mem1_reg[23][10]  ( .D(n14694), .SI(\mem1[23][9] ), .SE(test_se), 
        .CLK(n1565), .Q(\mem1[23][10] ), .QN(n27462) );
  SDFFX1 \mem1_reg[23][9]  ( .D(n14693), .SI(\mem1[23][8] ), .SE(test_se), 
        .CLK(n1565), .Q(\mem1[23][9] ), .QN(n27463) );
  SDFFX1 \mem1_reg[23][8]  ( .D(n14692), .SI(\mem1[22][15] ), .SE(test_se), 
        .CLK(n1565), .Q(\mem1[23][8] ), .QN(n27464) );
  SDFFX1 \mem1_reg[22][15]  ( .D(n14691), .SI(\mem1[22][14] ), .SE(test_se), 
        .CLK(n1565), .Q(\mem1[22][15] ), .QN(n27465) );
  SDFFX1 \mem1_reg[22][14]  ( .D(n14690), .SI(\mem1[22][13] ), .SE(test_se), 
        .CLK(n1565), .Q(\mem1[22][14] ), .QN(n27466) );
  SDFFX1 \mem1_reg[22][13]  ( .D(n14689), .SI(\mem1[22][12] ), .SE(test_se), 
        .CLK(n1566), .Q(\mem1[22][13] ), .QN(n27467) );
  SDFFX1 \mem1_reg[22][12]  ( .D(n14688), .SI(\mem1[22][11] ), .SE(test_se), 
        .CLK(n1566), .Q(\mem1[22][12] ), .QN(n27468) );
  SDFFX1 \mem1_reg[22][11]  ( .D(n14687), .SI(\mem1[22][10] ), .SE(test_se), 
        .CLK(n1566), .Q(\mem1[22][11] ), .QN(n27469) );
  SDFFX1 \mem1_reg[22][10]  ( .D(n14686), .SI(\mem1[22][9] ), .SE(test_se), 
        .CLK(n1566), .Q(\mem1[22][10] ), .QN(n27470) );
  SDFFX1 \mem1_reg[22][9]  ( .D(n14685), .SI(\mem1[22][8] ), .SE(test_se), 
        .CLK(n1566), .Q(\mem1[22][9] ), .QN(n27471) );
  SDFFX1 \mem1_reg[22][8]  ( .D(n14684), .SI(\mem1[21][15] ), .SE(test_se), 
        .CLK(n1566), .Q(\mem1[22][8] ), .QN(n27472) );
  SDFFX1 \mem1_reg[21][15]  ( .D(n14683), .SI(\mem1[21][14] ), .SE(test_se), 
        .CLK(n1566), .Q(\mem1[21][15] ), .QN(n27473) );
  SDFFX1 \mem1_reg[21][14]  ( .D(n14682), .SI(\mem1[21][13] ), .SE(test_se), 
        .CLK(n1566), .Q(\mem1[21][14] ), .QN(n27474) );
  SDFFX1 \mem1_reg[21][13]  ( .D(n14681), .SI(\mem1[21][12] ), .SE(test_se), 
        .CLK(n1566), .Q(\mem1[21][13] ), .QN(n27475) );
  SDFFX1 \mem1_reg[21][12]  ( .D(n14680), .SI(\mem1[21][11] ), .SE(test_se), 
        .CLK(n1566), .Q(\mem1[21][12] ), .QN(n27476) );
  SDFFX1 \mem1_reg[21][11]  ( .D(n14679), .SI(\mem1[21][10] ), .SE(test_se), 
        .CLK(n1566), .Q(\mem1[21][11] ), .QN(n27477) );
  SDFFX1 \mem1_reg[21][10]  ( .D(n14678), .SI(\mem1[21][9] ), .SE(test_se), 
        .CLK(n1566), .Q(\mem1[21][10] ), .QN(n27478) );
  SDFFX1 \mem1_reg[21][9]  ( .D(n14677), .SI(\mem1[21][8] ), .SE(test_se), 
        .CLK(n1567), .Q(\mem1[21][9] ), .QN(n27479) );
  SDFFX1 \mem1_reg[21][8]  ( .D(n14676), .SI(\mem1[20][15] ), .SE(test_se), 
        .CLK(n1567), .Q(\mem1[21][8] ), .QN(n27480) );
  SDFFX1 \mem1_reg[20][15]  ( .D(n14675), .SI(\mem1[20][14] ), .SE(test_se), 
        .CLK(n1567), .Q(\mem1[20][15] ), .QN(n27481) );
  SDFFX1 \mem1_reg[20][14]  ( .D(n14674), .SI(\mem1[20][13] ), .SE(test_se), 
        .CLK(n1567), .Q(\mem1[20][14] ), .QN(n27482) );
  SDFFX1 \mem1_reg[20][13]  ( .D(n14673), .SI(\mem1[20][12] ), .SE(test_se), 
        .CLK(n1567), .Q(\mem1[20][13] ), .QN(n27483) );
  SDFFX1 \mem1_reg[20][12]  ( .D(n14672), .SI(\mem1[20][11] ), .SE(test_se), 
        .CLK(n1567), .Q(\mem1[20][12] ), .QN(n27484) );
  SDFFX1 \mem1_reg[20][11]  ( .D(n14671), .SI(\mem1[20][10] ), .SE(test_se), 
        .CLK(n1567), .Q(\mem1[20][11] ), .QN(n27485) );
  SDFFX1 \mem1_reg[20][10]  ( .D(n14670), .SI(\mem1[20][9] ), .SE(test_se), 
        .CLK(n1567), .Q(\mem1[20][10] ), .QN(n27486) );
  SDFFX1 \mem1_reg[20][9]  ( .D(n14669), .SI(\mem1[20][8] ), .SE(test_se), 
        .CLK(n1567), .Q(\mem1[20][9] ), .QN(n27487) );
  SDFFX1 \mem1_reg[20][8]  ( .D(n14668), .SI(\mem1[19][15] ), .SE(test_se), 
        .CLK(n1567), .Q(\mem1[20][8] ), .QN(n27488) );
  SDFFX1 \mem1_reg[19][15]  ( .D(n14667), .SI(\mem1[19][14] ), .SE(test_se), 
        .CLK(n1567), .Q(\mem1[19][15] ), .QN(n27489) );
  SDFFX1 \mem1_reg[19][14]  ( .D(n14666), .SI(\mem1[19][13] ), .SE(test_se), 
        .CLK(n1567), .Q(\mem1[19][14] ), .QN(n27490) );
  SDFFX1 \mem1_reg[19][13]  ( .D(n14665), .SI(\mem1[19][12] ), .SE(test_se), 
        .CLK(n1568), .Q(\mem1[19][13] ), .QN(n27491) );
  SDFFX1 \mem1_reg[19][12]  ( .D(n14664), .SI(\mem1[19][11] ), .SE(test_se), 
        .CLK(n1568), .Q(\mem1[19][12] ), .QN(n27492) );
  SDFFX1 \mem1_reg[19][11]  ( .D(n14663), .SI(\mem1[19][10] ), .SE(test_se), 
        .CLK(n1568), .Q(\mem1[19][11] ), .QN(n27493) );
  SDFFX1 \mem1_reg[19][10]  ( .D(n14662), .SI(\mem1[19][9] ), .SE(test_se), 
        .CLK(n1568), .Q(\mem1[19][10] ), .QN(n27494) );
  SDFFX1 \mem1_reg[19][9]  ( .D(n14661), .SI(\mem1[19][8] ), .SE(test_se), 
        .CLK(n1568), .Q(\mem1[19][9] ), .QN(n27495) );
  SDFFX1 \mem1_reg[19][8]  ( .D(n14660), .SI(\mem1[18][15] ), .SE(test_se), 
        .CLK(n1568), .Q(\mem1[19][8] ), .QN(n27496) );
  SDFFX1 \mem1_reg[18][15]  ( .D(n14659), .SI(\mem1[18][14] ), .SE(test_se), 
        .CLK(n1568), .Q(\mem1[18][15] ), .QN(n27497) );
  SDFFX1 \mem1_reg[18][14]  ( .D(n14658), .SI(\mem1[18][13] ), .SE(test_se), 
        .CLK(n1568), .Q(\mem1[18][14] ), .QN(n27498) );
  SDFFX1 \mem1_reg[18][13]  ( .D(n14657), .SI(\mem1[18][12] ), .SE(test_se), 
        .CLK(n1568), .Q(\mem1[18][13] ), .QN(n27499) );
  SDFFX1 \mem1_reg[18][12]  ( .D(n14656), .SI(\mem1[18][11] ), .SE(test_se), 
        .CLK(n1568), .Q(\mem1[18][12] ), .QN(n27500) );
  SDFFX1 \mem1_reg[18][11]  ( .D(n14655), .SI(\mem1[18][10] ), .SE(test_se), 
        .CLK(n1568), .Q(\mem1[18][11] ), .QN(n27501) );
  SDFFX1 \mem1_reg[18][10]  ( .D(n14654), .SI(\mem1[18][9] ), .SE(test_se), 
        .CLK(n1568), .Q(\mem1[18][10] ), .QN(n27502) );
  SDFFX1 \mem1_reg[18][9]  ( .D(n14653), .SI(\mem1[18][8] ), .SE(test_se), 
        .CLK(n1569), .Q(\mem1[18][9] ), .QN(n27503) );
  SDFFX1 \mem1_reg[18][8]  ( .D(n14652), .SI(\mem1[17][15] ), .SE(test_se), 
        .CLK(n1569), .Q(\mem1[18][8] ), .QN(n27504) );
  SDFFX1 \mem1_reg[17][15]  ( .D(n14651), .SI(\mem1[17][14] ), .SE(test_se), 
        .CLK(n1569), .Q(\mem1[17][15] ), .QN(n27505) );
  SDFFX1 \mem1_reg[17][14]  ( .D(n14650), .SI(\mem1[17][13] ), .SE(test_se), 
        .CLK(n1569), .Q(\mem1[17][14] ), .QN(n27506) );
  SDFFX1 \mem1_reg[17][13]  ( .D(n14649), .SI(\mem1[17][12] ), .SE(test_se), 
        .CLK(n1569), .Q(\mem1[17][13] ), .QN(n27507) );
  SDFFX1 \mem1_reg[17][12]  ( .D(n14648), .SI(\mem1[17][11] ), .SE(test_se), 
        .CLK(n1569), .Q(\mem1[17][12] ), .QN(n27508) );
  SDFFX1 \mem1_reg[17][11]  ( .D(n14647), .SI(\mem1[17][10] ), .SE(test_se), 
        .CLK(n1569), .Q(\mem1[17][11] ), .QN(n27509) );
  SDFFX1 \mem1_reg[17][10]  ( .D(n14646), .SI(\mem1[17][9] ), .SE(test_se), 
        .CLK(n1569), .Q(\mem1[17][10] ), .QN(n27510) );
  SDFFX1 \mem1_reg[17][9]  ( .D(n14645), .SI(\mem1[17][8] ), .SE(test_se), 
        .CLK(n1569), .Q(\mem1[17][9] ), .QN(n27511) );
  SDFFX1 \mem1_reg[17][8]  ( .D(n14644), .SI(\mem1[16][15] ), .SE(test_se), 
        .CLK(n1569), .Q(\mem1[17][8] ), .QN(n27512) );
  SDFFX1 \mem1_reg[16][15]  ( .D(n14643), .SI(\mem1[16][14] ), .SE(test_se), 
        .CLK(n1569), .Q(\mem1[16][15] ), .QN(n27513) );
  SDFFX1 \mem1_reg[16][14]  ( .D(n14642), .SI(\mem1[16][13] ), .SE(test_se), 
        .CLK(n1569), .Q(\mem1[16][14] ), .QN(n27514) );
  SDFFX1 \mem1_reg[16][13]  ( .D(n14641), .SI(\mem1[16][12] ), .SE(test_se), 
        .CLK(n1570), .Q(\mem1[16][13] ), .QN(n27515) );
  SDFFX1 \mem1_reg[16][12]  ( .D(n14640), .SI(\mem1[16][11] ), .SE(test_se), 
        .CLK(n1570), .Q(\mem1[16][12] ), .QN(n27516) );
  SDFFX1 \mem1_reg[16][11]  ( .D(n14639), .SI(\mem1[16][10] ), .SE(test_se), 
        .CLK(n1570), .Q(\mem1[16][11] ), .QN(n27517) );
  SDFFX1 \mem1_reg[16][10]  ( .D(n14638), .SI(\mem1[16][9] ), .SE(test_se), 
        .CLK(n1570), .Q(\mem1[16][10] ), .QN(n27518) );
  SDFFX1 \mem1_reg[16][9]  ( .D(n14637), .SI(\mem1[16][8] ), .SE(test_se), 
        .CLK(n1570), .Q(\mem1[16][9] ), .QN(n27519) );
  SDFFX1 \mem1_reg[16][8]  ( .D(n14636), .SI(\mem1[15][15] ), .SE(test_se), 
        .CLK(n1570), .Q(\mem1[16][8] ), .QN(n27520) );
  SDFFX1 \mem1_reg[15][15]  ( .D(n14635), .SI(\mem1[15][14] ), .SE(test_se), 
        .CLK(n1570), .Q(\mem1[15][15] ), .QN(n27521) );
  SDFFX1 \mem1_reg[15][14]  ( .D(n14634), .SI(\mem1[15][13] ), .SE(test_se), 
        .CLK(n1570), .Q(\mem1[15][14] ), .QN(n27522) );
  SDFFX1 \mem1_reg[15][13]  ( .D(n14633), .SI(\mem1[15][12] ), .SE(test_se), 
        .CLK(n1570), .Q(\mem1[15][13] ), .QN(n27523) );
  SDFFX1 \mem1_reg[15][12]  ( .D(n14632), .SI(\mem1[15][11] ), .SE(test_se), 
        .CLK(n1570), .Q(\mem1[15][12] ), .QN(n27524) );
  SDFFX1 \mem1_reg[15][11]  ( .D(n14631), .SI(\mem1[15][10] ), .SE(test_se), 
        .CLK(n1570), .Q(\mem1[15][11] ), .QN(n27525) );
  SDFFX1 \mem1_reg[15][10]  ( .D(n14630), .SI(\mem1[15][9] ), .SE(test_se), 
        .CLK(n1570), .Q(\mem1[15][10] ), .QN(n27526) );
  SDFFX1 \mem1_reg[15][9]  ( .D(n14629), .SI(\mem1[15][8] ), .SE(test_se), 
        .CLK(n1571), .Q(\mem1[15][9] ), .QN(n27527) );
  SDFFX1 \mem1_reg[15][8]  ( .D(n14628), .SI(\mem1[14][15] ), .SE(test_se), 
        .CLK(n1571), .Q(\mem1[15][8] ), .QN(n27528) );
  SDFFX1 \mem1_reg[14][15]  ( .D(n14627), .SI(\mem1[14][14] ), .SE(test_se), 
        .CLK(n1571), .Q(\mem1[14][15] ), .QN(n27529) );
  SDFFX1 \mem1_reg[14][14]  ( .D(n14626), .SI(\mem1[14][13] ), .SE(test_se), 
        .CLK(n1571), .Q(\mem1[14][14] ), .QN(n27530) );
  SDFFX1 \mem1_reg[14][13]  ( .D(n14625), .SI(\mem1[14][12] ), .SE(test_se), 
        .CLK(n1571), .Q(\mem1[14][13] ), .QN(n27531) );
  SDFFX1 \mem1_reg[14][12]  ( .D(n14624), .SI(\mem1[14][11] ), .SE(test_se), 
        .CLK(n1571), .Q(\mem1[14][12] ), .QN(n27532) );
  SDFFX1 \mem1_reg[14][11]  ( .D(n14623), .SI(\mem1[14][10] ), .SE(test_se), 
        .CLK(n1571), .Q(\mem1[14][11] ), .QN(n27533) );
  SDFFX1 \mem1_reg[14][10]  ( .D(n14622), .SI(\mem1[14][9] ), .SE(test_se), 
        .CLK(n1571), .Q(\mem1[14][10] ), .QN(n27534) );
  SDFFX1 \mem1_reg[14][9]  ( .D(n14621), .SI(\mem1[14][8] ), .SE(test_se), 
        .CLK(n1571), .Q(\mem1[14][9] ), .QN(n27535) );
  SDFFX1 \mem1_reg[14][8]  ( .D(n14620), .SI(\mem1[13][15] ), .SE(test_se), 
        .CLK(n1571), .Q(\mem1[14][8] ), .QN(n27536) );
  SDFFX1 \mem1_reg[13][15]  ( .D(n14619), .SI(\mem1[13][14] ), .SE(test_se), 
        .CLK(n1571), .Q(\mem1[13][15] ), .QN(n27537) );
  SDFFX1 \mem1_reg[13][14]  ( .D(n14618), .SI(\mem1[13][13] ), .SE(test_se), 
        .CLK(n1571), .Q(\mem1[13][14] ), .QN(n27538) );
  SDFFX1 \mem1_reg[13][13]  ( .D(n14617), .SI(\mem1[13][12] ), .SE(test_se), 
        .CLK(n1572), .Q(\mem1[13][13] ), .QN(n27539) );
  SDFFX1 \mem1_reg[13][12]  ( .D(n14616), .SI(\mem1[13][11] ), .SE(test_se), 
        .CLK(n1572), .Q(\mem1[13][12] ), .QN(n27540) );
  SDFFX1 \mem1_reg[13][11]  ( .D(n14615), .SI(\mem1[13][10] ), .SE(test_se), 
        .CLK(n1572), .Q(\mem1[13][11] ), .QN(n27541) );
  SDFFX1 \mem1_reg[13][10]  ( .D(n14614), .SI(\mem1[13][9] ), .SE(test_se), 
        .CLK(n1572), .Q(\mem1[13][10] ), .QN(n27542) );
  SDFFX1 \mem1_reg[13][9]  ( .D(n14613), .SI(\mem1[13][8] ), .SE(test_se), 
        .CLK(n1572), .Q(\mem1[13][9] ), .QN(n27543) );
  SDFFX1 \mem1_reg[13][8]  ( .D(n14612), .SI(\mem1[12][15] ), .SE(test_se), 
        .CLK(n1572), .Q(\mem1[13][8] ), .QN(n27544) );
  SDFFX1 \mem1_reg[12][15]  ( .D(n14611), .SI(\mem1[12][14] ), .SE(test_se), 
        .CLK(n1572), .Q(\mem1[12][15] ), .QN(n27545) );
  SDFFX1 \mem1_reg[12][14]  ( .D(n14610), .SI(\mem1[12][13] ), .SE(test_se), 
        .CLK(n1572), .Q(\mem1[12][14] ), .QN(n27546) );
  SDFFX1 \mem1_reg[12][13]  ( .D(n14609), .SI(\mem1[12][12] ), .SE(test_se), 
        .CLK(n1572), .Q(\mem1[12][13] ), .QN(n27547) );
  SDFFX1 \mem1_reg[12][12]  ( .D(n14608), .SI(\mem1[12][11] ), .SE(test_se), 
        .CLK(n1572), .Q(\mem1[12][12] ), .QN(n27548) );
  SDFFX1 \mem1_reg[12][11]  ( .D(n14607), .SI(\mem1[12][10] ), .SE(test_se), 
        .CLK(n1572), .Q(\mem1[12][11] ), .QN(n27549) );
  SDFFX1 \mem1_reg[12][10]  ( .D(n14606), .SI(\mem1[12][9] ), .SE(test_se), 
        .CLK(n1572), .Q(\mem1[12][10] ), .QN(n27550) );
  SDFFX1 \mem1_reg[12][9]  ( .D(n14605), .SI(\mem1[12][8] ), .SE(test_se), 
        .CLK(n1573), .Q(\mem1[12][9] ), .QN(n27551) );
  SDFFX1 \mem1_reg[12][8]  ( .D(n14604), .SI(\mem1[11][15] ), .SE(test_se), 
        .CLK(n1573), .Q(\mem1[12][8] ), .QN(n27552) );
  SDFFX1 \mem1_reg[11][15]  ( .D(n14603), .SI(\mem1[11][14] ), .SE(test_se), 
        .CLK(n1573), .Q(\mem1[11][15] ), .QN(n27553) );
  SDFFX1 \mem1_reg[11][14]  ( .D(n14602), .SI(\mem1[11][13] ), .SE(test_se), 
        .CLK(n1573), .Q(\mem1[11][14] ), .QN(n27554) );
  SDFFX1 \mem1_reg[11][13]  ( .D(n14601), .SI(\mem1[11][12] ), .SE(test_se), 
        .CLK(n1573), .Q(\mem1[11][13] ), .QN(n27555) );
  SDFFX1 \mem1_reg[11][12]  ( .D(n14600), .SI(\mem1[11][11] ), .SE(test_se), 
        .CLK(n1573), .Q(\mem1[11][12] ), .QN(n27556) );
  SDFFX1 \mem1_reg[11][11]  ( .D(n14599), .SI(\mem1[11][10] ), .SE(test_se), 
        .CLK(n1573), .Q(\mem1[11][11] ), .QN(n27557) );
  SDFFX1 \mem1_reg[11][10]  ( .D(n14598), .SI(\mem1[11][9] ), .SE(test_se), 
        .CLK(n1573), .Q(\mem1[11][10] ), .QN(n27558) );
  SDFFX1 \mem1_reg[11][9]  ( .D(n14597), .SI(\mem1[11][8] ), .SE(test_se), 
        .CLK(n1573), .Q(\mem1[11][9] ), .QN(n27559) );
  SDFFX1 \mem1_reg[11][8]  ( .D(n14596), .SI(\mem1[10][15] ), .SE(test_se), 
        .CLK(n1573), .Q(\mem1[11][8] ), .QN(n27560) );
  SDFFX1 \mem1_reg[10][15]  ( .D(n14595), .SI(\mem1[10][14] ), .SE(test_se), 
        .CLK(n1573), .Q(\mem1[10][15] ), .QN(n27561) );
  SDFFX1 \mem1_reg[10][14]  ( .D(n14594), .SI(\mem1[10][13] ), .SE(test_se), 
        .CLK(n1573), .Q(\mem1[10][14] ), .QN(n27562) );
  SDFFX1 \mem1_reg[10][13]  ( .D(n14593), .SI(\mem1[10][12] ), .SE(test_se), 
        .CLK(n1574), .Q(\mem1[10][13] ), .QN(n27563) );
  SDFFX1 \mem1_reg[10][12]  ( .D(n14592), .SI(\mem1[10][11] ), .SE(test_se), 
        .CLK(n1574), .Q(\mem1[10][12] ), .QN(n27564) );
  SDFFX1 \mem1_reg[10][11]  ( .D(n14591), .SI(\mem1[10][10] ), .SE(test_se), 
        .CLK(n1574), .Q(\mem1[10][11] ), .QN(n27565) );
  SDFFX1 \mem1_reg[10][10]  ( .D(n14590), .SI(\mem1[10][9] ), .SE(test_se), 
        .CLK(n1574), .Q(\mem1[10][10] ), .QN(n27566) );
  SDFFX1 \mem1_reg[10][9]  ( .D(n14589), .SI(\mem1[10][8] ), .SE(test_se), 
        .CLK(n1574), .Q(\mem1[10][9] ), .QN(n27567) );
  SDFFX1 \mem1_reg[10][8]  ( .D(n14588), .SI(\mem1[9][15] ), .SE(test_se), 
        .CLK(n1574), .Q(\mem1[10][8] ), .QN(n27568) );
  SDFFX1 \mem1_reg[9][15]  ( .D(n14587), .SI(\mem1[9][14] ), .SE(test_se), 
        .CLK(n1574), .Q(\mem1[9][15] ), .QN(n27569) );
  SDFFX1 \mem1_reg[9][14]  ( .D(n14586), .SI(\mem1[9][13] ), .SE(test_se), 
        .CLK(n1574), .Q(\mem1[9][14] ), .QN(n27570) );
  SDFFX1 \mem1_reg[9][13]  ( .D(n14585), .SI(\mem1[9][12] ), .SE(test_se), 
        .CLK(n1574), .Q(\mem1[9][13] ), .QN(n27571) );
  SDFFX1 \mem1_reg[9][12]  ( .D(n14584), .SI(\mem1[9][11] ), .SE(test_se), 
        .CLK(n1574), .Q(\mem1[9][12] ), .QN(n27572) );
  SDFFX1 \mem1_reg[9][11]  ( .D(n14583), .SI(\mem1[9][10] ), .SE(test_se), 
        .CLK(n1574), .Q(\mem1[9][11] ), .QN(n27573) );
  SDFFX1 \mem1_reg[9][10]  ( .D(n14582), .SI(\mem1[9][9] ), .SE(test_se), 
        .CLK(n1574), .Q(\mem1[9][10] ), .QN(n27574) );
  SDFFX1 \mem1_reg[9][9]  ( .D(n14581), .SI(\mem1[9][8] ), .SE(test_se), .CLK(
        n1575), .Q(\mem1[9][9] ), .QN(n27575) );
  SDFFX1 \mem1_reg[9][8]  ( .D(n14580), .SI(\mem1[8][15] ), .SE(test_se), 
        .CLK(n1575), .Q(\mem1[9][8] ), .QN(n27576) );
  SDFFX1 \mem1_reg[8][15]  ( .D(n14579), .SI(\mem1[8][14] ), .SE(test_se), 
        .CLK(n1575), .Q(\mem1[8][15] ), .QN(n27577) );
  SDFFX1 \mem1_reg[8][14]  ( .D(n14578), .SI(\mem1[8][13] ), .SE(test_se), 
        .CLK(n1575), .Q(\mem1[8][14] ), .QN(n27578) );
  SDFFX1 \mem1_reg[8][13]  ( .D(n14577), .SI(\mem1[8][12] ), .SE(test_se), 
        .CLK(n1575), .Q(\mem1[8][13] ), .QN(n27579) );
  SDFFX1 \mem1_reg[8][12]  ( .D(n14576), .SI(\mem1[8][11] ), .SE(test_se), 
        .CLK(n1575), .Q(\mem1[8][12] ), .QN(n27580) );
  SDFFX1 \mem1_reg[8][11]  ( .D(n14575), .SI(\mem1[8][10] ), .SE(test_se), 
        .CLK(n1575), .Q(\mem1[8][11] ), .QN(n27581) );
  SDFFX1 \mem1_reg[8][10]  ( .D(n14574), .SI(\mem1[8][9] ), .SE(test_se), 
        .CLK(n1575), .Q(\mem1[8][10] ), .QN(n27582) );
  SDFFX1 \mem1_reg[8][9]  ( .D(n14573), .SI(\mem1[8][8] ), .SE(test_se), .CLK(
        n1575), .Q(\mem1[8][9] ), .QN(n27583) );
  SDFFX1 \mem1_reg[8][8]  ( .D(n14572), .SI(\mem1[7][15] ), .SE(test_se), 
        .CLK(n1575), .Q(\mem1[8][8] ), .QN(n27584) );
  SDFFX1 \mem1_reg[7][15]  ( .D(n14571), .SI(\mem1[7][14] ), .SE(test_se), 
        .CLK(n1575), .Q(\mem1[7][15] ), .QN(n27585) );
  SDFFX1 \mem1_reg[7][14]  ( .D(n14570), .SI(\mem1[7][13] ), .SE(test_se), 
        .CLK(n1575), .Q(\mem1[7][14] ), .QN(n27586) );
  SDFFX1 \mem1_reg[7][13]  ( .D(n14569), .SI(\mem1[7][12] ), .SE(test_se), 
        .CLK(n1576), .Q(\mem1[7][13] ), .QN(n27587) );
  SDFFX1 \mem1_reg[7][12]  ( .D(n14568), .SI(\mem1[7][11] ), .SE(test_se), 
        .CLK(n1576), .Q(\mem1[7][12] ), .QN(n27588) );
  SDFFX1 \mem1_reg[7][11]  ( .D(n14567), .SI(\mem1[7][10] ), .SE(test_se), 
        .CLK(n1576), .Q(\mem1[7][11] ), .QN(n27589) );
  SDFFX1 \mem1_reg[7][10]  ( .D(n14566), .SI(\mem1[7][9] ), .SE(test_se), 
        .CLK(n1576), .Q(\mem1[7][10] ), .QN(n27590) );
  SDFFX1 \mem1_reg[7][9]  ( .D(n14565), .SI(\mem1[7][8] ), .SE(test_se), .CLK(
        n1576), .Q(\mem1[7][9] ), .QN(n27591) );
  SDFFX1 \mem1_reg[7][8]  ( .D(n14564), .SI(\mem1[6][15] ), .SE(test_se), 
        .CLK(n1576), .Q(\mem1[7][8] ), .QN(n27592) );
  SDFFX1 \mem1_reg[6][15]  ( .D(n14563), .SI(\mem1[6][14] ), .SE(test_se), 
        .CLK(n1576), .Q(\mem1[6][15] ), .QN(n27593) );
  SDFFX1 \mem1_reg[6][14]  ( .D(n14562), .SI(\mem1[6][13] ), .SE(test_se), 
        .CLK(n1576), .Q(\mem1[6][14] ), .QN(n27594) );
  SDFFX1 \mem1_reg[6][13]  ( .D(n14561), .SI(\mem1[6][12] ), .SE(test_se), 
        .CLK(n1576), .Q(\mem1[6][13] ), .QN(n27595) );
  SDFFX1 \mem1_reg[6][12]  ( .D(n14560), .SI(\mem1[6][11] ), .SE(test_se), 
        .CLK(n1576), .Q(\mem1[6][12] ), .QN(n27596) );
  SDFFX1 \mem1_reg[6][11]  ( .D(n14559), .SI(\mem1[6][10] ), .SE(test_se), 
        .CLK(n1576), .Q(\mem1[6][11] ), .QN(n27597) );
  SDFFX1 \mem1_reg[6][10]  ( .D(n14558), .SI(\mem1[6][9] ), .SE(test_se), 
        .CLK(n1576), .Q(\mem1[6][10] ), .QN(n27598) );
  SDFFX1 \mem1_reg[6][9]  ( .D(n14557), .SI(\mem1[6][8] ), .SE(test_se), .CLK(
        n1577), .Q(\mem1[6][9] ), .QN(n27599) );
  SDFFX1 \mem1_reg[6][8]  ( .D(n14556), .SI(\mem1[5][15] ), .SE(test_se), 
        .CLK(n1577), .Q(\mem1[6][8] ), .QN(n27600) );
  SDFFX1 \mem1_reg[5][15]  ( .D(n14555), .SI(\mem1[5][14] ), .SE(test_se), 
        .CLK(n1577), .Q(\mem1[5][15] ), .QN(n27601) );
  SDFFX1 \mem1_reg[5][14]  ( .D(n14554), .SI(\mem1[5][13] ), .SE(test_se), 
        .CLK(n1577), .Q(\mem1[5][14] ), .QN(n27602) );
  SDFFX1 \mem1_reg[5][13]  ( .D(n14553), .SI(\mem1[5][12] ), .SE(test_se), 
        .CLK(n1577), .Q(\mem1[5][13] ), .QN(n27603) );
  SDFFX1 \mem1_reg[5][12]  ( .D(n14552), .SI(\mem1[5][11] ), .SE(test_se), 
        .CLK(n1577), .Q(\mem1[5][12] ), .QN(n27604) );
  SDFFX1 \mem1_reg[5][11]  ( .D(n14551), .SI(\mem1[5][10] ), .SE(test_se), 
        .CLK(n1577), .Q(\mem1[5][11] ), .QN(n27605) );
  SDFFX1 \mem1_reg[5][10]  ( .D(n14550), .SI(\mem1[5][9] ), .SE(test_se), 
        .CLK(n1577), .Q(\mem1[5][10] ), .QN(n27606) );
  SDFFX1 \mem1_reg[5][9]  ( .D(n14549), .SI(\mem1[5][8] ), .SE(test_se), .CLK(
        n1577), .Q(\mem1[5][9] ), .QN(n27607) );
  SDFFX1 \mem1_reg[5][8]  ( .D(n14548), .SI(\mem1[4][15] ), .SE(test_se), 
        .CLK(n1577), .Q(\mem1[5][8] ), .QN(n27608) );
  SDFFX1 \mem1_reg[4][15]  ( .D(n14547), .SI(\mem1[4][14] ), .SE(test_se), 
        .CLK(n1577), .Q(\mem1[4][15] ), .QN(n27609) );
  SDFFX1 \mem1_reg[4][14]  ( .D(n14546), .SI(\mem1[4][13] ), .SE(test_se), 
        .CLK(n1577), .Q(\mem1[4][14] ), .QN(n27610) );
  SDFFX1 \mem1_reg[4][13]  ( .D(n14545), .SI(\mem1[4][12] ), .SE(test_se), 
        .CLK(n1578), .Q(\mem1[4][13] ), .QN(n27611) );
  SDFFX1 \mem1_reg[4][12]  ( .D(n14544), .SI(\mem1[4][11] ), .SE(test_se), 
        .CLK(n1578), .Q(\mem1[4][12] ), .QN(n27612) );
  SDFFX1 \mem1_reg[4][11]  ( .D(n14543), .SI(\mem1[4][10] ), .SE(test_se), 
        .CLK(n1578), .Q(\mem1[4][11] ), .QN(n27613) );
  SDFFX1 \mem1_reg[4][10]  ( .D(n14542), .SI(\mem1[4][9] ), .SE(test_se), 
        .CLK(n1578), .Q(\mem1[4][10] ), .QN(n27614) );
  SDFFX1 \mem1_reg[4][9]  ( .D(n14541), .SI(\mem1[4][8] ), .SE(test_se), .CLK(
        n1578), .Q(\mem1[4][9] ), .QN(n27615) );
  SDFFX1 \mem1_reg[4][8]  ( .D(n14540), .SI(\mem1[3][15] ), .SE(test_se), 
        .CLK(n1578), .Q(\mem1[4][8] ), .QN(n27616) );
  SDFFX1 \mem1_reg[3][15]  ( .D(n14539), .SI(\mem1[3][14] ), .SE(test_se), 
        .CLK(n1578), .Q(\mem1[3][15] ), .QN(n27617) );
  SDFFX1 \mem1_reg[3][14]  ( .D(n14538), .SI(\mem1[3][13] ), .SE(test_se), 
        .CLK(n1578), .Q(\mem1[3][14] ), .QN(n27618) );
  SDFFX1 \mem1_reg[3][13]  ( .D(n14537), .SI(\mem1[3][12] ), .SE(test_se), 
        .CLK(n1578), .Q(\mem1[3][13] ), .QN(n27619) );
  SDFFX1 \mem1_reg[3][12]  ( .D(n14536), .SI(\mem1[3][11] ), .SE(test_se), 
        .CLK(n1578), .Q(\mem1[3][12] ), .QN(n27620) );
  SDFFX1 \mem1_reg[3][11]  ( .D(n14535), .SI(\mem1[3][10] ), .SE(test_se), 
        .CLK(n1578), .Q(\mem1[3][11] ), .QN(n27621) );
  SDFFX1 \mem1_reg[3][10]  ( .D(n14534), .SI(\mem1[3][9] ), .SE(test_se), 
        .CLK(n1578), .Q(\mem1[3][10] ), .QN(n27622) );
  SDFFX1 \mem1_reg[3][9]  ( .D(n14533), .SI(\mem1[3][8] ), .SE(test_se), .CLK(
        n1579), .Q(\mem1[3][9] ), .QN(n27623) );
  SDFFX1 \mem1_reg[3][8]  ( .D(n14532), .SI(\mem1[2][15] ), .SE(test_se), 
        .CLK(n1579), .Q(\mem1[3][8] ), .QN(n27624) );
  SDFFX1 \mem1_reg[2][15]  ( .D(n14531), .SI(\mem1[2][14] ), .SE(test_se), 
        .CLK(n1579), .Q(\mem1[2][15] ), .QN(n27625) );
  SDFFX1 \mem1_reg[2][14]  ( .D(n14530), .SI(\mem1[2][13] ), .SE(test_se), 
        .CLK(n1579), .Q(\mem1[2][14] ), .QN(n27626) );
  SDFFX1 \mem1_reg[2][13]  ( .D(n14529), .SI(\mem1[2][12] ), .SE(test_se), 
        .CLK(n1579), .Q(\mem1[2][13] ), .QN(n27627) );
  SDFFX1 \mem1_reg[2][12]  ( .D(n14528), .SI(\mem1[2][11] ), .SE(test_se), 
        .CLK(n1579), .Q(\mem1[2][12] ), .QN(n27628) );
  SDFFX1 \mem1_reg[2][11]  ( .D(n14527), .SI(\mem1[2][10] ), .SE(test_se), 
        .CLK(n1579), .Q(\mem1[2][11] ), .QN(n27629) );
  SDFFX1 \mem1_reg[2][10]  ( .D(n14526), .SI(\mem1[2][9] ), .SE(test_se), 
        .CLK(n1579), .Q(\mem1[2][10] ), .QN(n27630) );
  SDFFX1 \mem1_reg[2][9]  ( .D(n14525), .SI(\mem1[2][8] ), .SE(test_se), .CLK(
        n1579), .Q(\mem1[2][9] ), .QN(n27631) );
  SDFFX1 \mem1_reg[2][8]  ( .D(n14524), .SI(\mem1[1][15] ), .SE(test_se), 
        .CLK(n1579), .Q(\mem1[2][8] ), .QN(n27632) );
  SDFFX1 \mem1_reg[1][15]  ( .D(n14523), .SI(\mem1[1][14] ), .SE(test_se), 
        .CLK(n1579), .Q(\mem1[1][15] ), .QN(n27633) );
  SDFFX1 \mem1_reg[1][14]  ( .D(n14522), .SI(\mem1[1][13] ), .SE(test_se), 
        .CLK(n1579), .Q(\mem1[1][14] ), .QN(n27634) );
  SDFFX1 \mem1_reg[1][13]  ( .D(n14521), .SI(\mem1[1][12] ), .SE(test_se), 
        .CLK(n1580), .Q(\mem1[1][13] ), .QN(n27635) );
  SDFFX1 \mem1_reg[1][12]  ( .D(n14520), .SI(\mem1[1][11] ), .SE(test_se), 
        .CLK(n1580), .Q(\mem1[1][12] ), .QN(n27636) );
  SDFFX1 \mem1_reg[1][11]  ( .D(n14519), .SI(\mem1[1][10] ), .SE(test_se), 
        .CLK(n1580), .Q(\mem1[1][11] ), .QN(n27637) );
  SDFFX1 \mem1_reg[1][10]  ( .D(n14518), .SI(\mem1[1][9] ), .SE(test_se), 
        .CLK(n1580), .Q(\mem1[1][10] ), .QN(n27638) );
  SDFFX1 \mem1_reg[1][9]  ( .D(n14517), .SI(\mem1[1][8] ), .SE(test_se), .CLK(
        n1580), .Q(\mem1[1][9] ), .QN(n27639) );
  SDFFX1 \mem1_reg[1][8]  ( .D(n14516), .SI(\mem1[0][15] ), .SE(test_se), 
        .CLK(n1580), .Q(\mem1[1][8] ), .QN(n27640) );
  SDFFX1 \mem1_reg[0][15]  ( .D(n14515), .SI(\mem1[0][14] ), .SE(test_se), 
        .CLK(n1580), .Q(\mem1[0][15] ), .QN(n27641) );
  SDFFX1 \mem1_reg[0][14]  ( .D(n14514), .SI(\mem1[0][13] ), .SE(test_se), 
        .CLK(n1580), .Q(\mem1[0][14] ), .QN(n27642) );
  SDFFX1 \mem1_reg[0][13]  ( .D(n14513), .SI(\mem1[0][12] ), .SE(test_se), 
        .CLK(n1580), .Q(\mem1[0][13] ), .QN(n27643) );
  SDFFX1 \mem1_reg[0][12]  ( .D(n14512), .SI(\mem1[0][11] ), .SE(test_se), 
        .CLK(n1580), .Q(\mem1[0][12] ), .QN(n27644) );
  SDFFX1 \mem1_reg[0][11]  ( .D(n14511), .SI(\mem1[0][10] ), .SE(test_se), 
        .CLK(n1580), .Q(\mem1[0][11] ), .QN(n27645) );
  SDFFX1 \mem1_reg[0][10]  ( .D(n14510), .SI(\mem1[0][9] ), .SE(test_se), 
        .CLK(n1580), .Q(\mem1[0][10] ), .QN(n27646) );
  SDFFX1 \mem1_reg[0][9]  ( .D(n14509), .SI(\mem1[0][8] ), .SE(test_se), .CLK(
        n1581), .Q(\mem1[0][9] ), .QN(n27647) );
  SDFFX1 \mem1_reg[0][8]  ( .D(n14508), .SI(\mem0[255][7] ), .SE(test_se), 
        .CLK(n1581), .Q(\mem1[0][8] ), .QN(n27648) );
  SDFFX1 \mem3_reg[255][31]  ( .D(n14507), .SI(\mem3[255][30] ), .SE(test_se), 
        .CLK(n2076), .Q(\mem3[255][31] ), .QN(n27649) );
  SDFFX1 \mem3_reg[255][30]  ( .D(n14506), .SI(\mem3[255][29] ), .SE(test_se), 
        .CLK(n1737), .Q(\mem3[255][30] ), .QN(n27650) );
  SDFFX1 \mem3_reg[255][29]  ( .D(n14505), .SI(\mem3[255][28] ), .SE(test_se), 
        .CLK(n1737), .Q(\mem3[255][29] ), .QN(n27651) );
  SDFFX1 \mem3_reg[255][28]  ( .D(n14504), .SI(\mem3[255][27] ), .SE(test_se), 
        .CLK(n1738), .Q(\mem3[255][28] ), .QN(n27652) );
  SDFFX1 \mem3_reg[255][27]  ( .D(n14503), .SI(\mem3[255][26] ), .SE(test_se), 
        .CLK(n1738), .Q(\mem3[255][27] ), .QN(n27653) );
  SDFFX1 \mem3_reg[255][26]  ( .D(n14502), .SI(\mem3[255][25] ), .SE(test_se), 
        .CLK(n1738), .Q(\mem3[255][26] ), .QN(n27654) );
  SDFFX1 \mem3_reg[255][25]  ( .D(n14501), .SI(\mem3[255][24] ), .SE(test_se), 
        .CLK(n1738), .Q(\mem3[255][25] ), .QN(n27655) );
  SDFFX1 \mem3_reg[255][24]  ( .D(n14500), .SI(\mem3[254][31] ), .SE(test_se), 
        .CLK(n1738), .Q(\mem3[255][24] ), .QN(n27656) );
  SDFFX1 \mem3_reg[254][31]  ( .D(n14499), .SI(\mem3[254][30] ), .SE(test_se), 
        .CLK(n1738), .Q(\mem3[254][31] ), .QN(n27657) );
  SDFFX1 \mem3_reg[254][30]  ( .D(n14498), .SI(\mem3[254][29] ), .SE(test_se), 
        .CLK(n1738), .Q(\mem3[254][30] ), .QN(n27658) );
  SDFFX1 \mem3_reg[254][29]  ( .D(n14497), .SI(\mem3[254][28] ), .SE(test_se), 
        .CLK(n1738), .Q(\mem3[254][29] ), .QN(n27659) );
  SDFFX1 \mem3_reg[254][28]  ( .D(n14496), .SI(\mem3[254][27] ), .SE(test_se), 
        .CLK(n1738), .Q(\mem3[254][28] ), .QN(n27660) );
  SDFFX1 \mem3_reg[254][27]  ( .D(n14495), .SI(\mem3[254][26] ), .SE(test_se), 
        .CLK(n1738), .Q(\mem3[254][27] ), .QN(n27661) );
  SDFFX1 \mem3_reg[254][26]  ( .D(n14494), .SI(\mem3[254][25] ), .SE(test_se), 
        .CLK(n1738), .Q(\mem3[254][26] ), .QN(n27662) );
  SDFFX1 \mem3_reg[254][25]  ( .D(n14493), .SI(\mem3[254][24] ), .SE(test_se), 
        .CLK(n1738), .Q(\mem3[254][25] ), .QN(n27663) );
  SDFFX1 \mem3_reg[254][24]  ( .D(n14492), .SI(\mem3[253][31] ), .SE(test_se), 
        .CLK(n1739), .Q(\mem3[254][24] ), .QN(n27664) );
  SDFFX1 \mem3_reg[253][31]  ( .D(n14491), .SI(\mem3[253][30] ), .SE(test_se), 
        .CLK(n1739), .Q(\mem3[253][31] ), .QN(n27665) );
  SDFFX1 \mem3_reg[253][30]  ( .D(n14490), .SI(\mem3[253][29] ), .SE(test_se), 
        .CLK(n1739), .Q(\mem3[253][30] ), .QN(n27666) );
  SDFFX1 \mem3_reg[253][29]  ( .D(n14489), .SI(\mem3[253][28] ), .SE(test_se), 
        .CLK(n1739), .Q(\mem3[253][29] ), .QN(n27667) );
  SDFFX1 \mem3_reg[253][28]  ( .D(n14488), .SI(\mem3[253][27] ), .SE(test_se), 
        .CLK(n1739), .Q(\mem3[253][28] ), .QN(n27668) );
  SDFFX1 \mem3_reg[253][27]  ( .D(n14487), .SI(\mem3[253][26] ), .SE(test_se), 
        .CLK(n1739), .Q(\mem3[253][27] ), .QN(n27669) );
  SDFFX1 \mem3_reg[253][26]  ( .D(n14486), .SI(\mem3[253][25] ), .SE(test_se), 
        .CLK(n1739), .Q(\mem3[253][26] ), .QN(n27670) );
  SDFFX1 \mem3_reg[253][25]  ( .D(n14485), .SI(\mem3[253][24] ), .SE(test_se), 
        .CLK(n1739), .Q(\mem3[253][25] ), .QN(n27671) );
  SDFFX1 \mem3_reg[253][24]  ( .D(n14484), .SI(\mem3[252][31] ), .SE(test_se), 
        .CLK(n1739), .Q(\mem3[253][24] ), .QN(n27672) );
  SDFFX1 \mem3_reg[252][31]  ( .D(n14483), .SI(\mem3[252][30] ), .SE(test_se), 
        .CLK(n1739), .Q(\mem3[252][31] ), .QN(n27673) );
  SDFFX1 \mem3_reg[252][30]  ( .D(n14482), .SI(\mem3[252][29] ), .SE(test_se), 
        .CLK(n1739), .Q(\mem3[252][30] ), .QN(n27674) );
  SDFFX1 \mem3_reg[252][29]  ( .D(n14481), .SI(\mem3[252][28] ), .SE(test_se), 
        .CLK(n1739), .Q(\mem3[252][29] ), .QN(n27675) );
  SDFFX1 \mem3_reg[252][28]  ( .D(n14480), .SI(\mem3[252][27] ), .SE(test_se), 
        .CLK(n1740), .Q(\mem3[252][28] ), .QN(n27676) );
  SDFFX1 \mem3_reg[252][27]  ( .D(n14479), .SI(\mem3[252][26] ), .SE(test_se), 
        .CLK(n1740), .Q(\mem3[252][27] ), .QN(n27677) );
  SDFFX1 \mem3_reg[252][26]  ( .D(n14478), .SI(\mem3[252][25] ), .SE(test_se), 
        .CLK(n1740), .Q(\mem3[252][26] ), .QN(n27678) );
  SDFFX1 \mem3_reg[252][25]  ( .D(n14477), .SI(\mem3[252][24] ), .SE(test_se), 
        .CLK(n1740), .Q(\mem3[252][25] ), .QN(n27679) );
  SDFFX1 \mem3_reg[252][24]  ( .D(n14476), .SI(\mem3[251][31] ), .SE(test_se), 
        .CLK(n1740), .Q(\mem3[252][24] ), .QN(n27680) );
  SDFFX1 \mem3_reg[251][31]  ( .D(n14475), .SI(\mem3[251][30] ), .SE(test_se), 
        .CLK(n2045), .Q(\mem3[251][31] ), .QN(n27681) );
  SDFFX1 \mem3_reg[251][30]  ( .D(n14474), .SI(\mem3[251][29] ), .SE(test_se), 
        .CLK(n2045), .Q(\mem3[251][30] ), .QN(n27682) );
  SDFFX1 \mem3_reg[251][29]  ( .D(n14473), .SI(\mem3[251][28] ), .SE(test_se), 
        .CLK(n2045), .Q(\mem3[251][29] ), .QN(n27683) );
  SDFFX1 \mem3_reg[251][28]  ( .D(n14472), .SI(\mem3[251][27] ), .SE(test_se), 
        .CLK(n2045), .Q(\mem3[251][28] ), .QN(n27684) );
  SDFFX1 \mem3_reg[251][27]  ( .D(n14471), .SI(\mem3[251][26] ), .SE(test_se), 
        .CLK(n2045), .Q(\mem3[251][27] ), .QN(n27685) );
  SDFFX1 \mem3_reg[251][26]  ( .D(n14470), .SI(\mem3[251][25] ), .SE(test_se), 
        .CLK(n2045), .Q(\mem3[251][26] ), .QN(n27686) );
  SDFFX1 \mem3_reg[251][25]  ( .D(n14469), .SI(\mem3[251][24] ), .SE(test_se), 
        .CLK(n2045), .Q(\mem3[251][25] ), .QN(n27687) );
  SDFFX1 \mem3_reg[251][24]  ( .D(n14468), .SI(\mem3[250][31] ), .SE(test_se), 
        .CLK(n2045), .Q(\mem3[251][24] ), .QN(n27688) );
  SDFFX1 \mem3_reg[250][31]  ( .D(n14467), .SI(\mem3[250][30] ), .SE(test_se), 
        .CLK(n2045), .Q(\mem3[250][31] ), .QN(n27689) );
  SDFFX1 \mem3_reg[250][30]  ( .D(n14466), .SI(\mem3[250][29] ), .SE(test_se), 
        .CLK(n2045), .Q(\mem3[250][30] ), .QN(n27690) );
  SDFFX1 \mem3_reg[250][29]  ( .D(n14465), .SI(\mem3[250][28] ), .SE(test_se), 
        .CLK(n2046), .Q(\mem3[250][29] ), .QN(n27691) );
  SDFFX1 \mem3_reg[250][28]  ( .D(n14464), .SI(\mem3[250][27] ), .SE(test_se), 
        .CLK(n2046), .Q(\mem3[250][28] ), .QN(n27692) );
  SDFFX1 \mem3_reg[250][27]  ( .D(n14463), .SI(\mem3[250][26] ), .SE(test_se), 
        .CLK(n2046), .Q(\mem3[250][27] ), .QN(n27693) );
  SDFFX1 \mem3_reg[250][26]  ( .D(n14462), .SI(\mem3[250][25] ), .SE(test_se), 
        .CLK(n2046), .Q(\mem3[250][26] ), .QN(n27694) );
  SDFFX1 \mem3_reg[250][25]  ( .D(n14461), .SI(\mem3[250][24] ), .SE(test_se), 
        .CLK(n2046), .Q(\mem3[250][25] ), .QN(n27695) );
  SDFFX1 \mem3_reg[250][24]  ( .D(n14460), .SI(\mem3[249][31] ), .SE(test_se), 
        .CLK(n2046), .Q(\mem3[250][24] ), .QN(n27696) );
  SDFFX1 \mem3_reg[249][31]  ( .D(n14459), .SI(\mem3[249][30] ), .SE(test_se), 
        .CLK(n2046), .Q(\mem3[249][31] ), .QN(n27697) );
  SDFFX1 \mem3_reg[249][30]  ( .D(n14458), .SI(\mem3[249][29] ), .SE(test_se), 
        .CLK(n2046), .Q(\mem3[249][30] ), .QN(n27698) );
  SDFFX1 \mem3_reg[249][29]  ( .D(n14457), .SI(\mem3[249][28] ), .SE(test_se), 
        .CLK(n2046), .Q(\mem3[249][29] ), .QN(n27699) );
  SDFFX1 \mem3_reg[249][28]  ( .D(n14456), .SI(\mem3[249][27] ), .SE(test_se), 
        .CLK(n2046), .Q(\mem3[249][28] ), .QN(n27700) );
  SDFFX1 \mem3_reg[249][27]  ( .D(n14455), .SI(\mem3[249][26] ), .SE(test_se), 
        .CLK(n2046), .Q(\mem3[249][27] ), .QN(n27701) );
  SDFFX1 \mem3_reg[249][26]  ( .D(n14454), .SI(\mem3[249][25] ), .SE(test_se), 
        .CLK(n2046), .Q(\mem3[249][26] ), .QN(n27702) );
  SDFFX1 \mem3_reg[249][25]  ( .D(n14453), .SI(\mem3[249][24] ), .SE(test_se), 
        .CLK(n2047), .Q(\mem3[249][25] ), .QN(n27703) );
  SDFFX1 \mem3_reg[249][24]  ( .D(n14452), .SI(\mem3[248][31] ), .SE(test_se), 
        .CLK(n2047), .Q(\mem3[249][24] ), .QN(n27704) );
  SDFFX1 \mem3_reg[248][31]  ( .D(n14451), .SI(\mem3[248][30] ), .SE(test_se), 
        .CLK(n2047), .Q(\mem3[248][31] ), .QN(n27705) );
  SDFFX1 \mem3_reg[248][30]  ( .D(n14450), .SI(\mem3[248][29] ), .SE(test_se), 
        .CLK(n2047), .Q(\mem3[248][30] ), .QN(n27706) );
  SDFFX1 \mem3_reg[248][29]  ( .D(n14449), .SI(\mem3[248][28] ), .SE(test_se), 
        .CLK(n2047), .Q(\mem3[248][29] ), .QN(n27707) );
  SDFFX1 \mem3_reg[248][28]  ( .D(n14448), .SI(\mem3[248][27] ), .SE(test_se), 
        .CLK(n2047), .Q(\mem3[248][28] ), .QN(n27708) );
  SDFFX1 \mem3_reg[248][27]  ( .D(n14447), .SI(\mem3[248][26] ), .SE(test_se), 
        .CLK(n2047), .Q(\mem3[248][27] ), .QN(n27709) );
  SDFFX1 \mem3_reg[248][26]  ( .D(n14446), .SI(\mem3[248][25] ), .SE(test_se), 
        .CLK(n2047), .Q(\mem3[248][26] ), .QN(n27710) );
  SDFFX1 \mem3_reg[248][25]  ( .D(n14445), .SI(\mem3[248][24] ), .SE(test_se), 
        .CLK(n2047), .Q(\mem3[248][25] ), .QN(n27711) );
  SDFFX1 \mem3_reg[248][24]  ( .D(n14444), .SI(\mem3[247][31] ), .SE(test_se), 
        .CLK(n2047), .Q(\mem3[248][24] ), .QN(n27712) );
  SDFFX1 \mem3_reg[247][31]  ( .D(n14443), .SI(\mem3[247][30] ), .SE(test_se), 
        .CLK(n2055), .Q(\mem3[247][31] ), .QN(n27713) );
  SDFFX1 \mem3_reg[247][30]  ( .D(n14442), .SI(\mem3[247][29] ), .SE(test_se), 
        .CLK(n2055), .Q(\mem3[247][30] ), .QN(n27714) );
  SDFFX1 \mem3_reg[247][29]  ( .D(n14441), .SI(\mem3[247][28] ), .SE(test_se), 
        .CLK(n2056), .Q(\mem3[247][29] ), .QN(n27715) );
  SDFFX1 \mem3_reg[247][28]  ( .D(n14440), .SI(\mem3[247][27] ), .SE(test_se), 
        .CLK(n2056), .Q(\mem3[247][28] ), .QN(n27716) );
  SDFFX1 \mem3_reg[247][27]  ( .D(n14439), .SI(\mem3[247][26] ), .SE(test_se), 
        .CLK(n2056), .Q(\mem3[247][27] ), .QN(n27717) );
  SDFFX1 \mem3_reg[247][26]  ( .D(n14438), .SI(\mem3[247][25] ), .SE(test_se), 
        .CLK(n2056), .Q(\mem3[247][26] ), .QN(n27718) );
  SDFFX1 \mem3_reg[247][25]  ( .D(n14437), .SI(\mem3[247][24] ), .SE(test_se), 
        .CLK(n2056), .Q(\mem3[247][25] ), .QN(n27719) );
  SDFFX1 \mem3_reg[247][24]  ( .D(n14436), .SI(\mem3[246][31] ), .SE(test_se), 
        .CLK(n2056), .Q(\mem3[247][24] ), .QN(n27720) );
  SDFFX1 \mem3_reg[246][31]  ( .D(n14435), .SI(\mem3[246][30] ), .SE(test_se), 
        .CLK(n2056), .Q(\mem3[246][31] ), .QN(n27721) );
  SDFFX1 \mem3_reg[246][30]  ( .D(n14434), .SI(\mem3[246][29] ), .SE(test_se), 
        .CLK(n2056), .Q(\mem3[246][30] ), .QN(n27722) );
  SDFFX1 \mem3_reg[246][29]  ( .D(n14433), .SI(\mem3[246][28] ), .SE(test_se), 
        .CLK(n2056), .Q(\mem3[246][29] ), .QN(n27723) );
  SDFFX1 \mem3_reg[246][28]  ( .D(n14432), .SI(\mem3[246][27] ), .SE(test_se), 
        .CLK(n2056), .Q(\mem3[246][28] ), .QN(n27724) );
  SDFFX1 \mem3_reg[246][27]  ( .D(n14431), .SI(\mem3[246][26] ), .SE(test_se), 
        .CLK(n2056), .Q(\mem3[246][27] ), .QN(n27725) );
  SDFFX1 \mem3_reg[246][26]  ( .D(n14430), .SI(\mem3[246][25] ), .SE(test_se), 
        .CLK(n2056), .Q(\mem3[246][26] ), .QN(n27726) );
  SDFFX1 \mem3_reg[246][25]  ( .D(n14429), .SI(\mem3[246][24] ), .SE(test_se), 
        .CLK(n2057), .Q(\mem3[246][25] ), .QN(n27727) );
  SDFFX1 \mem3_reg[246][24]  ( .D(n14428), .SI(\mem3[245][31] ), .SE(test_se), 
        .CLK(n2057), .Q(\mem3[246][24] ), .QN(n27728) );
  SDFFX1 \mem3_reg[245][31]  ( .D(n14427), .SI(\mem3[245][30] ), .SE(test_se), 
        .CLK(n2057), .Q(\mem3[245][31] ), .QN(n27729) );
  SDFFX1 \mem3_reg[245][30]  ( .D(n14426), .SI(\mem3[245][29] ), .SE(test_se), 
        .CLK(n2057), .Q(\mem3[245][30] ), .QN(n27730) );
  SDFFX1 \mem3_reg[245][29]  ( .D(n14425), .SI(\mem3[245][28] ), .SE(test_se), 
        .CLK(n2057), .Q(\mem3[245][29] ), .QN(n27731) );
  SDFFX1 \mem3_reg[245][28]  ( .D(n14424), .SI(\mem3[245][27] ), .SE(test_se), 
        .CLK(n2057), .Q(\mem3[245][28] ), .QN(n27732) );
  SDFFX1 \mem3_reg[245][27]  ( .D(n14423), .SI(\mem3[245][26] ), .SE(test_se), 
        .CLK(n2057), .Q(\mem3[245][27] ), .QN(n27733) );
  SDFFX1 \mem3_reg[245][26]  ( .D(n14422), .SI(\mem3[245][25] ), .SE(test_se), 
        .CLK(n2057), .Q(\mem3[245][26] ), .QN(n27734) );
  SDFFX1 \mem3_reg[245][25]  ( .D(n14421), .SI(\mem3[245][24] ), .SE(test_se), 
        .CLK(n2057), .Q(\mem3[245][25] ), .QN(n27735) );
  SDFFX1 \mem3_reg[245][24]  ( .D(n14420), .SI(\mem3[244][31] ), .SE(test_se), 
        .CLK(n2057), .Q(\mem3[245][24] ), .QN(n27736) );
  SDFFX1 \mem3_reg[244][31]  ( .D(n14419), .SI(\mem3[244][30] ), .SE(test_se), 
        .CLK(n2057), .Q(\mem3[244][31] ), .QN(n27737) );
  SDFFX1 \mem3_reg[244][30]  ( .D(n14418), .SI(\mem3[244][29] ), .SE(test_se), 
        .CLK(n2057), .Q(\mem3[244][30] ), .QN(n27738) );
  SDFFX1 \mem3_reg[244][29]  ( .D(n14417), .SI(\mem3[244][28] ), .SE(test_se), 
        .CLK(n2058), .Q(\mem3[244][29] ), .QN(n27739) );
  SDFFX1 \mem3_reg[244][28]  ( .D(n14416), .SI(\mem3[244][27] ), .SE(test_se), 
        .CLK(n2058), .Q(\mem3[244][28] ), .QN(n27740) );
  SDFFX1 \mem3_reg[244][27]  ( .D(n14415), .SI(\mem3[244][26] ), .SE(test_se), 
        .CLK(n2058), .Q(\mem3[244][27] ), .QN(n27741) );
  SDFFX1 \mem3_reg[244][26]  ( .D(n14414), .SI(\mem3[244][25] ), .SE(test_se), 
        .CLK(n2058), .Q(\mem3[244][26] ), .QN(n27742) );
  SDFFX1 \mem3_reg[244][25]  ( .D(n14413), .SI(\mem3[244][24] ), .SE(test_se), 
        .CLK(n2058), .Q(\mem3[244][25] ), .QN(n27743) );
  SDFFX1 \mem3_reg[244][24]  ( .D(n14412), .SI(\mem3[243][31] ), .SE(test_se), 
        .CLK(n2058), .Q(\mem3[244][24] ), .QN(n27744) );
  SDFFX1 \mem3_reg[243][31]  ( .D(n14411), .SI(\mem3[243][30] ), .SE(test_se), 
        .CLK(n2072), .Q(\mem3[243][31] ), .QN(n27745) );
  SDFFX1 \mem3_reg[243][30]  ( .D(n14410), .SI(\mem3[243][29] ), .SE(test_se), 
        .CLK(n2073), .Q(\mem3[243][30] ), .QN(n27746) );
  SDFFX1 \mem3_reg[243][29]  ( .D(n14409), .SI(\mem3[243][28] ), .SE(test_se), 
        .CLK(n2073), .Q(\mem3[243][29] ), .QN(n27747) );
  SDFFX1 \mem3_reg[243][28]  ( .D(n14408), .SI(\mem3[243][27] ), .SE(test_se), 
        .CLK(n2073), .Q(\mem3[243][28] ), .QN(n27748) );
  SDFFX1 \mem3_reg[243][27]  ( .D(n14407), .SI(\mem3[243][26] ), .SE(test_se), 
        .CLK(n2073), .Q(\mem3[243][27] ), .QN(n27749) );
  SDFFX1 \mem3_reg[243][26]  ( .D(n14406), .SI(\mem3[243][25] ), .SE(test_se), 
        .CLK(n2073), .Q(\mem3[243][26] ), .QN(n27750) );
  SDFFX1 \mem3_reg[243][25]  ( .D(n14405), .SI(\mem3[243][24] ), .SE(test_se), 
        .CLK(n2073), .Q(\mem3[243][25] ), .QN(n27751) );
  SDFFX1 \mem3_reg[243][24]  ( .D(n14404), .SI(\mem3[242][31] ), .SE(test_se), 
        .CLK(n2073), .Q(\mem3[243][24] ), .QN(n27752) );
  SDFFX1 \mem3_reg[242][31]  ( .D(n14403), .SI(\mem3[242][30] ), .SE(test_se), 
        .CLK(n2075), .Q(\mem3[242][31] ), .QN(n27753) );
  SDFFX1 \mem3_reg[242][30]  ( .D(n14402), .SI(\mem3[242][29] ), .SE(test_se), 
        .CLK(n2075), .Q(\mem3[242][30] ), .QN(n27754) );
  SDFFX1 \mem3_reg[242][29]  ( .D(n14401), .SI(\mem3[242][28] ), .SE(test_se), 
        .CLK(n2075), .Q(\mem3[242][29] ), .QN(n27755) );
  SDFFX1 \mem3_reg[242][28]  ( .D(n14400), .SI(test_si8), .SE(test_se), .CLK(
        n2076), .Q(\mem3[242][28] ), .QN(n27756) );
  SDFFX1 \mem3_reg[242][27]  ( .D(n14399), .SI(\mem3[242][26] ), .SE(test_se), 
        .CLK(n1740), .Q(\mem3[242][27] ), .QN(n27757) );
  SDFFX1 \mem3_reg[242][26]  ( .D(n14398), .SI(\mem3[242][25] ), .SE(test_se), 
        .CLK(n1740), .Q(\mem3[242][26] ), .QN(n27758) );
  SDFFX1 \mem3_reg[242][25]  ( .D(n14397), .SI(\mem3[242][24] ), .SE(test_se), 
        .CLK(n1740), .Q(\mem3[242][25] ), .QN(n27759) );
  SDFFX1 \mem3_reg[242][24]  ( .D(n14396), .SI(\mem3[241][31] ), .SE(test_se), 
        .CLK(n1740), .Q(\mem3[242][24] ), .QN(n27760) );
  SDFFX1 \mem3_reg[241][31]  ( .D(n14395), .SI(\mem3[241][30] ), .SE(test_se), 
        .CLK(n1740), .Q(\mem3[241][31] ), .QN(n27761) );
  SDFFX1 \mem3_reg[241][30]  ( .D(n14394), .SI(\mem3[241][29] ), .SE(test_se), 
        .CLK(n1740), .Q(\mem3[241][30] ), .QN(n27762) );
  SDFFX1 \mem3_reg[241][29]  ( .D(n14393), .SI(\mem3[241][28] ), .SE(test_se), 
        .CLK(n1740), .Q(\mem3[241][29] ), .QN(n27763) );
  SDFFX1 \mem3_reg[241][28]  ( .D(n14392), .SI(\mem3[241][27] ), .SE(test_se), 
        .CLK(n1741), .Q(\mem3[241][28] ), .QN(n27764) );
  SDFFX1 \mem3_reg[241][27]  ( .D(n14391), .SI(\mem3[241][26] ), .SE(test_se), 
        .CLK(n1741), .Q(\mem3[241][27] ), .QN(n27765) );
  SDFFX1 \mem3_reg[241][26]  ( .D(n14390), .SI(\mem3[241][25] ), .SE(test_se), 
        .CLK(n1741), .Q(\mem3[241][26] ), .QN(n27766) );
  SDFFX1 \mem3_reg[241][25]  ( .D(n14389), .SI(\mem3[241][24] ), .SE(test_se), 
        .CLK(n1741), .Q(\mem3[241][25] ), .QN(n27767) );
  SDFFX1 \mem3_reg[241][24]  ( .D(n14388), .SI(\mem3[240][31] ), .SE(test_se), 
        .CLK(n1741), .Q(\mem3[241][24] ), .QN(n27768) );
  SDFFX1 \mem3_reg[240][31]  ( .D(n14387), .SI(\mem3[240][30] ), .SE(test_se), 
        .CLK(n1741), .Q(\mem3[240][31] ), .QN(n27769) );
  SDFFX1 \mem3_reg[240][30]  ( .D(n14386), .SI(\mem3[240][29] ), .SE(test_se), 
        .CLK(n1741), .Q(\mem3[240][30] ), .QN(n27770) );
  SDFFX1 \mem3_reg[240][29]  ( .D(n14385), .SI(\mem3[240][28] ), .SE(test_se), 
        .CLK(n1741), .Q(\mem3[240][29] ), .QN(n27771) );
  SDFFX1 \mem3_reg[240][28]  ( .D(n14384), .SI(\mem3[240][27] ), .SE(test_se), 
        .CLK(n1741), .Q(\mem3[240][28] ), .QN(n27772) );
  SDFFX1 \mem3_reg[240][27]  ( .D(n14383), .SI(\mem3[240][26] ), .SE(test_se), 
        .CLK(n1741), .Q(\mem3[240][27] ), .QN(n27773) );
  SDFFX1 \mem3_reg[240][26]  ( .D(n14382), .SI(\mem3[240][25] ), .SE(test_se), 
        .CLK(n1741), .Q(\mem3[240][26] ), .QN(n27774) );
  SDFFX1 \mem3_reg[240][25]  ( .D(n14381), .SI(\mem3[240][24] ), .SE(test_se), 
        .CLK(n1741), .Q(\mem3[240][25] ), .QN(n27775) );
  SDFFX1 \mem3_reg[240][24]  ( .D(n14380), .SI(\mem3[239][31] ), .SE(test_se), 
        .CLK(n1742), .Q(\mem3[240][24] ), .QN(n27776) );
  SDFFX1 \mem3_reg[239][31]  ( .D(n14379), .SI(\mem3[239][30] ), .SE(test_se), 
        .CLK(n1742), .Q(\mem3[239][31] ), .QN(n27777) );
  SDFFX1 \mem3_reg[239][30]  ( .D(n14378), .SI(\mem3[239][29] ), .SE(test_se), 
        .CLK(n1742), .Q(\mem3[239][30] ), .QN(n27778) );
  SDFFX1 \mem3_reg[239][29]  ( .D(n14377), .SI(\mem3[239][28] ), .SE(test_se), 
        .CLK(n1742), .Q(\mem3[239][29] ), .QN(n27779) );
  SDFFX1 \mem3_reg[239][28]  ( .D(n14376), .SI(\mem3[239][27] ), .SE(test_se), 
        .CLK(n1742), .Q(\mem3[239][28] ), .QN(n27780) );
  SDFFX1 \mem3_reg[239][27]  ( .D(n14375), .SI(\mem3[239][26] ), .SE(test_se), 
        .CLK(n1742), .Q(\mem3[239][27] ), .QN(n27781) );
  SDFFX1 \mem3_reg[239][26]  ( .D(n14374), .SI(\mem3[239][25] ), .SE(test_se), 
        .CLK(n1742), .Q(\mem3[239][26] ), .QN(n27782) );
  SDFFX1 \mem3_reg[239][25]  ( .D(n14373), .SI(\mem3[239][24] ), .SE(test_se), 
        .CLK(n1742), .Q(\mem3[239][25] ), .QN(n27783) );
  SDFFX1 \mem3_reg[239][24]  ( .D(n14372), .SI(\mem3[238][31] ), .SE(test_se), 
        .CLK(n1742), .Q(\mem3[239][24] ), .QN(n27784) );
  SDFFX1 \mem3_reg[238][31]  ( .D(n14371), .SI(\mem3[238][30] ), .SE(test_se), 
        .CLK(n1742), .Q(\mem3[238][31] ), .QN(n27785) );
  SDFFX1 \mem3_reg[238][30]  ( .D(n14370), .SI(\mem3[238][29] ), .SE(test_se), 
        .CLK(n1742), .Q(\mem3[238][30] ), .QN(n27786) );
  SDFFX1 \mem3_reg[238][29]  ( .D(n14369), .SI(\mem3[238][28] ), .SE(test_se), 
        .CLK(n1742), .Q(\mem3[238][29] ), .QN(n27787) );
  SDFFX1 \mem3_reg[238][28]  ( .D(n14368), .SI(\mem3[238][27] ), .SE(test_se), 
        .CLK(n1743), .Q(\mem3[238][28] ), .QN(n27788) );
  SDFFX1 \mem3_reg[238][27]  ( .D(n14367), .SI(\mem3[238][26] ), .SE(test_se), 
        .CLK(n1743), .Q(\mem3[238][27] ), .QN(n27789) );
  SDFFX1 \mem3_reg[238][26]  ( .D(n14366), .SI(\mem3[238][25] ), .SE(test_se), 
        .CLK(n1743), .Q(\mem3[238][26] ), .QN(n27790) );
  SDFFX1 \mem3_reg[238][25]  ( .D(n14365), .SI(\mem3[238][24] ), .SE(test_se), 
        .CLK(n1743), .Q(\mem3[238][25] ), .QN(n27791) );
  SDFFX1 \mem3_reg[238][24]  ( .D(n14364), .SI(\mem3[237][31] ), .SE(test_se), 
        .CLK(n1743), .Q(\mem3[238][24] ), .QN(n27792) );
  SDFFX1 \mem3_reg[237][31]  ( .D(n14363), .SI(\mem3[237][30] ), .SE(test_se), 
        .CLK(n1743), .Q(\mem3[237][31] ), .QN(n27793) );
  SDFFX1 \mem3_reg[237][30]  ( .D(n14362), .SI(\mem3[237][29] ), .SE(test_se), 
        .CLK(n1743), .Q(\mem3[237][30] ), .QN(n27794) );
  SDFFX1 \mem3_reg[237][29]  ( .D(n14361), .SI(\mem3[237][28] ), .SE(test_se), 
        .CLK(n1743), .Q(\mem3[237][29] ), .QN(n27795) );
  SDFFX1 \mem3_reg[237][28]  ( .D(n14360), .SI(\mem3[237][27] ), .SE(test_se), 
        .CLK(n1743), .Q(\mem3[237][28] ), .QN(n27796) );
  SDFFX1 \mem3_reg[237][27]  ( .D(n14359), .SI(\mem3[237][26] ), .SE(test_se), 
        .CLK(n1743), .Q(\mem3[237][27] ), .QN(n27797) );
  SDFFX1 \mem3_reg[237][26]  ( .D(n14358), .SI(\mem3[237][25] ), .SE(test_se), 
        .CLK(n1743), .Q(\mem3[237][26] ), .QN(n27798) );
  SDFFX1 \mem3_reg[237][25]  ( .D(n14357), .SI(\mem3[237][24] ), .SE(test_se), 
        .CLK(n1743), .Q(\mem3[237][25] ), .QN(n27799) );
  SDFFX1 \mem3_reg[237][24]  ( .D(n14356), .SI(\mem3[236][31] ), .SE(test_se), 
        .CLK(n1744), .Q(\mem3[237][24] ), .QN(n27800) );
  SDFFX1 \mem3_reg[236][31]  ( .D(n14355), .SI(\mem3[236][30] ), .SE(test_se), 
        .CLK(n1744), .Q(\mem3[236][31] ), .QN(n27801) );
  SDFFX1 \mem3_reg[236][30]  ( .D(n14354), .SI(\mem3[236][29] ), .SE(test_se), 
        .CLK(n1744), .Q(\mem3[236][30] ), .QN(n27802) );
  SDFFX1 \mem3_reg[236][29]  ( .D(n14353), .SI(\mem3[236][28] ), .SE(test_se), 
        .CLK(n1744), .Q(\mem3[236][29] ), .QN(n27803) );
  SDFFX1 \mem3_reg[236][28]  ( .D(n14352), .SI(\mem3[236][27] ), .SE(test_se), 
        .CLK(n1744), .Q(\mem3[236][28] ), .QN(n27804) );
  SDFFX1 \mem3_reg[236][27]  ( .D(n14351), .SI(\mem3[236][26] ), .SE(test_se), 
        .CLK(n1744), .Q(\mem3[236][27] ), .QN(n27805) );
  SDFFX1 \mem3_reg[236][26]  ( .D(n14350), .SI(\mem3[236][25] ), .SE(test_se), 
        .CLK(n1744), .Q(\mem3[236][26] ), .QN(n27806) );
  SDFFX1 \mem3_reg[236][25]  ( .D(n14349), .SI(\mem3[236][24] ), .SE(test_se), 
        .CLK(n1744), .Q(\mem3[236][25] ), .QN(n27807) );
  SDFFX1 \mem3_reg[236][24]  ( .D(n14348), .SI(\mem3[235][31] ), .SE(test_se), 
        .CLK(n1744), .Q(\mem3[236][24] ), .QN(n27808) );
  SDFFX1 \mem3_reg[235][31]  ( .D(n14347), .SI(\mem3[235][30] ), .SE(test_se), 
        .CLK(n1744), .Q(\mem3[235][31] ), .QN(n27809) );
  SDFFX1 \mem3_reg[235][30]  ( .D(n14346), .SI(\mem3[235][29] ), .SE(test_se), 
        .CLK(n1744), .Q(\mem3[235][30] ), .QN(n27810) );
  SDFFX1 \mem3_reg[235][29]  ( .D(n14345), .SI(\mem3[235][28] ), .SE(test_se), 
        .CLK(n1744), .Q(\mem3[235][29] ), .QN(n27811) );
  SDFFX1 \mem3_reg[235][28]  ( .D(n14344), .SI(\mem3[235][27] ), .SE(test_se), 
        .CLK(n1745), .Q(\mem3[235][28] ), .QN(n27812) );
  SDFFX1 \mem3_reg[235][27]  ( .D(n14343), .SI(\mem3[235][26] ), .SE(test_se), 
        .CLK(n1745), .Q(\mem3[235][27] ), .QN(n27813) );
  SDFFX1 \mem3_reg[235][26]  ( .D(n14342), .SI(\mem3[235][25] ), .SE(test_se), 
        .CLK(n1745), .Q(\mem3[235][26] ), .QN(n27814) );
  SDFFX1 \mem3_reg[235][25]  ( .D(n14341), .SI(\mem3[235][24] ), .SE(test_se), 
        .CLK(n1745), .Q(\mem3[235][25] ), .QN(n27815) );
  SDFFX1 \mem3_reg[235][24]  ( .D(n14340), .SI(\mem3[234][31] ), .SE(test_se), 
        .CLK(n1745), .Q(\mem3[235][24] ), .QN(n27816) );
  SDFFX1 \mem3_reg[234][31]  ( .D(n14339), .SI(\mem3[234][30] ), .SE(test_se), 
        .CLK(n1745), .Q(\mem3[234][31] ), .QN(n27817) );
  SDFFX1 \mem3_reg[234][30]  ( .D(n14338), .SI(\mem3[234][29] ), .SE(test_se), 
        .CLK(n1745), .Q(\mem3[234][30] ), .QN(n27818) );
  SDFFX1 \mem3_reg[234][29]  ( .D(n14337), .SI(\mem3[234][28] ), .SE(test_se), 
        .CLK(n1745), .Q(\mem3[234][29] ), .QN(n27819) );
  SDFFX1 \mem3_reg[234][28]  ( .D(n14336), .SI(\mem3[234][27] ), .SE(test_se), 
        .CLK(n1745), .Q(\mem3[234][28] ), .QN(n27820) );
  SDFFX1 \mem3_reg[234][27]  ( .D(n14335), .SI(\mem3[234][26] ), .SE(test_se), 
        .CLK(n1745), .Q(\mem3[234][27] ), .QN(n27821) );
  SDFFX1 \mem3_reg[234][26]  ( .D(n14334), .SI(\mem3[234][25] ), .SE(test_se), 
        .CLK(n1745), .Q(\mem3[234][26] ), .QN(n27822) );
  SDFFX1 \mem3_reg[234][25]  ( .D(n14333), .SI(\mem3[234][24] ), .SE(test_se), 
        .CLK(n1745), .Q(\mem3[234][25] ), .QN(n27823) );
  SDFFX1 \mem3_reg[234][24]  ( .D(n14332), .SI(\mem3[233][31] ), .SE(test_se), 
        .CLK(n1746), .Q(\mem3[234][24] ), .QN(n27824) );
  SDFFX1 \mem3_reg[233][31]  ( .D(n14331), .SI(\mem3[233][30] ), .SE(test_se), 
        .CLK(n1746), .Q(\mem3[233][31] ), .QN(n27825) );
  SDFFX1 \mem3_reg[233][30]  ( .D(n14330), .SI(\mem3[233][29] ), .SE(test_se), 
        .CLK(n1746), .Q(\mem3[233][30] ), .QN(n27826) );
  SDFFX1 \mem3_reg[233][29]  ( .D(n14329), .SI(\mem3[233][28] ), .SE(test_se), 
        .CLK(n1746), .Q(\mem3[233][29] ), .QN(n27827) );
  SDFFX1 \mem3_reg[233][28]  ( .D(n14328), .SI(\mem3[233][27] ), .SE(test_se), 
        .CLK(n1746), .Q(\mem3[233][28] ), .QN(n27828) );
  SDFFX1 \mem3_reg[233][27]  ( .D(n14327), .SI(\mem3[233][26] ), .SE(test_se), 
        .CLK(n1746), .Q(\mem3[233][27] ), .QN(n27829) );
  SDFFX1 \mem3_reg[233][26]  ( .D(n14326), .SI(\mem3[233][25] ), .SE(test_se), 
        .CLK(n1746), .Q(\mem3[233][26] ), .QN(n27830) );
  SDFFX1 \mem3_reg[233][25]  ( .D(n14325), .SI(\mem3[233][24] ), .SE(test_se), 
        .CLK(n1746), .Q(\mem3[233][25] ), .QN(n27831) );
  SDFFX1 \mem3_reg[233][24]  ( .D(n14324), .SI(\mem3[232][31] ), .SE(test_se), 
        .CLK(n1746), .Q(\mem3[233][24] ), .QN(n27832) );
  SDFFX1 \mem3_reg[232][31]  ( .D(n14323), .SI(\mem3[232][30] ), .SE(test_se), 
        .CLK(n1746), .Q(\mem3[232][31] ), .QN(n27833) );
  SDFFX1 \mem3_reg[232][30]  ( .D(n14322), .SI(\mem3[232][29] ), .SE(test_se), 
        .CLK(n1746), .Q(\mem3[232][30] ), .QN(n27834) );
  SDFFX1 \mem3_reg[232][29]  ( .D(n14321), .SI(\mem3[232][28] ), .SE(test_se), 
        .CLK(n1746), .Q(\mem3[232][29] ), .QN(n27835) );
  SDFFX1 \mem3_reg[232][28]  ( .D(n14320), .SI(\mem3[232][27] ), .SE(test_se), 
        .CLK(n1747), .Q(\mem3[232][28] ), .QN(n27836) );
  SDFFX1 \mem3_reg[232][27]  ( .D(n14319), .SI(\mem3[232][26] ), .SE(test_se), 
        .CLK(n1747), .Q(\mem3[232][27] ), .QN(n27837) );
  SDFFX1 \mem3_reg[232][26]  ( .D(n14318), .SI(\mem3[232][25] ), .SE(test_se), 
        .CLK(n1747), .Q(\mem3[232][26] ), .QN(n27838) );
  SDFFX1 \mem3_reg[232][25]  ( .D(n14317), .SI(\mem3[232][24] ), .SE(test_se), 
        .CLK(n1747), .Q(\mem3[232][25] ), .QN(n27839) );
  SDFFX1 \mem3_reg[232][24]  ( .D(n14316), .SI(\mem3[231][31] ), .SE(test_se), 
        .CLK(n1747), .Q(\mem3[232][24] ), .QN(n27840) );
  SDFFX1 \mem3_reg[231][31]  ( .D(n14315), .SI(\mem3[231][30] ), .SE(test_se), 
        .CLK(n1747), .Q(\mem3[231][31] ), .QN(n27841) );
  SDFFX1 \mem3_reg[231][30]  ( .D(n14314), .SI(\mem3[231][29] ), .SE(test_se), 
        .CLK(n1747), .Q(\mem3[231][30] ), .QN(n27842) );
  SDFFX1 \mem3_reg[231][29]  ( .D(n14313), .SI(\mem3[231][28] ), .SE(test_se), 
        .CLK(n1747), .Q(\mem3[231][29] ), .QN(n27843) );
  SDFFX1 \mem3_reg[231][28]  ( .D(n14312), .SI(\mem3[231][27] ), .SE(test_se), 
        .CLK(n1747), .Q(\mem3[231][28] ), .QN(n27844) );
  SDFFX1 \mem3_reg[231][27]  ( .D(n14311), .SI(\mem3[231][26] ), .SE(test_se), 
        .CLK(n1747), .Q(\mem3[231][27] ), .QN(n27845) );
  SDFFX1 \mem3_reg[231][26]  ( .D(n14310), .SI(\mem3[231][25] ), .SE(test_se), 
        .CLK(n1747), .Q(\mem3[231][26] ), .QN(n27846) );
  SDFFX1 \mem3_reg[231][25]  ( .D(n14309), .SI(\mem3[231][24] ), .SE(test_se), 
        .CLK(n1747), .Q(\mem3[231][25] ), .QN(n27847) );
  SDFFX1 \mem3_reg[231][24]  ( .D(n14308), .SI(\mem3[230][31] ), .SE(test_se), 
        .CLK(n1748), .Q(\mem3[231][24] ), .QN(n27848) );
  SDFFX1 \mem3_reg[230][31]  ( .D(n14307), .SI(\mem3[230][30] ), .SE(test_se), 
        .CLK(n1748), .Q(\mem3[230][31] ), .QN(n27849) );
  SDFFX1 \mem3_reg[230][30]  ( .D(n14306), .SI(\mem3[230][29] ), .SE(test_se), 
        .CLK(n1748), .Q(\mem3[230][30] ), .QN(n27850) );
  SDFFX1 \mem3_reg[230][29]  ( .D(n14305), .SI(\mem3[230][28] ), .SE(test_se), 
        .CLK(n1748), .Q(\mem3[230][29] ), .QN(n27851) );
  SDFFX1 \mem3_reg[230][28]  ( .D(n14304), .SI(\mem3[230][27] ), .SE(test_se), 
        .CLK(n1748), .Q(\mem3[230][28] ), .QN(n27852) );
  SDFFX1 \mem3_reg[230][27]  ( .D(n14303), .SI(\mem3[230][26] ), .SE(test_se), 
        .CLK(n1748), .Q(\mem3[230][27] ), .QN(n27853) );
  SDFFX1 \mem3_reg[230][26]  ( .D(n14302), .SI(\mem3[230][25] ), .SE(test_se), 
        .CLK(n1748), .Q(\mem3[230][26] ), .QN(n27854) );
  SDFFX1 \mem3_reg[230][25]  ( .D(n14301), .SI(\mem3[230][24] ), .SE(test_se), 
        .CLK(n1748), .Q(\mem3[230][25] ), .QN(n27855) );
  SDFFX1 \mem3_reg[230][24]  ( .D(n14300), .SI(\mem3[229][31] ), .SE(test_se), 
        .CLK(n1748), .Q(\mem3[230][24] ), .QN(n27856) );
  SDFFX1 \mem3_reg[229][31]  ( .D(n14299), .SI(\mem3[229][30] ), .SE(test_se), 
        .CLK(n1748), .Q(\mem3[229][31] ), .QN(n27857) );
  SDFFX1 \mem3_reg[229][30]  ( .D(n14298), .SI(\mem3[229][29] ), .SE(test_se), 
        .CLK(n1748), .Q(\mem3[229][30] ), .QN(n27858) );
  SDFFX1 \mem3_reg[229][29]  ( .D(n14297), .SI(\mem3[229][28] ), .SE(test_se), 
        .CLK(n1748), .Q(\mem3[229][29] ), .QN(n27859) );
  SDFFX1 \mem3_reg[229][28]  ( .D(n14296), .SI(\mem3[229][27] ), .SE(test_se), 
        .CLK(n1749), .Q(\mem3[229][28] ), .QN(n27860) );
  SDFFX1 \mem3_reg[229][27]  ( .D(n14295), .SI(\mem3[229][26] ), .SE(test_se), 
        .CLK(n1749), .Q(\mem3[229][27] ), .QN(n27861) );
  SDFFX1 \mem3_reg[229][26]  ( .D(n14294), .SI(\mem3[229][25] ), .SE(test_se), 
        .CLK(n1749), .Q(\mem3[229][26] ), .QN(n27862) );
  SDFFX1 \mem3_reg[229][25]  ( .D(n14293), .SI(\mem3[229][24] ), .SE(test_se), 
        .CLK(n1749), .Q(\mem3[229][25] ), .QN(n27863) );
  SDFFX1 \mem3_reg[229][24]  ( .D(n14292), .SI(\mem3[228][31] ), .SE(test_se), 
        .CLK(n1749), .Q(\mem3[229][24] ), .QN(n27864) );
  SDFFX1 \mem3_reg[228][31]  ( .D(n14291), .SI(\mem3[228][30] ), .SE(test_se), 
        .CLK(n1749), .Q(\mem3[228][31] ), .QN(n27865) );
  SDFFX1 \mem3_reg[228][30]  ( .D(n14290), .SI(\mem3[228][29] ), .SE(test_se), 
        .CLK(n1749), .Q(\mem3[228][30] ), .QN(n27866) );
  SDFFX1 \mem3_reg[228][29]  ( .D(n14289), .SI(\mem3[228][28] ), .SE(test_se), 
        .CLK(n1749), .Q(\mem3[228][29] ), .QN(n27867) );
  SDFFX1 \mem3_reg[228][28]  ( .D(n14288), .SI(\mem3[228][27] ), .SE(test_se), 
        .CLK(n1749), .Q(\mem3[228][28] ), .QN(n27868) );
  SDFFX1 \mem3_reg[228][27]  ( .D(n14287), .SI(\mem3[228][26] ), .SE(test_se), 
        .CLK(n1749), .Q(\mem3[228][27] ), .QN(n27869) );
  SDFFX1 \mem3_reg[228][26]  ( .D(n14286), .SI(\mem3[228][25] ), .SE(test_se), 
        .CLK(n1749), .Q(\mem3[228][26] ), .QN(n27870) );
  SDFFX1 \mem3_reg[228][25]  ( .D(n14285), .SI(\mem3[228][24] ), .SE(test_se), 
        .CLK(n1749), .Q(\mem3[228][25] ), .QN(n27871) );
  SDFFX1 \mem3_reg[228][24]  ( .D(n14284), .SI(\mem3[227][31] ), .SE(test_se), 
        .CLK(n1750), .Q(\mem3[228][24] ), .QN(n27872) );
  SDFFX1 \mem3_reg[227][31]  ( .D(n14283), .SI(\mem3[227][30] ), .SE(test_se), 
        .CLK(n1750), .Q(\mem3[227][31] ), .QN(n27873) );
  SDFFX1 \mem3_reg[227][30]  ( .D(n14282), .SI(\mem3[227][29] ), .SE(test_se), 
        .CLK(n1750), .Q(\mem3[227][30] ), .QN(n27874) );
  SDFFX1 \mem3_reg[227][29]  ( .D(n14281), .SI(\mem3[227][28] ), .SE(test_se), 
        .CLK(n1750), .Q(\mem3[227][29] ), .QN(n27875) );
  SDFFX1 \mem3_reg[227][28]  ( .D(n14280), .SI(\mem3[227][27] ), .SE(test_se), 
        .CLK(n1750), .Q(\mem3[227][28] ), .QN(n27876) );
  SDFFX1 \mem3_reg[227][27]  ( .D(n14279), .SI(\mem3[227][26] ), .SE(test_se), 
        .CLK(n1750), .Q(\mem3[227][27] ), .QN(n27877) );
  SDFFX1 \mem3_reg[227][26]  ( .D(n14278), .SI(\mem3[227][25] ), .SE(test_se), 
        .CLK(n1750), .Q(\mem3[227][26] ), .QN(n27878) );
  SDFFX1 \mem3_reg[227][25]  ( .D(n14277), .SI(\mem3[227][24] ), .SE(test_se), 
        .CLK(n1750), .Q(\mem3[227][25] ), .QN(n27879) );
  SDFFX1 \mem3_reg[227][24]  ( .D(n14276), .SI(\mem3[226][31] ), .SE(test_se), 
        .CLK(n1750), .Q(\mem3[227][24] ), .QN(n27880) );
  SDFFX1 \mem3_reg[226][31]  ( .D(n14275), .SI(\mem3[226][30] ), .SE(test_se), 
        .CLK(n1750), .Q(\mem3[226][31] ), .QN(n27881) );
  SDFFX1 \mem3_reg[226][30]  ( .D(n14274), .SI(\mem3[226][29] ), .SE(test_se), 
        .CLK(n1750), .Q(\mem3[226][30] ), .QN(n27882) );
  SDFFX1 \mem3_reg[226][29]  ( .D(n14273), .SI(\mem3[226][28] ), .SE(test_se), 
        .CLK(n1750), .Q(\mem3[226][29] ), .QN(n27883) );
  SDFFX1 \mem3_reg[226][28]  ( .D(n14272), .SI(\mem3[226][27] ), .SE(test_se), 
        .CLK(n1751), .Q(\mem3[226][28] ), .QN(n27884) );
  SDFFX1 \mem3_reg[226][27]  ( .D(n14271), .SI(\mem3[226][26] ), .SE(test_se), 
        .CLK(n1751), .Q(\mem3[226][27] ), .QN(n27885) );
  SDFFX1 \mem3_reg[226][26]  ( .D(n14270), .SI(\mem3[226][25] ), .SE(test_se), 
        .CLK(n1751), .Q(\mem3[226][26] ), .QN(n27886) );
  SDFFX1 \mem3_reg[226][25]  ( .D(n14269), .SI(\mem3[226][24] ), .SE(test_se), 
        .CLK(n1751), .Q(\mem3[226][25] ), .QN(n27887) );
  SDFFX1 \mem3_reg[226][24]  ( .D(n14268), .SI(\mem3[225][31] ), .SE(test_se), 
        .CLK(n1751), .Q(\mem3[226][24] ), .QN(n27888) );
  SDFFX1 \mem3_reg[225][31]  ( .D(n14267), .SI(\mem3[225][30] ), .SE(test_se), 
        .CLK(n1751), .Q(\mem3[225][31] ), .QN(n27889) );
  SDFFX1 \mem3_reg[225][30]  ( .D(n14266), .SI(\mem3[225][29] ), .SE(test_se), 
        .CLK(n1751), .Q(\mem3[225][30] ), .QN(n27890) );
  SDFFX1 \mem3_reg[225][29]  ( .D(n14265), .SI(\mem3[225][28] ), .SE(test_se), 
        .CLK(n1751), .Q(\mem3[225][29] ), .QN(n27891) );
  SDFFX1 \mem3_reg[225][28]  ( .D(n14264), .SI(\mem3[225][27] ), .SE(test_se), 
        .CLK(n1751), .Q(\mem3[225][28] ), .QN(n27892) );
  SDFFX1 \mem3_reg[225][27]  ( .D(n14263), .SI(\mem3[225][26] ), .SE(test_se), 
        .CLK(n1751), .Q(\mem3[225][27] ), .QN(n27893) );
  SDFFX1 \mem3_reg[225][26]  ( .D(n14262), .SI(\mem3[225][25] ), .SE(test_se), 
        .CLK(n1751), .Q(\mem3[225][26] ), .QN(n27894) );
  SDFFX1 \mem3_reg[225][25]  ( .D(n14261), .SI(\mem3[225][24] ), .SE(test_se), 
        .CLK(n1751), .Q(\mem3[225][25] ), .QN(n27895) );
  SDFFX1 \mem3_reg[225][24]  ( .D(n14260), .SI(\mem3[224][31] ), .SE(test_se), 
        .CLK(n1752), .Q(\mem3[225][24] ), .QN(n27896) );
  SDFFX1 \mem3_reg[224][31]  ( .D(n14259), .SI(\mem3[224][30] ), .SE(test_se), 
        .CLK(n1752), .Q(\mem3[224][31] ), .QN(n27897) );
  SDFFX1 \mem3_reg[224][30]  ( .D(n14258), .SI(\mem3[224][29] ), .SE(test_se), 
        .CLK(n1752), .Q(\mem3[224][30] ), .QN(n27898) );
  SDFFX1 \mem3_reg[224][29]  ( .D(n14257), .SI(\mem3[224][28] ), .SE(test_se), 
        .CLK(n1752), .Q(\mem3[224][29] ), .QN(n27899) );
  SDFFX1 \mem3_reg[224][28]  ( .D(n14256), .SI(\mem3[224][27] ), .SE(test_se), 
        .CLK(n1752), .Q(\mem3[224][28] ), .QN(n27900) );
  SDFFX1 \mem3_reg[224][27]  ( .D(n14255), .SI(\mem3[224][26] ), .SE(test_se), 
        .CLK(n1752), .Q(\mem3[224][27] ), .QN(n27901) );
  SDFFX1 \mem3_reg[224][26]  ( .D(n14254), .SI(\mem3[224][25] ), .SE(test_se), 
        .CLK(n1752), .Q(\mem3[224][26] ), .QN(n27902) );
  SDFFX1 \mem3_reg[224][25]  ( .D(n14253), .SI(\mem3[224][24] ), .SE(test_se), 
        .CLK(n1752), .Q(\mem3[224][25] ), .QN(n27903) );
  SDFFX1 \mem3_reg[224][24]  ( .D(n14252), .SI(\mem3[223][31] ), .SE(test_se), 
        .CLK(n1752), .Q(\mem3[224][24] ), .QN(n27904) );
  SDFFX1 \mem3_reg[223][31]  ( .D(n14251), .SI(\mem3[223][30] ), .SE(test_se), 
        .CLK(n1752), .Q(\mem3[223][31] ), .QN(n27905) );
  SDFFX1 \mem3_reg[223][30]  ( .D(n14250), .SI(\mem3[223][29] ), .SE(test_se), 
        .CLK(n1752), .Q(\mem3[223][30] ), .QN(n27906) );
  SDFFX1 \mem3_reg[223][29]  ( .D(n14249), .SI(\mem3[223][28] ), .SE(test_se), 
        .CLK(n1752), .Q(\mem3[223][29] ), .QN(n27907) );
  SDFFX1 \mem3_reg[223][28]  ( .D(n14248), .SI(\mem3[223][27] ), .SE(test_se), 
        .CLK(n1753), .Q(\mem3[223][28] ), .QN(n27908) );
  SDFFX1 \mem3_reg[223][27]  ( .D(n14247), .SI(\mem3[223][26] ), .SE(test_se), 
        .CLK(n1753), .Q(\mem3[223][27] ), .QN(n27909) );
  SDFFX1 \mem3_reg[223][26]  ( .D(n14246), .SI(\mem3[223][25] ), .SE(test_se), 
        .CLK(n1753), .Q(\mem3[223][26] ), .QN(n27910) );
  SDFFX1 \mem3_reg[223][25]  ( .D(n14245), .SI(\mem3[223][24] ), .SE(test_se), 
        .CLK(n1753), .Q(\mem3[223][25] ), .QN(n27911) );
  SDFFX1 \mem3_reg[223][24]  ( .D(n14244), .SI(\mem3[222][31] ), .SE(test_se), 
        .CLK(n1753), .Q(\mem3[223][24] ), .QN(n27912) );
  SDFFX1 \mem3_reg[222][31]  ( .D(n14243), .SI(\mem3[222][30] ), .SE(test_se), 
        .CLK(n1753), .Q(\mem3[222][31] ), .QN(n27913) );
  SDFFX1 \mem3_reg[222][30]  ( .D(n14242), .SI(\mem3[222][29] ), .SE(test_se), 
        .CLK(n1753), .Q(\mem3[222][30] ), .QN(n27914) );
  SDFFX1 \mem3_reg[222][29]  ( .D(n14241), .SI(\mem3[222][28] ), .SE(test_se), 
        .CLK(n1753), .Q(\mem3[222][29] ), .QN(n27915) );
  SDFFX1 \mem3_reg[222][28]  ( .D(n14240), .SI(\mem3[222][27] ), .SE(test_se), 
        .CLK(n1753), .Q(\mem3[222][28] ), .QN(n27916) );
  SDFFX1 \mem3_reg[222][27]  ( .D(n14239), .SI(\mem3[222][26] ), .SE(test_se), 
        .CLK(n1753), .Q(\mem3[222][27] ), .QN(n27917) );
  SDFFX1 \mem3_reg[222][26]  ( .D(n14238), .SI(\mem3[222][25] ), .SE(test_se), 
        .CLK(n1753), .Q(\mem3[222][26] ), .QN(n27918) );
  SDFFX1 \mem3_reg[222][25]  ( .D(n14237), .SI(\mem3[222][24] ), .SE(test_se), 
        .CLK(n1753), .Q(\mem3[222][25] ), .QN(n27919) );
  SDFFX1 \mem3_reg[222][24]  ( .D(n14236), .SI(\mem3[221][31] ), .SE(test_se), 
        .CLK(n1754), .Q(\mem3[222][24] ), .QN(n27920) );
  SDFFX1 \mem3_reg[221][31]  ( .D(n14235), .SI(\mem3[221][30] ), .SE(test_se), 
        .CLK(n1754), .Q(\mem3[221][31] ), .QN(n27921) );
  SDFFX1 \mem3_reg[221][30]  ( .D(n14234), .SI(\mem3[221][29] ), .SE(test_se), 
        .CLK(n1754), .Q(\mem3[221][30] ), .QN(n27922) );
  SDFFX1 \mem3_reg[221][29]  ( .D(n14233), .SI(\mem3[221][28] ), .SE(test_se), 
        .CLK(n1754), .Q(\mem3[221][29] ), .QN(n27923) );
  SDFFX1 \mem3_reg[221][28]  ( .D(n14232), .SI(\mem3[221][27] ), .SE(test_se), 
        .CLK(n1754), .Q(\mem3[221][28] ), .QN(n27924) );
  SDFFX1 \mem3_reg[221][27]  ( .D(n14231), .SI(\mem3[221][26] ), .SE(test_se), 
        .CLK(n1754), .Q(\mem3[221][27] ), .QN(n27925) );
  SDFFX1 \mem3_reg[221][26]  ( .D(n14230), .SI(\mem3[221][25] ), .SE(test_se), 
        .CLK(n1754), .Q(\mem3[221][26] ), .QN(n27926) );
  SDFFX1 \mem3_reg[221][25]  ( .D(n14229), .SI(\mem3[221][24] ), .SE(test_se), 
        .CLK(n1754), .Q(\mem3[221][25] ), .QN(n27927) );
  SDFFX1 \mem3_reg[221][24]  ( .D(n14228), .SI(\mem3[220][31] ), .SE(test_se), 
        .CLK(n1754), .Q(\mem3[221][24] ), .QN(n27928) );
  SDFFX1 \mem3_reg[220][31]  ( .D(n14227), .SI(\mem3[220][30] ), .SE(test_se), 
        .CLK(n1754), .Q(\mem3[220][31] ), .QN(n27929) );
  SDFFX1 \mem3_reg[220][30]  ( .D(n14226), .SI(\mem3[220][29] ), .SE(test_se), 
        .CLK(n1754), .Q(\mem3[220][30] ), .QN(n27930) );
  SDFFX1 \mem3_reg[220][29]  ( .D(n14225), .SI(\mem3[220][28] ), .SE(test_se), 
        .CLK(n1754), .Q(\mem3[220][29] ), .QN(n27931) );
  SDFFX1 \mem3_reg[220][28]  ( .D(n14224), .SI(\mem3[220][27] ), .SE(test_se), 
        .CLK(n1755), .Q(\mem3[220][28] ), .QN(n27932) );
  SDFFX1 \mem3_reg[220][27]  ( .D(n14223), .SI(\mem3[220][26] ), .SE(test_se), 
        .CLK(n1755), .Q(\mem3[220][27] ), .QN(n27933) );
  SDFFX1 \mem3_reg[220][26]  ( .D(n14222), .SI(\mem3[220][25] ), .SE(test_se), 
        .CLK(n1755), .Q(\mem3[220][26] ), .QN(n27934) );
  SDFFX1 \mem3_reg[220][25]  ( .D(n14221), .SI(\mem3[220][24] ), .SE(test_se), 
        .CLK(n1755), .Q(\mem3[220][25] ), .QN(n27935) );
  SDFFX1 \mem3_reg[220][24]  ( .D(n14220), .SI(\mem3[219][31] ), .SE(test_se), 
        .CLK(n1755), .Q(\mem3[220][24] ), .QN(n27936) );
  SDFFX1 \mem3_reg[219][31]  ( .D(n14219), .SI(\mem3[219][30] ), .SE(test_se), 
        .CLK(n1755), .Q(\mem3[219][31] ), .QN(n27937) );
  SDFFX1 \mem3_reg[219][30]  ( .D(n14218), .SI(\mem3[219][29] ), .SE(test_se), 
        .CLK(n1755), .Q(\mem3[219][30] ), .QN(n27938) );
  SDFFX1 \mem3_reg[219][29]  ( .D(n14217), .SI(\mem3[219][28] ), .SE(test_se), 
        .CLK(n1755), .Q(\mem3[219][29] ), .QN(n27939) );
  SDFFX1 \mem3_reg[219][28]  ( .D(n14216), .SI(\mem3[219][27] ), .SE(test_se), 
        .CLK(n1755), .Q(\mem3[219][28] ), .QN(n27940) );
  SDFFX1 \mem3_reg[219][27]  ( .D(n14215), .SI(\mem3[219][26] ), .SE(test_se), 
        .CLK(n1755), .Q(\mem3[219][27] ), .QN(n27941) );
  SDFFX1 \mem3_reg[219][26]  ( .D(n14214), .SI(\mem3[219][25] ), .SE(test_se), 
        .CLK(n1755), .Q(\mem3[219][26] ), .QN(n27942) );
  SDFFX1 \mem3_reg[219][25]  ( .D(n14213), .SI(\mem3[219][24] ), .SE(test_se), 
        .CLK(n1755), .Q(\mem3[219][25] ), .QN(n27943) );
  SDFFX1 \mem3_reg[219][24]  ( .D(n14212), .SI(\mem3[218][31] ), .SE(test_se), 
        .CLK(n1756), .Q(\mem3[219][24] ), .QN(n27944) );
  SDFFX1 \mem3_reg[218][31]  ( .D(n14211), .SI(\mem3[218][30] ), .SE(test_se), 
        .CLK(n1756), .Q(\mem3[218][31] ), .QN(n27945) );
  SDFFX1 \mem3_reg[218][30]  ( .D(n14210), .SI(\mem3[218][29] ), .SE(test_se), 
        .CLK(n1756), .Q(\mem3[218][30] ), .QN(n27946) );
  SDFFX1 \mem3_reg[218][29]  ( .D(n14209), .SI(\mem3[218][28] ), .SE(test_se), 
        .CLK(n1756), .Q(\mem3[218][29] ), .QN(n27947) );
  SDFFX1 \mem3_reg[218][28]  ( .D(n14208), .SI(\mem3[218][27] ), .SE(test_se), 
        .CLK(n1756), .Q(\mem3[218][28] ), .QN(n27948) );
  SDFFX1 \mem3_reg[218][27]  ( .D(n14207), .SI(\mem3[218][26] ), .SE(test_se), 
        .CLK(n1756), .Q(\mem3[218][27] ), .QN(n27949) );
  SDFFX1 \mem3_reg[218][26]  ( .D(n14206), .SI(\mem3[218][25] ), .SE(test_se), 
        .CLK(n1756), .Q(\mem3[218][26] ), .QN(n27950) );
  SDFFX1 \mem3_reg[218][25]  ( .D(n14205), .SI(\mem3[218][24] ), .SE(test_se), 
        .CLK(n1756), .Q(\mem3[218][25] ), .QN(n27951) );
  SDFFX1 \mem3_reg[218][24]  ( .D(n14204), .SI(\mem3[217][31] ), .SE(test_se), 
        .CLK(n1756), .Q(\mem3[218][24] ), .QN(n27952) );
  SDFFX1 \mem3_reg[217][31]  ( .D(n14203), .SI(\mem3[217][30] ), .SE(test_se), 
        .CLK(n1756), .Q(\mem3[217][31] ), .QN(n27953) );
  SDFFX1 \mem3_reg[217][30]  ( .D(n14202), .SI(\mem3[217][29] ), .SE(test_se), 
        .CLK(n1756), .Q(\mem3[217][30] ), .QN(n27954) );
  SDFFX1 \mem3_reg[217][29]  ( .D(n14201), .SI(\mem3[217][28] ), .SE(test_se), 
        .CLK(n1756), .Q(\mem3[217][29] ), .QN(n27955) );
  SDFFX1 \mem3_reg[217][28]  ( .D(n14200), .SI(\mem3[217][27] ), .SE(test_se), 
        .CLK(n1757), .Q(\mem3[217][28] ), .QN(n27956) );
  SDFFX1 \mem3_reg[217][27]  ( .D(n14199), .SI(\mem3[217][26] ), .SE(test_se), 
        .CLK(n1757), .Q(\mem3[217][27] ), .QN(n27957) );
  SDFFX1 \mem3_reg[217][26]  ( .D(n14198), .SI(\mem3[217][25] ), .SE(test_se), 
        .CLK(n1757), .Q(\mem3[217][26] ), .QN(n27958) );
  SDFFX1 \mem3_reg[217][25]  ( .D(n14197), .SI(\mem3[217][24] ), .SE(test_se), 
        .CLK(n1757), .Q(\mem3[217][25] ), .QN(n27959) );
  SDFFX1 \mem3_reg[217][24]  ( .D(n14196), .SI(\mem3[216][31] ), .SE(test_se), 
        .CLK(n1757), .Q(\mem3[217][24] ), .QN(n27960) );
  SDFFX1 \mem3_reg[216][31]  ( .D(n14195), .SI(\mem3[216][30] ), .SE(test_se), 
        .CLK(n1757), .Q(\mem3[216][31] ), .QN(n27961) );
  SDFFX1 \mem3_reg[216][30]  ( .D(n14194), .SI(\mem3[216][29] ), .SE(test_se), 
        .CLK(n1757), .Q(\mem3[216][30] ), .QN(n27962) );
  SDFFX1 \mem3_reg[216][29]  ( .D(n14193), .SI(\mem3[216][28] ), .SE(test_se), 
        .CLK(n1757), .Q(\mem3[216][29] ), .QN(n27963) );
  SDFFX1 \mem3_reg[216][28]  ( .D(n14192), .SI(\mem3[216][27] ), .SE(test_se), 
        .CLK(n1757), .Q(\mem3[216][28] ), .QN(n27964) );
  SDFFX1 \mem3_reg[216][27]  ( .D(n14191), .SI(\mem3[216][26] ), .SE(test_se), 
        .CLK(n1757), .Q(\mem3[216][27] ), .QN(n27965) );
  SDFFX1 \mem3_reg[216][26]  ( .D(n14190), .SI(\mem3[216][25] ), .SE(test_se), 
        .CLK(n1757), .Q(\mem3[216][26] ), .QN(n27966) );
  SDFFX1 \mem3_reg[216][25]  ( .D(n14189), .SI(\mem3[216][24] ), .SE(test_se), 
        .CLK(n1757), .Q(\mem3[216][25] ), .QN(n27967) );
  SDFFX1 \mem3_reg[216][24]  ( .D(n14188), .SI(\mem3[215][31] ), .SE(test_se), 
        .CLK(n1758), .Q(\mem3[216][24] ), .QN(n27968) );
  SDFFX1 \mem3_reg[215][31]  ( .D(n14187), .SI(\mem3[215][30] ), .SE(test_se), 
        .CLK(n1758), .Q(\mem3[215][31] ), .QN(n27969) );
  SDFFX1 \mem3_reg[215][30]  ( .D(n14186), .SI(\mem3[215][29] ), .SE(test_se), 
        .CLK(n1758), .Q(\mem3[215][30] ), .QN(n27970) );
  SDFFX1 \mem3_reg[215][29]  ( .D(n14185), .SI(\mem3[215][28] ), .SE(test_se), 
        .CLK(n1758), .Q(\mem3[215][29] ), .QN(n27971) );
  SDFFX1 \mem3_reg[215][28]  ( .D(n14184), .SI(\mem3[215][27] ), .SE(test_se), 
        .CLK(n1758), .Q(\mem3[215][28] ), .QN(n27972) );
  SDFFX1 \mem3_reg[215][27]  ( .D(n14183), .SI(\mem3[215][26] ), .SE(test_se), 
        .CLK(n1758), .Q(\mem3[215][27] ), .QN(n27973) );
  SDFFX1 \mem3_reg[215][26]  ( .D(n14182), .SI(\mem3[215][25] ), .SE(test_se), 
        .CLK(n1758), .Q(\mem3[215][26] ), .QN(n27974) );
  SDFFX1 \mem3_reg[215][25]  ( .D(n14181), .SI(\mem3[215][24] ), .SE(test_se), 
        .CLK(n1758), .Q(\mem3[215][25] ), .QN(n27975) );
  SDFFX1 \mem3_reg[215][24]  ( .D(n14180), .SI(\mem3[214][31] ), .SE(test_se), 
        .CLK(n1758), .Q(\mem3[215][24] ), .QN(n27976) );
  SDFFX1 \mem3_reg[214][31]  ( .D(n14179), .SI(\mem3[214][30] ), .SE(test_se), 
        .CLK(n1758), .Q(\mem3[214][31] ), .QN(n27977) );
  SDFFX1 \mem3_reg[214][30]  ( .D(n14178), .SI(\mem3[214][29] ), .SE(test_se), 
        .CLK(n1758), .Q(\mem3[214][30] ), .QN(n27978) );
  SDFFX1 \mem3_reg[214][29]  ( .D(n14177), .SI(\mem3[214][28] ), .SE(test_se), 
        .CLK(n1758), .Q(\mem3[214][29] ), .QN(n27979) );
  SDFFX1 \mem3_reg[214][28]  ( .D(n14176), .SI(\mem3[214][27] ), .SE(test_se), 
        .CLK(n1759), .Q(\mem3[214][28] ), .QN(n27980) );
  SDFFX1 \mem3_reg[214][27]  ( .D(n14175), .SI(\mem3[214][26] ), .SE(test_se), 
        .CLK(n1759), .Q(\mem3[214][27] ), .QN(n27981) );
  SDFFX1 \mem3_reg[214][26]  ( .D(n14174), .SI(\mem3[214][25] ), .SE(test_se), 
        .CLK(n1759), .Q(\mem3[214][26] ), .QN(n27982) );
  SDFFX1 \mem3_reg[214][25]  ( .D(n14173), .SI(\mem3[214][24] ), .SE(test_se), 
        .CLK(n1759), .Q(\mem3[214][25] ), .QN(n27983) );
  SDFFX1 \mem3_reg[214][24]  ( .D(n14172), .SI(\mem3[213][31] ), .SE(test_se), 
        .CLK(n1759), .Q(\mem3[214][24] ), .QN(n27984) );
  SDFFX1 \mem3_reg[213][31]  ( .D(n14171), .SI(\mem3[213][30] ), .SE(test_se), 
        .CLK(n1759), .Q(\mem3[213][31] ), .QN(n27985) );
  SDFFX1 \mem3_reg[213][30]  ( .D(n14170), .SI(\mem3[213][29] ), .SE(test_se), 
        .CLK(n1759), .Q(\mem3[213][30] ), .QN(n27986) );
  SDFFX1 \mem3_reg[213][29]  ( .D(n14169), .SI(\mem3[213][28] ), .SE(test_se), 
        .CLK(n1759), .Q(\mem3[213][29] ), .QN(n27987) );
  SDFFX1 \mem3_reg[213][28]  ( .D(n14168), .SI(\mem3[213][27] ), .SE(test_se), 
        .CLK(n1759), .Q(\mem3[213][28] ), .QN(n27988) );
  SDFFX1 \mem3_reg[213][27]  ( .D(n14167), .SI(\mem3[213][26] ), .SE(test_se), 
        .CLK(n1759), .Q(\mem3[213][27] ), .QN(n27989) );
  SDFFX1 \mem3_reg[213][26]  ( .D(n14166), .SI(\mem3[213][25] ), .SE(test_se), 
        .CLK(n1759), .Q(\mem3[213][26] ), .QN(n27990) );
  SDFFX1 \mem3_reg[213][25]  ( .D(n14165), .SI(\mem3[213][24] ), .SE(test_se), 
        .CLK(n1759), .Q(\mem3[213][25] ), .QN(n27991) );
  SDFFX1 \mem3_reg[213][24]  ( .D(n14164), .SI(\mem3[212][31] ), .SE(test_se), 
        .CLK(n1760), .Q(\mem3[213][24] ), .QN(n27992) );
  SDFFX1 \mem3_reg[212][31]  ( .D(n14163), .SI(\mem3[212][30] ), .SE(test_se), 
        .CLK(n1760), .Q(\mem3[212][31] ), .QN(n27993) );
  SDFFX1 \mem3_reg[212][30]  ( .D(n14162), .SI(\mem3[212][29] ), .SE(test_se), 
        .CLK(n1760), .Q(\mem3[212][30] ), .QN(n27994) );
  SDFFX1 \mem3_reg[212][29]  ( .D(n14161), .SI(\mem3[212][28] ), .SE(test_se), 
        .CLK(n1760), .Q(\mem3[212][29] ), .QN(n27995) );
  SDFFX1 \mem3_reg[212][28]  ( .D(n14160), .SI(\mem3[212][27] ), .SE(test_se), 
        .CLK(n1760), .Q(\mem3[212][28] ), .QN(n27996) );
  SDFFX1 \mem3_reg[212][27]  ( .D(n14159), .SI(\mem3[212][26] ), .SE(test_se), 
        .CLK(n1760), .Q(\mem3[212][27] ), .QN(n27997) );
  SDFFX1 \mem3_reg[212][26]  ( .D(n14158), .SI(\mem3[212][25] ), .SE(test_se), 
        .CLK(n1760), .Q(\mem3[212][26] ), .QN(n27998) );
  SDFFX1 \mem3_reg[212][25]  ( .D(n14157), .SI(\mem3[212][24] ), .SE(test_se), 
        .CLK(n1760), .Q(\mem3[212][25] ), .QN(n27999) );
  SDFFX1 \mem3_reg[212][24]  ( .D(n14156), .SI(\mem3[211][31] ), .SE(test_se), 
        .CLK(n1760), .Q(\mem3[212][24] ), .QN(n28000) );
  SDFFX1 \mem3_reg[211][31]  ( .D(n14155), .SI(\mem3[211][30] ), .SE(test_se), 
        .CLK(n1760), .Q(\mem3[211][31] ), .QN(n28001) );
  SDFFX1 \mem3_reg[211][30]  ( .D(n14154), .SI(\mem3[211][29] ), .SE(test_se), 
        .CLK(n1760), .Q(\mem3[211][30] ), .QN(n28002) );
  SDFFX1 \mem3_reg[211][29]  ( .D(n14153), .SI(\mem3[211][28] ), .SE(test_se), 
        .CLK(n1760), .Q(\mem3[211][29] ), .QN(n28003) );
  SDFFX1 \mem3_reg[211][28]  ( .D(n14152), .SI(\mem3[211][27] ), .SE(test_se), 
        .CLK(n1761), .Q(\mem3[211][28] ), .QN(n28004) );
  SDFFX1 \mem3_reg[211][27]  ( .D(n14151), .SI(\mem3[211][26] ), .SE(test_se), 
        .CLK(n1761), .Q(\mem3[211][27] ), .QN(n28005) );
  SDFFX1 \mem3_reg[211][26]  ( .D(n14150), .SI(\mem3[211][25] ), .SE(test_se), 
        .CLK(n1761), .Q(\mem3[211][26] ), .QN(n28006) );
  SDFFX1 \mem3_reg[211][25]  ( .D(n14149), .SI(\mem3[211][24] ), .SE(test_se), 
        .CLK(n1761), .Q(\mem3[211][25] ), .QN(n28007) );
  SDFFX1 \mem3_reg[211][24]  ( .D(n14148), .SI(\mem3[210][31] ), .SE(test_se), 
        .CLK(n1761), .Q(\mem3[211][24] ), .QN(n28008) );
  SDFFX1 \mem3_reg[210][31]  ( .D(n14147), .SI(\mem3[210][30] ), .SE(test_se), 
        .CLK(n1761), .Q(\mem3[210][31] ), .QN(n28009) );
  SDFFX1 \mem3_reg[210][30]  ( .D(n14146), .SI(\mem3[210][29] ), .SE(test_se), 
        .CLK(n1761), .Q(\mem3[210][30] ), .QN(n28010) );
  SDFFX1 \mem3_reg[210][29]  ( .D(n14145), .SI(\mem3[210][28] ), .SE(test_se), 
        .CLK(n1761), .Q(\mem3[210][29] ), .QN(n28011) );
  SDFFX1 \mem3_reg[210][28]  ( .D(n14144), .SI(\mem3[210][27] ), .SE(test_se), 
        .CLK(n1761), .Q(\mem3[210][28] ), .QN(n28012) );
  SDFFX1 \mem3_reg[210][27]  ( .D(n14143), .SI(\mem3[210][26] ), .SE(test_se), 
        .CLK(n1761), .Q(\mem3[210][27] ), .QN(n28013) );
  SDFFX1 \mem3_reg[210][26]  ( .D(n14142), .SI(\mem3[210][25] ), .SE(test_se), 
        .CLK(n1761), .Q(\mem3[210][26] ), .QN(n28014) );
  SDFFX1 \mem3_reg[210][25]  ( .D(n14141), .SI(\mem3[210][24] ), .SE(test_se), 
        .CLK(n1761), .Q(\mem3[210][25] ), .QN(n28015) );
  SDFFX1 \mem3_reg[210][24]  ( .D(n14140), .SI(\mem3[209][31] ), .SE(test_se), 
        .CLK(n1762), .Q(\mem3[210][24] ), .QN(n28016) );
  SDFFX1 \mem3_reg[209][31]  ( .D(n14139), .SI(\mem3[209][30] ), .SE(test_se), 
        .CLK(n1762), .Q(\mem3[209][31] ), .QN(n28017) );
  SDFFX1 \mem3_reg[209][30]  ( .D(n14138), .SI(\mem3[209][29] ), .SE(test_se), 
        .CLK(n1762), .Q(\mem3[209][30] ), .QN(n28018) );
  SDFFX1 \mem3_reg[209][29]  ( .D(n14137), .SI(\mem3[209][28] ), .SE(test_se), 
        .CLK(n1762), .Q(\mem3[209][29] ), .QN(n28019) );
  SDFFX1 \mem3_reg[209][28]  ( .D(n14136), .SI(\mem3[209][27] ), .SE(test_se), 
        .CLK(n1762), .Q(\mem3[209][28] ), .QN(n28020) );
  SDFFX1 \mem3_reg[209][27]  ( .D(n14135), .SI(\mem3[209][26] ), .SE(test_se), 
        .CLK(n1762), .Q(\mem3[209][27] ), .QN(n28021) );
  SDFFX1 \mem3_reg[209][26]  ( .D(n14134), .SI(\mem3[209][25] ), .SE(test_se), 
        .CLK(n1762), .Q(\mem3[209][26] ), .QN(n28022) );
  SDFFX1 \mem3_reg[209][25]  ( .D(n14133), .SI(\mem3[209][24] ), .SE(test_se), 
        .CLK(n1762), .Q(\mem3[209][25] ), .QN(n28023) );
  SDFFX1 \mem3_reg[209][24]  ( .D(n14132), .SI(\mem3[208][31] ), .SE(test_se), 
        .CLK(n1762), .Q(\mem3[209][24] ), .QN(n28024) );
  SDFFX1 \mem3_reg[208][31]  ( .D(n14131), .SI(\mem3[208][30] ), .SE(test_se), 
        .CLK(n1762), .Q(\mem3[208][31] ), .QN(n28025) );
  SDFFX1 \mem3_reg[208][30]  ( .D(n14130), .SI(\mem3[208][29] ), .SE(test_se), 
        .CLK(n1762), .Q(\mem3[208][30] ), .QN(n28026) );
  SDFFX1 \mem3_reg[208][29]  ( .D(n14129), .SI(\mem3[208][28] ), .SE(test_se), 
        .CLK(n1762), .Q(\mem3[208][29] ), .QN(n28027) );
  SDFFX1 \mem3_reg[208][28]  ( .D(n14128), .SI(\mem3[208][27] ), .SE(test_se), 
        .CLK(n1763), .Q(\mem3[208][28] ), .QN(n28028) );
  SDFFX1 \mem3_reg[208][27]  ( .D(n14127), .SI(\mem3[208][26] ), .SE(test_se), 
        .CLK(n1763), .Q(\mem3[208][27] ), .QN(n28029) );
  SDFFX1 \mem3_reg[208][26]  ( .D(n14126), .SI(\mem3[208][25] ), .SE(test_se), 
        .CLK(n1763), .Q(\mem3[208][26] ), .QN(n28030) );
  SDFFX1 \mem3_reg[208][25]  ( .D(n14125), .SI(\mem3[208][24] ), .SE(test_se), 
        .CLK(n1763), .Q(\mem3[208][25] ), .QN(n28031) );
  SDFFX1 \mem3_reg[208][24]  ( .D(n14124), .SI(\mem3[207][31] ), .SE(test_se), 
        .CLK(n1763), .Q(\mem3[208][24] ), .QN(n28032) );
  SDFFX1 \mem3_reg[207][31]  ( .D(n14123), .SI(\mem3[207][30] ), .SE(test_se), 
        .CLK(n1763), .Q(\mem3[207][31] ), .QN(n28033) );
  SDFFX1 \mem3_reg[207][30]  ( .D(n14122), .SI(\mem3[207][29] ), .SE(test_se), 
        .CLK(n1763), .Q(\mem3[207][30] ), .QN(n28034) );
  SDFFX1 \mem3_reg[207][29]  ( .D(n14121), .SI(\mem3[207][28] ), .SE(test_se), 
        .CLK(n1763), .Q(\mem3[207][29] ), .QN(n28035) );
  SDFFX1 \mem3_reg[207][28]  ( .D(n14120), .SI(\mem3[207][27] ), .SE(test_se), 
        .CLK(n1763), .Q(\mem3[207][28] ), .QN(n28036) );
  SDFFX1 \mem3_reg[207][27]  ( .D(n14119), .SI(\mem3[207][26] ), .SE(test_se), 
        .CLK(n1763), .Q(\mem3[207][27] ), .QN(n28037) );
  SDFFX1 \mem3_reg[207][26]  ( .D(n14118), .SI(\mem3[207][25] ), .SE(test_se), 
        .CLK(n1763), .Q(\mem3[207][26] ), .QN(n28038) );
  SDFFX1 \mem3_reg[207][25]  ( .D(n14117), .SI(\mem3[207][24] ), .SE(test_se), 
        .CLK(n1763), .Q(\mem3[207][25] ), .QN(n28039) );
  SDFFX1 \mem3_reg[207][24]  ( .D(n14116), .SI(\mem3[206][31] ), .SE(test_se), 
        .CLK(n1764), .Q(\mem3[207][24] ), .QN(n28040) );
  SDFFX1 \mem3_reg[206][31]  ( .D(n14115), .SI(\mem3[206][30] ), .SE(test_se), 
        .CLK(n1764), .Q(\mem3[206][31] ), .QN(n28041) );
  SDFFX1 \mem3_reg[206][30]  ( .D(n14114), .SI(\mem3[206][29] ), .SE(test_se), 
        .CLK(n1764), .Q(\mem3[206][30] ), .QN(n28042) );
  SDFFX1 \mem3_reg[206][29]  ( .D(n14113), .SI(\mem3[206][28] ), .SE(test_se), 
        .CLK(n1764), .Q(\mem3[206][29] ), .QN(n28043) );
  SDFFX1 \mem3_reg[206][28]  ( .D(n14112), .SI(\mem3[206][27] ), .SE(test_se), 
        .CLK(n1764), .Q(\mem3[206][28] ), .QN(n28044) );
  SDFFX1 \mem3_reg[206][27]  ( .D(n14111), .SI(\mem3[206][26] ), .SE(test_se), 
        .CLK(n1764), .Q(\mem3[206][27] ), .QN(n28045) );
  SDFFX1 \mem3_reg[206][26]  ( .D(n14110), .SI(\mem3[206][25] ), .SE(test_se), 
        .CLK(n1764), .Q(\mem3[206][26] ), .QN(n28046) );
  SDFFX1 \mem3_reg[206][25]  ( .D(n14109), .SI(\mem3[206][24] ), .SE(test_se), 
        .CLK(n1764), .Q(\mem3[206][25] ), .QN(n28047) );
  SDFFX1 \mem3_reg[206][24]  ( .D(n14108), .SI(\mem3[205][31] ), .SE(test_se), 
        .CLK(n1764), .Q(\mem3[206][24] ), .QN(n28048) );
  SDFFX1 \mem3_reg[205][31]  ( .D(n14107), .SI(\mem3[205][30] ), .SE(test_se), 
        .CLK(n1764), .Q(\mem3[205][31] ), .QN(n28049) );
  SDFFX1 \mem3_reg[205][30]  ( .D(n14106), .SI(\mem3[205][29] ), .SE(test_se), 
        .CLK(n1764), .Q(\mem3[205][30] ), .QN(n28050) );
  SDFFX1 \mem3_reg[205][29]  ( .D(n14105), .SI(\mem3[205][28] ), .SE(test_se), 
        .CLK(n1764), .Q(\mem3[205][29] ), .QN(n28051) );
  SDFFX1 \mem3_reg[205][28]  ( .D(n14104), .SI(\mem3[205][27] ), .SE(test_se), 
        .CLK(n1765), .Q(\mem3[205][28] ), .QN(n28052) );
  SDFFX1 \mem3_reg[205][27]  ( .D(n14103), .SI(\mem3[205][26] ), .SE(test_se), 
        .CLK(n1765), .Q(\mem3[205][27] ), .QN(n28053) );
  SDFFX1 \mem3_reg[205][26]  ( .D(n14102), .SI(\mem3[205][25] ), .SE(test_se), 
        .CLK(n1765), .Q(\mem3[205][26] ), .QN(n28054) );
  SDFFX1 \mem3_reg[205][25]  ( .D(n14101), .SI(\mem3[205][24] ), .SE(test_se), 
        .CLK(n1765), .Q(\mem3[205][25] ), .QN(n28055) );
  SDFFX1 \mem3_reg[205][24]  ( .D(n14100), .SI(\mem3[204][31] ), .SE(test_se), 
        .CLK(n1765), .Q(\mem3[205][24] ), .QN(n28056) );
  SDFFX1 \mem3_reg[204][31]  ( .D(n14099), .SI(\mem3[204][30] ), .SE(test_se), 
        .CLK(n1765), .Q(\mem3[204][31] ), .QN(n28057) );
  SDFFX1 \mem3_reg[204][30]  ( .D(n14098), .SI(\mem3[204][29] ), .SE(test_se), 
        .CLK(n1765), .Q(\mem3[204][30] ), .QN(n28058) );
  SDFFX1 \mem3_reg[204][29]  ( .D(n14097), .SI(\mem3[204][28] ), .SE(test_se), 
        .CLK(n1765), .Q(\mem3[204][29] ), .QN(n28059) );
  SDFFX1 \mem3_reg[204][28]  ( .D(n14096), .SI(\mem3[204][27] ), .SE(test_se), 
        .CLK(n1765), .Q(\mem3[204][28] ), .QN(n28060) );
  SDFFX1 \mem3_reg[204][27]  ( .D(n14095), .SI(\mem3[204][26] ), .SE(test_se), 
        .CLK(n1765), .Q(\mem3[204][27] ), .QN(n28061) );
  SDFFX1 \mem3_reg[204][26]  ( .D(n14094), .SI(\mem3[204][25] ), .SE(test_se), 
        .CLK(n1765), .Q(\mem3[204][26] ), .QN(n28062) );
  SDFFX1 \mem3_reg[204][25]  ( .D(n14093), .SI(\mem3[204][24] ), .SE(test_se), 
        .CLK(n1765), .Q(\mem3[204][25] ), .QN(n28063) );
  SDFFX1 \mem3_reg[204][24]  ( .D(n14092), .SI(\mem3[203][31] ), .SE(test_se), 
        .CLK(n1766), .Q(\mem3[204][24] ), .QN(n28064) );
  SDFFX1 \mem3_reg[203][31]  ( .D(n14091), .SI(\mem3[203][30] ), .SE(test_se), 
        .CLK(n1766), .Q(\mem3[203][31] ), .QN(n28065) );
  SDFFX1 \mem3_reg[203][30]  ( .D(n14090), .SI(\mem3[203][29] ), .SE(test_se), 
        .CLK(n1766), .Q(\mem3[203][30] ), .QN(n28066) );
  SDFFX1 \mem3_reg[203][29]  ( .D(n14089), .SI(\mem3[203][28] ), .SE(test_se), 
        .CLK(n1766), .Q(\mem3[203][29] ), .QN(n28067) );
  SDFFX1 \mem3_reg[203][28]  ( .D(n14088), .SI(\mem3[203][27] ), .SE(test_se), 
        .CLK(n1766), .Q(\mem3[203][28] ), .QN(n28068) );
  SDFFX1 \mem3_reg[203][27]  ( .D(n14087), .SI(\mem3[203][26] ), .SE(test_se), 
        .CLK(n1766), .Q(\mem3[203][27] ), .QN(n28069) );
  SDFFX1 \mem3_reg[203][26]  ( .D(n14086), .SI(\mem3[203][25] ), .SE(test_se), 
        .CLK(n1766), .Q(\mem3[203][26] ), .QN(n28070) );
  SDFFX1 \mem3_reg[203][25]  ( .D(n14085), .SI(\mem3[203][24] ), .SE(test_se), 
        .CLK(n1766), .Q(\mem3[203][25] ), .QN(n28071) );
  SDFFX1 \mem3_reg[203][24]  ( .D(n14084), .SI(\mem3[202][31] ), .SE(test_se), 
        .CLK(n1766), .Q(\mem3[203][24] ), .QN(n28072) );
  SDFFX1 \mem3_reg[202][31]  ( .D(n14083), .SI(\mem3[202][30] ), .SE(test_se), 
        .CLK(n1766), .Q(\mem3[202][31] ), .QN(n28073) );
  SDFFX1 \mem3_reg[202][30]  ( .D(n14082), .SI(\mem3[202][29] ), .SE(test_se), 
        .CLK(n1766), .Q(\mem3[202][30] ), .QN(n28074) );
  SDFFX1 \mem3_reg[202][29]  ( .D(n14081), .SI(\mem3[202][28] ), .SE(test_se), 
        .CLK(n1766), .Q(\mem3[202][29] ), .QN(n28075) );
  SDFFX1 \mem3_reg[202][28]  ( .D(n14080), .SI(\mem3[202][27] ), .SE(test_se), 
        .CLK(n1767), .Q(\mem3[202][28] ), .QN(n28076) );
  SDFFX1 \mem3_reg[202][27]  ( .D(n14079), .SI(\mem3[202][26] ), .SE(test_se), 
        .CLK(n1767), .Q(\mem3[202][27] ), .QN(n28077) );
  SDFFX1 \mem3_reg[202][26]  ( .D(n14078), .SI(\mem3[202][25] ), .SE(test_se), 
        .CLK(n1767), .Q(\mem3[202][26] ), .QN(n28078) );
  SDFFX1 \mem3_reg[202][25]  ( .D(n14077), .SI(\mem3[202][24] ), .SE(test_se), 
        .CLK(n1767), .Q(\mem3[202][25] ), .QN(n28079) );
  SDFFX1 \mem3_reg[202][24]  ( .D(n14076), .SI(\mem3[201][31] ), .SE(test_se), 
        .CLK(n1767), .Q(\mem3[202][24] ), .QN(n28080) );
  SDFFX1 \mem3_reg[201][31]  ( .D(n14075), .SI(\mem3[201][30] ), .SE(test_se), 
        .CLK(n1767), .Q(\mem3[201][31] ), .QN(n28081) );
  SDFFX1 \mem3_reg[201][30]  ( .D(n14074), .SI(\mem3[201][29] ), .SE(test_se), 
        .CLK(n1767), .Q(\mem3[201][30] ), .QN(n28082) );
  SDFFX1 \mem3_reg[201][29]  ( .D(n14073), .SI(\mem3[201][28] ), .SE(test_se), 
        .CLK(n1767), .Q(\mem3[201][29] ), .QN(n28083) );
  SDFFX1 \mem3_reg[201][28]  ( .D(n14072), .SI(\mem3[201][27] ), .SE(test_se), 
        .CLK(n1767), .Q(\mem3[201][28] ), .QN(n28084) );
  SDFFX1 \mem3_reg[201][27]  ( .D(n14071), .SI(\mem3[201][26] ), .SE(test_se), 
        .CLK(n1767), .Q(\mem3[201][27] ), .QN(n28085) );
  SDFFX1 \mem3_reg[201][26]  ( .D(n14070), .SI(\mem3[201][25] ), .SE(test_se), 
        .CLK(n1767), .Q(\mem3[201][26] ), .QN(n28086) );
  SDFFX1 \mem3_reg[201][25]  ( .D(n14069), .SI(\mem3[201][24] ), .SE(test_se), 
        .CLK(n1767), .Q(\mem3[201][25] ), .QN(n28087) );
  SDFFX1 \mem3_reg[201][24]  ( .D(n14068), .SI(\mem3[200][31] ), .SE(test_se), 
        .CLK(n1768), .Q(\mem3[201][24] ), .QN(n28088) );
  SDFFX1 \mem3_reg[200][31]  ( .D(n14067), .SI(\mem3[200][30] ), .SE(test_se), 
        .CLK(n1768), .Q(\mem3[200][31] ), .QN(n28089) );
  SDFFX1 \mem3_reg[200][30]  ( .D(n14066), .SI(\mem3[200][29] ), .SE(test_se), 
        .CLK(n1768), .Q(\mem3[200][30] ), .QN(n28090) );
  SDFFX1 \mem3_reg[200][29]  ( .D(n14065), .SI(\mem3[200][28] ), .SE(test_se), 
        .CLK(n1768), .Q(\mem3[200][29] ), .QN(n28091) );
  SDFFX1 \mem3_reg[200][28]  ( .D(n14064), .SI(\mem3[200][27] ), .SE(test_se), 
        .CLK(n1768), .Q(\mem3[200][28] ), .QN(n28092) );
  SDFFX1 \mem3_reg[200][27]  ( .D(n14063), .SI(\mem3[200][26] ), .SE(test_se), 
        .CLK(n1768), .Q(\mem3[200][27] ), .QN(n28093) );
  SDFFX1 \mem3_reg[200][26]  ( .D(n14062), .SI(\mem3[200][25] ), .SE(test_se), 
        .CLK(n1768), .Q(\mem3[200][26] ), .QN(n28094) );
  SDFFX1 \mem3_reg[200][25]  ( .D(n14061), .SI(\mem3[200][24] ), .SE(test_se), 
        .CLK(n1768), .Q(\mem3[200][25] ), .QN(n28095) );
  SDFFX1 \mem3_reg[200][24]  ( .D(n14060), .SI(\mem3[199][31] ), .SE(test_se), 
        .CLK(n1768), .Q(\mem3[200][24] ), .QN(n28096) );
  SDFFX1 \mem3_reg[199][31]  ( .D(n14059), .SI(\mem3[199][30] ), .SE(test_se), 
        .CLK(n1768), .Q(\mem3[199][31] ), .QN(n28097) );
  SDFFX1 \mem3_reg[199][30]  ( .D(n14058), .SI(\mem3[199][29] ), .SE(test_se), 
        .CLK(n1768), .Q(\mem3[199][30] ), .QN(n28098) );
  SDFFX1 \mem3_reg[199][29]  ( .D(n14057), .SI(\mem3[199][28] ), .SE(test_se), 
        .CLK(n1768), .Q(\mem3[199][29] ), .QN(n28099) );
  SDFFX1 \mem3_reg[199][28]  ( .D(n14056), .SI(\mem3[199][27] ), .SE(test_se), 
        .CLK(n1769), .Q(\mem3[199][28] ), .QN(n28100) );
  SDFFX1 \mem3_reg[199][27]  ( .D(n14055), .SI(\mem3[199][26] ), .SE(test_se), 
        .CLK(n1769), .Q(\mem3[199][27] ), .QN(n28101) );
  SDFFX1 \mem3_reg[199][26]  ( .D(n14054), .SI(\mem3[199][25] ), .SE(test_se), 
        .CLK(n1769), .Q(\mem3[199][26] ), .QN(n28102) );
  SDFFX1 \mem3_reg[199][25]  ( .D(n14053), .SI(\mem3[199][24] ), .SE(test_se), 
        .CLK(n1769), .Q(\mem3[199][25] ), .QN(n28103) );
  SDFFX1 \mem3_reg[199][24]  ( .D(n14052), .SI(\mem3[198][31] ), .SE(test_se), 
        .CLK(n1769), .Q(\mem3[199][24] ), .QN(n28104) );
  SDFFX1 \mem3_reg[198][31]  ( .D(n14051), .SI(\mem3[198][30] ), .SE(test_se), 
        .CLK(n1769), .Q(\mem3[198][31] ), .QN(n28105) );
  SDFFX1 \mem3_reg[198][30]  ( .D(n14050), .SI(\mem3[198][29] ), .SE(test_se), 
        .CLK(n1769), .Q(\mem3[198][30] ), .QN(n28106) );
  SDFFX1 \mem3_reg[198][29]  ( .D(n14049), .SI(\mem3[198][28] ), .SE(test_se), 
        .CLK(n1769), .Q(\mem3[198][29] ), .QN(n28107) );
  SDFFX1 \mem3_reg[198][28]  ( .D(n14048), .SI(\mem3[198][27] ), .SE(test_se), 
        .CLK(n1769), .Q(\mem3[198][28] ), .QN(n28108) );
  SDFFX1 \mem3_reg[198][27]  ( .D(n14047), .SI(\mem3[198][26] ), .SE(test_se), 
        .CLK(n1769), .Q(\mem3[198][27] ), .QN(n28109) );
  SDFFX1 \mem3_reg[198][26]  ( .D(n14046), .SI(\mem3[198][25] ), .SE(test_se), 
        .CLK(n1769), .Q(\mem3[198][26] ), .QN(n28110) );
  SDFFX1 \mem3_reg[198][25]  ( .D(n14045), .SI(\mem3[198][24] ), .SE(test_se), 
        .CLK(n1769), .Q(\mem3[198][25] ), .QN(n28111) );
  SDFFX1 \mem3_reg[198][24]  ( .D(n14044), .SI(\mem3[197][31] ), .SE(test_se), 
        .CLK(n1770), .Q(\mem3[198][24] ), .QN(n28112) );
  SDFFX1 \mem3_reg[197][31]  ( .D(n14043), .SI(\mem3[197][30] ), .SE(test_se), 
        .CLK(n1770), .Q(\mem3[197][31] ), .QN(n28113) );
  SDFFX1 \mem3_reg[197][30]  ( .D(n14042), .SI(\mem3[197][29] ), .SE(test_se), 
        .CLK(n1770), .Q(\mem3[197][30] ), .QN(n28114) );
  SDFFX1 \mem3_reg[197][29]  ( .D(n14041), .SI(\mem3[197][28] ), .SE(test_se), 
        .CLK(n1770), .Q(\mem3[197][29] ), .QN(n28115) );
  SDFFX1 \mem3_reg[197][28]  ( .D(n14040), .SI(\mem3[197][27] ), .SE(test_se), 
        .CLK(n1770), .Q(\mem3[197][28] ), .QN(n28116) );
  SDFFX1 \mem3_reg[197][27]  ( .D(n14039), .SI(\mem3[197][26] ), .SE(test_se), 
        .CLK(n1770), .Q(\mem3[197][27] ), .QN(n28117) );
  SDFFX1 \mem3_reg[197][26]  ( .D(n14038), .SI(\mem3[197][25] ), .SE(test_se), 
        .CLK(n1770), .Q(\mem3[197][26] ), .QN(n28118) );
  SDFFX1 \mem3_reg[197][25]  ( .D(n14037), .SI(\mem3[197][24] ), .SE(test_se), 
        .CLK(n1770), .Q(\mem3[197][25] ), .QN(n28119) );
  SDFFX1 \mem3_reg[197][24]  ( .D(n14036), .SI(\mem3[196][31] ), .SE(test_se), 
        .CLK(n1770), .Q(\mem3[197][24] ), .QN(n28120) );
  SDFFX1 \mem3_reg[196][31]  ( .D(n14035), .SI(\mem3[196][30] ), .SE(test_se), 
        .CLK(n1770), .Q(\mem3[196][31] ), .QN(n28121) );
  SDFFX1 \mem3_reg[196][30]  ( .D(n14034), .SI(\mem3[196][29] ), .SE(test_se), 
        .CLK(n1770), .Q(\mem3[196][30] ), .QN(n28122) );
  SDFFX1 \mem3_reg[196][29]  ( .D(n14033), .SI(\mem3[196][28] ), .SE(test_se), 
        .CLK(n1770), .Q(\mem3[196][29] ), .QN(n28123) );
  SDFFX1 \mem3_reg[196][28]  ( .D(n14032), .SI(\mem3[196][27] ), .SE(test_se), 
        .CLK(n1771), .Q(\mem3[196][28] ), .QN(n28124) );
  SDFFX1 \mem3_reg[196][27]  ( .D(n14031), .SI(\mem3[196][26] ), .SE(test_se), 
        .CLK(n1771), .Q(\mem3[196][27] ), .QN(n28125) );
  SDFFX1 \mem3_reg[196][26]  ( .D(n14030), .SI(\mem3[196][25] ), .SE(test_se), 
        .CLK(n1771), .Q(\mem3[196][26] ), .QN(n28126) );
  SDFFX1 \mem3_reg[196][25]  ( .D(n14029), .SI(\mem3[196][24] ), .SE(test_se), 
        .CLK(n1771), .Q(\mem3[196][25] ), .QN(n28127) );
  SDFFX1 \mem3_reg[196][24]  ( .D(n14028), .SI(\mem3[195][31] ), .SE(test_se), 
        .CLK(n1771), .Q(\mem3[196][24] ), .QN(n28128) );
  SDFFX1 \mem3_reg[195][31]  ( .D(n14027), .SI(\mem3[195][30] ), .SE(test_se), 
        .CLK(n1771), .Q(\mem3[195][31] ), .QN(n28129) );
  SDFFX1 \mem3_reg[195][30]  ( .D(n14026), .SI(\mem3[195][29] ), .SE(test_se), 
        .CLK(n1771), .Q(\mem3[195][30] ), .QN(n28130) );
  SDFFX1 \mem3_reg[195][29]  ( .D(n14025), .SI(\mem3[195][28] ), .SE(test_se), 
        .CLK(n1771), .Q(\mem3[195][29] ), .QN(n28131) );
  SDFFX1 \mem3_reg[195][28]  ( .D(n14024), .SI(\mem3[195][27] ), .SE(test_se), 
        .CLK(n1771), .Q(\mem3[195][28] ), .QN(n28132) );
  SDFFX1 \mem3_reg[195][27]  ( .D(n14023), .SI(\mem3[195][26] ), .SE(test_se), 
        .CLK(n1771), .Q(\mem3[195][27] ), .QN(n28133) );
  SDFFX1 \mem3_reg[195][26]  ( .D(n14022), .SI(\mem3[195][25] ), .SE(test_se), 
        .CLK(n1771), .Q(\mem3[195][26] ), .QN(n28134) );
  SDFFX1 \mem3_reg[195][25]  ( .D(n14021), .SI(\mem3[195][24] ), .SE(test_se), 
        .CLK(n1771), .Q(\mem3[195][25] ), .QN(n28135) );
  SDFFX1 \mem3_reg[195][24]  ( .D(n14020), .SI(\mem3[194][31] ), .SE(test_se), 
        .CLK(n1772), .Q(\mem3[195][24] ), .QN(n28136) );
  SDFFX1 \mem3_reg[194][31]  ( .D(n14019), .SI(\mem3[194][30] ), .SE(test_se), 
        .CLK(n1772), .Q(\mem3[194][31] ), .QN(n28137) );
  SDFFX1 \mem3_reg[194][30]  ( .D(n14018), .SI(\mem3[194][29] ), .SE(test_se), 
        .CLK(n1772), .Q(\mem3[194][30] ), .QN(n28138) );
  SDFFX1 \mem3_reg[194][29]  ( .D(n14017), .SI(\mem3[194][28] ), .SE(test_se), 
        .CLK(n1772), .Q(\mem3[194][29] ), .QN(n28139) );
  SDFFX1 \mem3_reg[194][28]  ( .D(n14016), .SI(\mem3[194][27] ), .SE(test_se), 
        .CLK(n1772), .Q(\mem3[194][28] ), .QN(n28140) );
  SDFFX1 \mem3_reg[194][27]  ( .D(n14015), .SI(\mem3[194][26] ), .SE(test_se), 
        .CLK(n1772), .Q(\mem3[194][27] ), .QN(n28141) );
  SDFFX1 \mem3_reg[194][26]  ( .D(n14014), .SI(\mem3[194][25] ), .SE(test_se), 
        .CLK(n1772), .Q(\mem3[194][26] ), .QN(n28142) );
  SDFFX1 \mem3_reg[194][25]  ( .D(n14013), .SI(\mem3[194][24] ), .SE(test_se), 
        .CLK(n1772), .Q(\mem3[194][25] ), .QN(n28143) );
  SDFFX1 \mem3_reg[194][24]  ( .D(n14012), .SI(\mem3[193][31] ), .SE(test_se), 
        .CLK(n1772), .Q(\mem3[194][24] ), .QN(n28144) );
  SDFFX1 \mem3_reg[193][31]  ( .D(n14011), .SI(\mem3[193][30] ), .SE(test_se), 
        .CLK(n1772), .Q(\mem3[193][31] ), .QN(n28145) );
  SDFFX1 \mem3_reg[193][30]  ( .D(n14010), .SI(\mem3[193][29] ), .SE(test_se), 
        .CLK(n1772), .Q(\mem3[193][30] ), .QN(n28146) );
  SDFFX1 \mem3_reg[193][29]  ( .D(n14009), .SI(\mem3[193][28] ), .SE(test_se), 
        .CLK(n1772), .Q(\mem3[193][29] ), .QN(n28147) );
  SDFFX1 \mem3_reg[193][28]  ( .D(n14008), .SI(\mem3[193][27] ), .SE(test_se), 
        .CLK(n1773), .Q(\mem3[193][28] ), .QN(n28148) );
  SDFFX1 \mem3_reg[193][27]  ( .D(n14007), .SI(\mem3[193][26] ), .SE(test_se), 
        .CLK(n1773), .Q(\mem3[193][27] ), .QN(n28149) );
  SDFFX1 \mem3_reg[193][26]  ( .D(n14006), .SI(\mem3[193][25] ), .SE(test_se), 
        .CLK(n1773), .Q(\mem3[193][26] ), .QN(n28150) );
  SDFFX1 \mem3_reg[193][25]  ( .D(n14005), .SI(\mem3[193][24] ), .SE(test_se), 
        .CLK(n1773), .Q(\mem3[193][25] ), .QN(n28151) );
  SDFFX1 \mem3_reg[193][24]  ( .D(n14004), .SI(\mem3[192][31] ), .SE(test_se), 
        .CLK(n1773), .Q(\mem3[193][24] ), .QN(n28152) );
  SDFFX1 \mem3_reg[192][31]  ( .D(n14003), .SI(\mem3[192][30] ), .SE(test_se), 
        .CLK(n1773), .Q(\mem3[192][31] ), .QN(n28153) );
  SDFFX1 \mem3_reg[192][30]  ( .D(n14002), .SI(\mem3[192][29] ), .SE(test_se), 
        .CLK(n1773), .Q(\mem3[192][30] ), .QN(n28154) );
  SDFFX1 \mem3_reg[192][29]  ( .D(n14001), .SI(\mem3[192][28] ), .SE(test_se), 
        .CLK(n1773), .Q(\mem3[192][29] ), .QN(n28155) );
  SDFFX1 \mem3_reg[192][28]  ( .D(n14000), .SI(\mem3[192][27] ), .SE(test_se), 
        .CLK(n1773), .Q(\mem3[192][28] ), .QN(n28156) );
  SDFFX1 \mem3_reg[192][27]  ( .D(n13999), .SI(\mem3[192][26] ), .SE(test_se), 
        .CLK(n1773), .Q(\mem3[192][27] ), .QN(n28157) );
  SDFFX1 \mem3_reg[192][26]  ( .D(n13998), .SI(\mem3[192][25] ), .SE(test_se), 
        .CLK(n1773), .Q(\mem3[192][26] ), .QN(n28158) );
  SDFFX1 \mem3_reg[192][25]  ( .D(n13997), .SI(\mem3[192][24] ), .SE(test_se), 
        .CLK(n1773), .Q(\mem3[192][25] ), .QN(n28159) );
  SDFFX1 \mem3_reg[192][24]  ( .D(n13996), .SI(\mem3[191][31] ), .SE(test_se), 
        .CLK(n1774), .Q(\mem3[192][24] ), .QN(n28160) );
  SDFFX1 \mem3_reg[191][31]  ( .D(n13995), .SI(\mem3[191][30] ), .SE(test_se), 
        .CLK(n1774), .Q(\mem3[191][31] ), .QN(n28161) );
  SDFFX1 \mem3_reg[191][30]  ( .D(n13994), .SI(\mem3[191][29] ), .SE(test_se), 
        .CLK(n1774), .Q(\mem3[191][30] ), .QN(n28162) );
  SDFFX1 \mem3_reg[191][29]  ( .D(n13993), .SI(\mem3[191][28] ), .SE(test_se), 
        .CLK(n1774), .Q(\mem3[191][29] ), .QN(n28163) );
  SDFFX1 \mem3_reg[191][28]  ( .D(n13992), .SI(\mem3[191][27] ), .SE(test_se), 
        .CLK(n1774), .Q(\mem3[191][28] ), .QN(n28164) );
  SDFFX1 \mem3_reg[191][27]  ( .D(n13991), .SI(\mem3[191][26] ), .SE(test_se), 
        .CLK(n1774), .Q(\mem3[191][27] ), .QN(n28165) );
  SDFFX1 \mem3_reg[191][26]  ( .D(n13990), .SI(\mem3[191][25] ), .SE(test_se), 
        .CLK(n1774), .Q(\mem3[191][26] ), .QN(n28166) );
  SDFFX1 \mem3_reg[191][25]  ( .D(n13989), .SI(\mem3[191][24] ), .SE(test_se), 
        .CLK(n1774), .Q(\mem3[191][25] ), .QN(n28167) );
  SDFFX1 \mem3_reg[191][24]  ( .D(n13988), .SI(\mem3[190][31] ), .SE(test_se), 
        .CLK(n1774), .Q(\mem3[191][24] ), .QN(n28168) );
  SDFFX1 \mem3_reg[190][31]  ( .D(n13987), .SI(\mem3[190][30] ), .SE(test_se), 
        .CLK(n1774), .Q(\mem3[190][31] ), .QN(n28169) );
  SDFFX1 \mem3_reg[190][30]  ( .D(n13986), .SI(\mem3[190][29] ), .SE(test_se), 
        .CLK(n1774), .Q(\mem3[190][30] ), .QN(n28170) );
  SDFFX1 \mem3_reg[190][29]  ( .D(n13985), .SI(\mem3[190][28] ), .SE(test_se), 
        .CLK(n1774), .Q(\mem3[190][29] ), .QN(n28171) );
  SDFFX1 \mem3_reg[190][28]  ( .D(n13984), .SI(\mem3[190][27] ), .SE(test_se), 
        .CLK(n1775), .Q(\mem3[190][28] ), .QN(n28172) );
  SDFFX1 \mem3_reg[190][27]  ( .D(n13983), .SI(\mem3[190][26] ), .SE(test_se), 
        .CLK(n1775), .Q(\mem3[190][27] ), .QN(n28173) );
  SDFFX1 \mem3_reg[190][26]  ( .D(n13982), .SI(\mem3[190][25] ), .SE(test_se), 
        .CLK(n1775), .Q(\mem3[190][26] ), .QN(n28174) );
  SDFFX1 \mem3_reg[190][25]  ( .D(n13981), .SI(\mem3[190][24] ), .SE(test_se), 
        .CLK(n1775), .Q(\mem3[190][25] ), .QN(n28175) );
  SDFFX1 \mem3_reg[190][24]  ( .D(n13980), .SI(\mem3[189][31] ), .SE(test_se), 
        .CLK(n1775), .Q(\mem3[190][24] ), .QN(n28176) );
  SDFFX1 \mem3_reg[189][31]  ( .D(n13979), .SI(\mem3[189][30] ), .SE(test_se), 
        .CLK(n1775), .Q(\mem3[189][31] ), .QN(n28177) );
  SDFFX1 \mem3_reg[189][30]  ( .D(n13978), .SI(\mem3[189][29] ), .SE(test_se), 
        .CLK(n1775), .Q(\mem3[189][30] ), .QN(n28178) );
  SDFFX1 \mem3_reg[189][29]  ( .D(n13977), .SI(\mem3[189][28] ), .SE(test_se), 
        .CLK(n1775), .Q(\mem3[189][29] ), .QN(n28179) );
  SDFFX1 \mem3_reg[189][28]  ( .D(n13976), .SI(\mem3[189][27] ), .SE(test_se), 
        .CLK(n1775), .Q(\mem3[189][28] ), .QN(n28180) );
  SDFFX1 \mem3_reg[189][27]  ( .D(n13975), .SI(\mem3[189][26] ), .SE(test_se), 
        .CLK(n1775), .Q(\mem3[189][27] ), .QN(n28181) );
  SDFFX1 \mem3_reg[189][26]  ( .D(n13974), .SI(\mem3[189][25] ), .SE(test_se), 
        .CLK(n1775), .Q(\mem3[189][26] ), .QN(n28182) );
  SDFFX1 \mem3_reg[189][25]  ( .D(n13973), .SI(\mem3[189][24] ), .SE(test_se), 
        .CLK(n1775), .Q(\mem3[189][25] ), .QN(n28183) );
  SDFFX1 \mem3_reg[189][24]  ( .D(n13972), .SI(\mem3[188][31] ), .SE(test_se), 
        .CLK(n1776), .Q(\mem3[189][24] ), .QN(n28184) );
  SDFFX1 \mem3_reg[188][31]  ( .D(n13971), .SI(\mem3[188][30] ), .SE(test_se), 
        .CLK(n1776), .Q(\mem3[188][31] ), .QN(n28185) );
  SDFFX1 \mem3_reg[188][30]  ( .D(n13970), .SI(\mem3[188][29] ), .SE(test_se), 
        .CLK(n1776), .Q(\mem3[188][30] ), .QN(n28186) );
  SDFFX1 \mem3_reg[188][29]  ( .D(n13969), .SI(\mem3[188][28] ), .SE(test_se), 
        .CLK(n1776), .Q(\mem3[188][29] ), .QN(n28187) );
  SDFFX1 \mem3_reg[188][28]  ( .D(n13968), .SI(\mem3[188][27] ), .SE(test_se), 
        .CLK(n1776), .Q(\mem3[188][28] ), .QN(n28188) );
  SDFFX1 \mem3_reg[188][27]  ( .D(n13967), .SI(\mem3[188][26] ), .SE(test_se), 
        .CLK(n1776), .Q(\mem3[188][27] ), .QN(n28189) );
  SDFFX1 \mem3_reg[188][26]  ( .D(n13966), .SI(\mem3[188][25] ), .SE(test_se), 
        .CLK(n1776), .Q(\mem3[188][26] ), .QN(n28190) );
  SDFFX1 \mem3_reg[188][25]  ( .D(n13965), .SI(\mem3[188][24] ), .SE(test_se), 
        .CLK(n1776), .Q(\mem3[188][25] ), .QN(n28191) );
  SDFFX1 \mem3_reg[188][24]  ( .D(n13964), .SI(\mem3[187][31] ), .SE(test_se), 
        .CLK(n1776), .Q(\mem3[188][24] ), .QN(n28192) );
  SDFFX1 \mem3_reg[187][31]  ( .D(n13963), .SI(\mem3[187][30] ), .SE(test_se), 
        .CLK(n1776), .Q(\mem3[187][31] ), .QN(n28193) );
  SDFFX1 \mem3_reg[187][30]  ( .D(n13962), .SI(\mem3[187][29] ), .SE(test_se), 
        .CLK(n1776), .Q(\mem3[187][30] ), .QN(n28194) );
  SDFFX1 \mem3_reg[187][29]  ( .D(n13961), .SI(\mem3[187][28] ), .SE(test_se), 
        .CLK(n1776), .Q(\mem3[187][29] ), .QN(n28195) );
  SDFFX1 \mem3_reg[187][28]  ( .D(n13960), .SI(\mem3[187][27] ), .SE(test_se), 
        .CLK(n1777), .Q(\mem3[187][28] ), .QN(n28196) );
  SDFFX1 \mem3_reg[187][27]  ( .D(n13959), .SI(\mem3[187][26] ), .SE(test_se), 
        .CLK(n1777), .Q(\mem3[187][27] ), .QN(n28197) );
  SDFFX1 \mem3_reg[187][26]  ( .D(n13958), .SI(\mem3[187][25] ), .SE(test_se), 
        .CLK(n1777), .Q(\mem3[187][26] ), .QN(n28198) );
  SDFFX1 \mem3_reg[187][25]  ( .D(n13957), .SI(\mem3[187][24] ), .SE(test_se), 
        .CLK(n1777), .Q(\mem3[187][25] ), .QN(n28199) );
  SDFFX1 \mem3_reg[187][24]  ( .D(n13956), .SI(\mem3[186][31] ), .SE(test_se), 
        .CLK(n1777), .Q(\mem3[187][24] ), .QN(n28200) );
  SDFFX1 \mem3_reg[186][31]  ( .D(n13955), .SI(\mem3[186][30] ), .SE(test_se), 
        .CLK(n1777), .Q(\mem3[186][31] ), .QN(n28201) );
  SDFFX1 \mem3_reg[186][30]  ( .D(n13954), .SI(\mem3[186][29] ), .SE(test_se), 
        .CLK(n1777), .Q(\mem3[186][30] ), .QN(n28202) );
  SDFFX1 \mem3_reg[186][29]  ( .D(n13953), .SI(\mem3[186][28] ), .SE(test_se), 
        .CLK(n1777), .Q(\mem3[186][29] ), .QN(n28203) );
  SDFFX1 \mem3_reg[186][28]  ( .D(n13952), .SI(\mem3[186][27] ), .SE(test_se), 
        .CLK(n1777), .Q(\mem3[186][28] ), .QN(n28204) );
  SDFFX1 \mem3_reg[186][27]  ( .D(n13951), .SI(\mem3[186][26] ), .SE(test_se), 
        .CLK(n1777), .Q(\mem3[186][27] ), .QN(n28205) );
  SDFFX1 \mem3_reg[186][26]  ( .D(n13950), .SI(\mem3[186][25] ), .SE(test_se), 
        .CLK(n1777), .Q(\mem3[186][26] ), .QN(n28206) );
  SDFFX1 \mem3_reg[186][25]  ( .D(n13949), .SI(\mem3[186][24] ), .SE(test_se), 
        .CLK(n1777), .Q(\mem3[186][25] ), .QN(n28207) );
  SDFFX1 \mem3_reg[186][24]  ( .D(n13948), .SI(\mem3[185][31] ), .SE(test_se), 
        .CLK(n1778), .Q(\mem3[186][24] ), .QN(n28208) );
  SDFFX1 \mem3_reg[185][31]  ( .D(n13947), .SI(\mem3[185][30] ), .SE(test_se), 
        .CLK(n1778), .Q(\mem3[185][31] ), .QN(n28209) );
  SDFFX1 \mem3_reg[185][30]  ( .D(n13946), .SI(\mem3[185][29] ), .SE(test_se), 
        .CLK(n1778), .Q(\mem3[185][30] ), .QN(n28210) );
  SDFFX1 \mem3_reg[185][29]  ( .D(n13945), .SI(\mem3[185][28] ), .SE(test_se), 
        .CLK(n1778), .Q(\mem3[185][29] ), .QN(n28211) );
  SDFFX1 \mem3_reg[185][28]  ( .D(n13944), .SI(\mem3[185][27] ), .SE(test_se), 
        .CLK(n1778), .Q(\mem3[185][28] ), .QN(n28212) );
  SDFFX1 \mem3_reg[185][27]  ( .D(n13943), .SI(\mem3[185][26] ), .SE(test_se), 
        .CLK(n1778), .Q(\mem3[185][27] ), .QN(n28213) );
  SDFFX1 \mem3_reg[185][26]  ( .D(n13942), .SI(\mem3[185][25] ), .SE(test_se), 
        .CLK(n1778), .Q(\mem3[185][26] ), .QN(n28214) );
  SDFFX1 \mem3_reg[185][25]  ( .D(n13941), .SI(\mem3[185][24] ), .SE(test_se), 
        .CLK(n1778), .Q(\mem3[185][25] ), .QN(n28215) );
  SDFFX1 \mem3_reg[185][24]  ( .D(n13940), .SI(\mem3[184][31] ), .SE(test_se), 
        .CLK(n1778), .Q(\mem3[185][24] ), .QN(n28216) );
  SDFFX1 \mem3_reg[184][31]  ( .D(n13939), .SI(\mem3[184][30] ), .SE(test_se), 
        .CLK(n1778), .Q(\mem3[184][31] ), .QN(n28217) );
  SDFFX1 \mem3_reg[184][30]  ( .D(n13938), .SI(\mem3[184][29] ), .SE(test_se), 
        .CLK(n1778), .Q(\mem3[184][30] ), .QN(n28218) );
  SDFFX1 \mem3_reg[184][29]  ( .D(n13937), .SI(\mem3[184][28] ), .SE(test_se), 
        .CLK(n1778), .Q(\mem3[184][29] ), .QN(n28219) );
  SDFFX1 \mem3_reg[184][28]  ( .D(n13936), .SI(\mem3[184][27] ), .SE(test_se), 
        .CLK(n1779), .Q(\mem3[184][28] ), .QN(n28220) );
  SDFFX1 \mem3_reg[184][27]  ( .D(n13935), .SI(\mem3[184][26] ), .SE(test_se), 
        .CLK(n1779), .Q(\mem3[184][27] ), .QN(n28221) );
  SDFFX1 \mem3_reg[184][26]  ( .D(n13934), .SI(\mem3[184][25] ), .SE(test_se), 
        .CLK(n1779), .Q(\mem3[184][26] ), .QN(n28222) );
  SDFFX1 \mem3_reg[184][25]  ( .D(n13933), .SI(\mem3[184][24] ), .SE(test_se), 
        .CLK(n1779), .Q(\mem3[184][25] ), .QN(n28223) );
  SDFFX1 \mem3_reg[184][24]  ( .D(n13932), .SI(\mem3[183][31] ), .SE(test_se), 
        .CLK(n1779), .Q(\mem3[184][24] ), .QN(n28224) );
  SDFFX1 \mem3_reg[183][31]  ( .D(n13931), .SI(\mem3[183][30] ), .SE(test_se), 
        .CLK(n1779), .Q(\mem3[183][31] ), .QN(n28225) );
  SDFFX1 \mem3_reg[183][30]  ( .D(n13930), .SI(\mem3[183][29] ), .SE(test_se), 
        .CLK(n1779), .Q(\mem3[183][30] ), .QN(n28226) );
  SDFFX1 \mem3_reg[183][29]  ( .D(n13929), .SI(\mem3[183][28] ), .SE(test_se), 
        .CLK(n1779), .Q(\mem3[183][29] ), .QN(n28227) );
  SDFFX1 \mem3_reg[183][28]  ( .D(n13928), .SI(\mem3[183][27] ), .SE(test_se), 
        .CLK(n1779), .Q(\mem3[183][28] ), .QN(n28228) );
  SDFFX1 \mem3_reg[183][27]  ( .D(n13927), .SI(\mem3[183][26] ), .SE(test_se), 
        .CLK(n1779), .Q(\mem3[183][27] ), .QN(n28229) );
  SDFFX1 \mem3_reg[183][26]  ( .D(n13926), .SI(\mem3[183][25] ), .SE(test_se), 
        .CLK(n1779), .Q(\mem3[183][26] ), .QN(n28230) );
  SDFFX1 \mem3_reg[183][25]  ( .D(n13925), .SI(\mem3[183][24] ), .SE(test_se), 
        .CLK(n1779), .Q(\mem3[183][25] ), .QN(n28231) );
  SDFFX1 \mem3_reg[183][24]  ( .D(n13924), .SI(\mem3[182][31] ), .SE(test_se), 
        .CLK(n1780), .Q(\mem3[183][24] ), .QN(n28232) );
  SDFFX1 \mem3_reg[182][31]  ( .D(n13923), .SI(\mem3[182][30] ), .SE(test_se), 
        .CLK(n1780), .Q(\mem3[182][31] ), .QN(n28233) );
  SDFFX1 \mem3_reg[182][30]  ( .D(n13922), .SI(\mem3[182][29] ), .SE(test_se), 
        .CLK(n1780), .Q(\mem3[182][30] ), .QN(n28234) );
  SDFFX1 \mem3_reg[182][29]  ( .D(n13921), .SI(\mem3[182][28] ), .SE(test_se), 
        .CLK(n1780), .Q(\mem3[182][29] ), .QN(n28235) );
  SDFFX1 \mem3_reg[182][28]  ( .D(n13920), .SI(\mem3[182][27] ), .SE(test_se), 
        .CLK(n1780), .Q(\mem3[182][28] ), .QN(n28236) );
  SDFFX1 \mem3_reg[182][27]  ( .D(n13919), .SI(\mem3[182][26] ), .SE(test_se), 
        .CLK(n1780), .Q(\mem3[182][27] ), .QN(n28237) );
  SDFFX1 \mem3_reg[182][26]  ( .D(n13918), .SI(\mem3[182][25] ), .SE(test_se), 
        .CLK(n1780), .Q(\mem3[182][26] ), .QN(n28238) );
  SDFFX1 \mem3_reg[182][25]  ( .D(n13917), .SI(\mem3[182][24] ), .SE(test_se), 
        .CLK(n1780), .Q(\mem3[182][25] ), .QN(n28239) );
  SDFFX1 \mem3_reg[182][24]  ( .D(n13916), .SI(\mem3[181][31] ), .SE(test_se), 
        .CLK(n1780), .Q(\mem3[182][24] ), .QN(n28240) );
  SDFFX1 \mem3_reg[181][31]  ( .D(n13915), .SI(\mem3[181][30] ), .SE(test_se), 
        .CLK(n1780), .Q(\mem3[181][31] ), .QN(n28241) );
  SDFFX1 \mem3_reg[181][30]  ( .D(n13914), .SI(\mem3[181][29] ), .SE(test_se), 
        .CLK(n1780), .Q(\mem3[181][30] ), .QN(n28242) );
  SDFFX1 \mem3_reg[181][29]  ( .D(n13913), .SI(\mem3[181][28] ), .SE(test_se), 
        .CLK(n1780), .Q(\mem3[181][29] ), .QN(n28243) );
  SDFFX1 \mem3_reg[181][28]  ( .D(n13912), .SI(\mem3[181][27] ), .SE(test_se), 
        .CLK(n1781), .Q(\mem3[181][28] ), .QN(n28244) );
  SDFFX1 \mem3_reg[181][27]  ( .D(n13911), .SI(\mem3[181][26] ), .SE(test_se), 
        .CLK(n1781), .Q(\mem3[181][27] ), .QN(n28245) );
  SDFFX1 \mem3_reg[181][26]  ( .D(n13910), .SI(\mem3[181][25] ), .SE(test_se), 
        .CLK(n1781), .Q(\mem3[181][26] ), .QN(n28246) );
  SDFFX1 \mem3_reg[181][25]  ( .D(n13909), .SI(\mem3[181][24] ), .SE(test_se), 
        .CLK(n1781), .Q(\mem3[181][25] ), .QN(n28247) );
  SDFFX1 \mem3_reg[181][24]  ( .D(n13908), .SI(\mem3[180][31] ), .SE(test_se), 
        .CLK(n1781), .Q(\mem3[181][24] ), .QN(n28248) );
  SDFFX1 \mem3_reg[180][31]  ( .D(n13907), .SI(\mem3[180][30] ), .SE(test_se), 
        .CLK(n1781), .Q(\mem3[180][31] ), .QN(n28249) );
  SDFFX1 \mem3_reg[180][30]  ( .D(n13906), .SI(\mem3[180][29] ), .SE(test_se), 
        .CLK(n1781), .Q(\mem3[180][30] ), .QN(n28250) );
  SDFFX1 \mem3_reg[180][29]  ( .D(n13905), .SI(\mem3[180][28] ), .SE(test_se), 
        .CLK(n1781), .Q(\mem3[180][29] ), .QN(n28251) );
  SDFFX1 \mem3_reg[180][28]  ( .D(n13904), .SI(\mem3[180][27] ), .SE(test_se), 
        .CLK(n1781), .Q(\mem3[180][28] ), .QN(n28252) );
  SDFFX1 \mem3_reg[180][27]  ( .D(n13903), .SI(\mem3[180][26] ), .SE(test_se), 
        .CLK(n1781), .Q(\mem3[180][27] ), .QN(n28253) );
  SDFFX1 \mem3_reg[180][26]  ( .D(n13902), .SI(\mem3[180][25] ), .SE(test_se), 
        .CLK(n1781), .Q(\mem3[180][26] ), .QN(n28254) );
  SDFFX1 \mem3_reg[180][25]  ( .D(n13901), .SI(\mem3[180][24] ), .SE(test_se), 
        .CLK(n1781), .Q(\mem3[180][25] ), .QN(n28255) );
  SDFFX1 \mem3_reg[180][24]  ( .D(n13900), .SI(\mem3[179][31] ), .SE(test_se), 
        .CLK(n1782), .Q(\mem3[180][24] ), .QN(n28256) );
  SDFFX1 \mem3_reg[179][31]  ( .D(n13899), .SI(\mem3[179][30] ), .SE(test_se), 
        .CLK(n1782), .Q(\mem3[179][31] ), .QN(n28257) );
  SDFFX1 \mem3_reg[179][30]  ( .D(n13898), .SI(\mem3[179][29] ), .SE(test_se), 
        .CLK(n1782), .Q(\mem3[179][30] ), .QN(n28258) );
  SDFFX1 \mem3_reg[179][29]  ( .D(n13897), .SI(\mem3[179][28] ), .SE(test_se), 
        .CLK(n1782), .Q(\mem3[179][29] ), .QN(n28259) );
  SDFFX1 \mem3_reg[179][28]  ( .D(n13896), .SI(\mem3[179][27] ), .SE(test_se), 
        .CLK(n1782), .Q(\mem3[179][28] ), .QN(n28260) );
  SDFFX1 \mem3_reg[179][27]  ( .D(n13895), .SI(\mem3[179][26] ), .SE(test_se), 
        .CLK(n1782), .Q(\mem3[179][27] ), .QN(n28261) );
  SDFFX1 \mem3_reg[179][26]  ( .D(n13894), .SI(\mem3[179][25] ), .SE(test_se), 
        .CLK(n1782), .Q(\mem3[179][26] ), .QN(n28262) );
  SDFFX1 \mem3_reg[179][25]  ( .D(n13893), .SI(\mem3[179][24] ), .SE(test_se), 
        .CLK(n1782), .Q(\mem3[179][25] ), .QN(n28263) );
  SDFFX1 \mem3_reg[179][24]  ( .D(n13892), .SI(\mem3[178][31] ), .SE(test_se), 
        .CLK(n1782), .Q(\mem3[179][24] ), .QN(n28264) );
  SDFFX1 \mem3_reg[178][31]  ( .D(n13891), .SI(\mem3[178][30] ), .SE(test_se), 
        .CLK(n1782), .Q(\mem3[178][31] ), .QN(n28265) );
  SDFFX1 \mem3_reg[178][30]  ( .D(n13890), .SI(\mem3[178][29] ), .SE(test_se), 
        .CLK(n1782), .Q(\mem3[178][30] ), .QN(n28266) );
  SDFFX1 \mem3_reg[178][29]  ( .D(n13889), .SI(\mem3[178][28] ), .SE(test_se), 
        .CLK(n1782), .Q(\mem3[178][29] ), .QN(n28267) );
  SDFFX1 \mem3_reg[178][28]  ( .D(n13888), .SI(\mem3[178][27] ), .SE(test_se), 
        .CLK(n1783), .Q(\mem3[178][28] ), .QN(n28268) );
  SDFFX1 \mem3_reg[178][27]  ( .D(n13887), .SI(\mem3[178][26] ), .SE(test_se), 
        .CLK(n1783), .Q(\mem3[178][27] ), .QN(n28269) );
  SDFFX1 \mem3_reg[178][26]  ( .D(n13886), .SI(\mem3[178][25] ), .SE(test_se), 
        .CLK(n1783), .Q(\mem3[178][26] ), .QN(n28270) );
  SDFFX1 \mem3_reg[178][25]  ( .D(n13885), .SI(\mem3[178][24] ), .SE(test_se), 
        .CLK(n1783), .Q(\mem3[178][25] ), .QN(n28271) );
  SDFFX1 \mem3_reg[178][24]  ( .D(n13884), .SI(\mem3[177][31] ), .SE(test_se), 
        .CLK(n1783), .Q(\mem3[178][24] ), .QN(n28272) );
  SDFFX1 \mem3_reg[177][31]  ( .D(n13883), .SI(\mem3[177][30] ), .SE(test_se), 
        .CLK(n1783), .Q(\mem3[177][31] ), .QN(n28273) );
  SDFFX1 \mem3_reg[177][30]  ( .D(n13882), .SI(\mem3[177][29] ), .SE(test_se), 
        .CLK(n1783), .Q(\mem3[177][30] ), .QN(n28274) );
  SDFFX1 \mem3_reg[177][29]  ( .D(n13881), .SI(\mem3[177][28] ), .SE(test_se), 
        .CLK(n1783), .Q(\mem3[177][29] ), .QN(n28275) );
  SDFFX1 \mem3_reg[177][28]  ( .D(n13880), .SI(\mem3[177][27] ), .SE(test_se), 
        .CLK(n1783), .Q(\mem3[177][28] ), .QN(n28276) );
  SDFFX1 \mem3_reg[177][27]  ( .D(n13879), .SI(\mem3[177][26] ), .SE(test_se), 
        .CLK(n1783), .Q(\mem3[177][27] ), .QN(n28277) );
  SDFFX1 \mem3_reg[177][26]  ( .D(n13878), .SI(\mem3[177][25] ), .SE(test_se), 
        .CLK(n1783), .Q(\mem3[177][26] ), .QN(n28278) );
  SDFFX1 \mem3_reg[177][25]  ( .D(n13877), .SI(\mem3[177][24] ), .SE(test_se), 
        .CLK(n1783), .Q(\mem3[177][25] ), .QN(n28279) );
  SDFFX1 \mem3_reg[177][24]  ( .D(n13876), .SI(\mem3[176][31] ), .SE(test_se), 
        .CLK(n1784), .Q(\mem3[177][24] ), .QN(n28280) );
  SDFFX1 \mem3_reg[176][31]  ( .D(n13875), .SI(\mem3[176][30] ), .SE(test_se), 
        .CLK(n1784), .Q(\mem3[176][31] ), .QN(n28281) );
  SDFFX1 \mem3_reg[176][30]  ( .D(n13874), .SI(\mem3[176][29] ), .SE(test_se), 
        .CLK(n1784), .Q(\mem3[176][30] ), .QN(n28282) );
  SDFFX1 \mem3_reg[176][29]  ( .D(n13873), .SI(\mem3[176][28] ), .SE(test_se), 
        .CLK(n1784), .Q(\mem3[176][29] ), .QN(n28283) );
  SDFFX1 \mem3_reg[176][28]  ( .D(n13872), .SI(\mem3[176][27] ), .SE(test_se), 
        .CLK(n1784), .Q(\mem3[176][28] ), .QN(n28284) );
  SDFFX1 \mem3_reg[176][27]  ( .D(n13871), .SI(\mem3[176][26] ), .SE(test_se), 
        .CLK(n1784), .Q(\mem3[176][27] ), .QN(n28285) );
  SDFFX1 \mem3_reg[176][26]  ( .D(n13870), .SI(\mem3[176][25] ), .SE(test_se), 
        .CLK(n1784), .Q(\mem3[176][26] ), .QN(n28286) );
  SDFFX1 \mem3_reg[176][25]  ( .D(n13869), .SI(\mem3[176][24] ), .SE(test_se), 
        .CLK(n1784), .Q(\mem3[176][25] ), .QN(n28287) );
  SDFFX1 \mem3_reg[176][24]  ( .D(n13868), .SI(\mem3[175][31] ), .SE(test_se), 
        .CLK(n1784), .Q(\mem3[176][24] ), .QN(n28288) );
  SDFFX1 \mem3_reg[175][31]  ( .D(n13867), .SI(\mem3[175][30] ), .SE(test_se), 
        .CLK(n1784), .Q(\mem3[175][31] ), .QN(n28289) );
  SDFFX1 \mem3_reg[175][30]  ( .D(n13866), .SI(\mem3[175][29] ), .SE(test_se), 
        .CLK(n1784), .Q(\mem3[175][30] ), .QN(n28290) );
  SDFFX1 \mem3_reg[175][29]  ( .D(n13865), .SI(\mem3[175][28] ), .SE(test_se), 
        .CLK(n1784), .Q(\mem3[175][29] ), .QN(n28291) );
  SDFFX1 \mem3_reg[175][28]  ( .D(n13864), .SI(\mem3[175][27] ), .SE(test_se), 
        .CLK(n1785), .Q(\mem3[175][28] ), .QN(n28292) );
  SDFFX1 \mem3_reg[175][27]  ( .D(n13863), .SI(\mem3[175][26] ), .SE(test_se), 
        .CLK(n1785), .Q(\mem3[175][27] ), .QN(n28293) );
  SDFFX1 \mem3_reg[175][26]  ( .D(n13862), .SI(\mem3[175][25] ), .SE(test_se), 
        .CLK(n1785), .Q(\mem3[175][26] ), .QN(n28294) );
  SDFFX1 \mem3_reg[175][25]  ( .D(n13861), .SI(\mem3[175][24] ), .SE(test_se), 
        .CLK(n1785), .Q(\mem3[175][25] ), .QN(n28295) );
  SDFFX1 \mem3_reg[175][24]  ( .D(n13860), .SI(\mem3[174][31] ), .SE(test_se), 
        .CLK(n1785), .Q(\mem3[175][24] ), .QN(n28296) );
  SDFFX1 \mem3_reg[174][31]  ( .D(n13859), .SI(\mem3[174][30] ), .SE(test_se), 
        .CLK(n1785), .Q(\mem3[174][31] ), .QN(n28297) );
  SDFFX1 \mem3_reg[174][30]  ( .D(n13858), .SI(\mem3[174][29] ), .SE(test_se), 
        .CLK(n1785), .Q(\mem3[174][30] ), .QN(n28298) );
  SDFFX1 \mem3_reg[174][29]  ( .D(n13857), .SI(\mem3[174][28] ), .SE(test_se), 
        .CLK(n1785), .Q(\mem3[174][29] ), .QN(n28299) );
  SDFFX1 \mem3_reg[174][28]  ( .D(n13856), .SI(\mem3[174][27] ), .SE(test_se), 
        .CLK(n1785), .Q(\mem3[174][28] ), .QN(n28300) );
  SDFFX1 \mem3_reg[174][27]  ( .D(n13855), .SI(\mem3[174][26] ), .SE(test_se), 
        .CLK(n1785), .Q(\mem3[174][27] ), .QN(n28301) );
  SDFFX1 \mem3_reg[174][26]  ( .D(n13854), .SI(\mem3[174][25] ), .SE(test_se), 
        .CLK(n1785), .Q(\mem3[174][26] ), .QN(n28302) );
  SDFFX1 \mem3_reg[174][25]  ( .D(n13853), .SI(\mem3[174][24] ), .SE(test_se), 
        .CLK(n1785), .Q(\mem3[174][25] ), .QN(n28303) );
  SDFFX1 \mem3_reg[174][24]  ( .D(n13852), .SI(\mem3[173][31] ), .SE(test_se), 
        .CLK(n1786), .Q(\mem3[174][24] ), .QN(n28304) );
  SDFFX1 \mem3_reg[173][31]  ( .D(n13851), .SI(\mem3[173][30] ), .SE(test_se), 
        .CLK(n1786), .Q(\mem3[173][31] ), .QN(n28305) );
  SDFFX1 \mem3_reg[173][30]  ( .D(n13850), .SI(\mem3[173][29] ), .SE(test_se), 
        .CLK(n1786), .Q(\mem3[173][30] ), .QN(n28306) );
  SDFFX1 \mem3_reg[173][29]  ( .D(n13849), .SI(\mem3[173][28] ), .SE(test_se), 
        .CLK(n1786), .Q(\mem3[173][29] ), .QN(n28307) );
  SDFFX1 \mem3_reg[173][28]  ( .D(n13848), .SI(\mem3[173][27] ), .SE(test_se), 
        .CLK(n1786), .Q(\mem3[173][28] ), .QN(n28308) );
  SDFFX1 \mem3_reg[173][27]  ( .D(n13847), .SI(\mem3[173][26] ), .SE(test_se), 
        .CLK(n1786), .Q(\mem3[173][27] ), .QN(n28309) );
  SDFFX1 \mem3_reg[173][26]  ( .D(n13846), .SI(\mem3[173][25] ), .SE(test_se), 
        .CLK(n1786), .Q(\mem3[173][26] ), .QN(n28310) );
  SDFFX1 \mem3_reg[173][25]  ( .D(n13845), .SI(\mem3[173][24] ), .SE(test_se), 
        .CLK(n1786), .Q(\mem3[173][25] ), .QN(n28311) );
  SDFFX1 \mem3_reg[173][24]  ( .D(n13844), .SI(\mem3[172][31] ), .SE(test_se), 
        .CLK(n1786), .Q(\mem3[173][24] ), .QN(n28312) );
  SDFFX1 \mem3_reg[172][31]  ( .D(n13843), .SI(\mem3[172][30] ), .SE(test_se), 
        .CLK(n1786), .Q(\mem3[172][31] ), .QN(n28313) );
  SDFFX1 \mem3_reg[172][30]  ( .D(n13842), .SI(\mem3[172][29] ), .SE(test_se), 
        .CLK(n1786), .Q(\mem3[172][30] ), .QN(n28314) );
  SDFFX1 \mem3_reg[172][29]  ( .D(n13841), .SI(\mem3[172][28] ), .SE(test_se), 
        .CLK(n1786), .Q(\mem3[172][29] ), .QN(n28315) );
  SDFFX1 \mem3_reg[172][28]  ( .D(n13840), .SI(\mem3[172][27] ), .SE(test_se), 
        .CLK(n1787), .Q(\mem3[172][28] ), .QN(n28316) );
  SDFFX1 \mem3_reg[172][27]  ( .D(n13839), .SI(\mem3[172][26] ), .SE(test_se), 
        .CLK(n1787), .Q(\mem3[172][27] ), .QN(n28317) );
  SDFFX1 \mem3_reg[172][26]  ( .D(n13838), .SI(\mem3[172][25] ), .SE(test_se), 
        .CLK(n1787), .Q(\mem3[172][26] ), .QN(n28318) );
  SDFFX1 \mem3_reg[172][25]  ( .D(n13837), .SI(\mem3[172][24] ), .SE(test_se), 
        .CLK(n1787), .Q(\mem3[172][25] ), .QN(n28319) );
  SDFFX1 \mem3_reg[172][24]  ( .D(n13836), .SI(\mem3[171][31] ), .SE(test_se), 
        .CLK(n1787), .Q(\mem3[172][24] ), .QN(n28320) );
  SDFFX1 \mem3_reg[171][31]  ( .D(n13835), .SI(\mem3[171][30] ), .SE(test_se), 
        .CLK(n1787), .Q(\mem3[171][31] ), .QN(n28321) );
  SDFFX1 \mem3_reg[171][30]  ( .D(n13834), .SI(\mem3[171][29] ), .SE(test_se), 
        .CLK(n1787), .Q(\mem3[171][30] ), .QN(n28322) );
  SDFFX1 \mem3_reg[171][29]  ( .D(n13833), .SI(\mem3[171][28] ), .SE(test_se), 
        .CLK(n1787), .Q(\mem3[171][29] ), .QN(n28323) );
  SDFFX1 \mem3_reg[171][28]  ( .D(n13832), .SI(\mem3[171][27] ), .SE(test_se), 
        .CLK(n1787), .Q(\mem3[171][28] ), .QN(n28324) );
  SDFFX1 \mem3_reg[171][27]  ( .D(n13831), .SI(\mem3[171][26] ), .SE(test_se), 
        .CLK(n1787), .Q(\mem3[171][27] ), .QN(n28325) );
  SDFFX1 \mem3_reg[171][26]  ( .D(n13830), .SI(\mem3[171][25] ), .SE(test_se), 
        .CLK(n1787), .Q(\mem3[171][26] ), .QN(n28326) );
  SDFFX1 \mem3_reg[171][25]  ( .D(n13829), .SI(\mem3[171][24] ), .SE(test_se), 
        .CLK(n1787), .Q(\mem3[171][25] ), .QN(n28327) );
  SDFFX1 \mem3_reg[171][24]  ( .D(n13828), .SI(\mem3[170][31] ), .SE(test_se), 
        .CLK(n1788), .Q(\mem3[171][24] ), .QN(n28328) );
  SDFFX1 \mem3_reg[170][31]  ( .D(n13827), .SI(\mem3[170][30] ), .SE(test_se), 
        .CLK(n1788), .Q(\mem3[170][31] ), .QN(n28329) );
  SDFFX1 \mem3_reg[170][30]  ( .D(n13826), .SI(\mem3[170][29] ), .SE(test_se), 
        .CLK(n1788), .Q(\mem3[170][30] ), .QN(n28330) );
  SDFFX1 \mem3_reg[170][29]  ( .D(n13825), .SI(\mem3[170][28] ), .SE(test_se), 
        .CLK(n1788), .Q(\mem3[170][29] ), .QN(n28331) );
  SDFFX1 \mem3_reg[170][28]  ( .D(n13824), .SI(\mem3[170][27] ), .SE(test_se), 
        .CLK(n1788), .Q(\mem3[170][28] ), .QN(n28332) );
  SDFFX1 \mem3_reg[170][27]  ( .D(n13823), .SI(\mem3[170][26] ), .SE(test_se), 
        .CLK(n1788), .Q(\mem3[170][27] ), .QN(n28333) );
  SDFFX1 \mem3_reg[170][26]  ( .D(n13822), .SI(\mem3[170][25] ), .SE(test_se), 
        .CLK(n1788), .Q(\mem3[170][26] ), .QN(n28334) );
  SDFFX1 \mem3_reg[170][25]  ( .D(n13821), .SI(\mem3[170][24] ), .SE(test_se), 
        .CLK(n1788), .Q(\mem3[170][25] ), .QN(n28335) );
  SDFFX1 \mem3_reg[170][24]  ( .D(n13820), .SI(\mem3[169][31] ), .SE(test_se), 
        .CLK(n1788), .Q(\mem3[170][24] ), .QN(n28336) );
  SDFFX1 \mem3_reg[169][31]  ( .D(n13819), .SI(\mem3[169][30] ), .SE(test_se), 
        .CLK(n1788), .Q(\mem3[169][31] ), .QN(n28337) );
  SDFFX1 \mem3_reg[169][30]  ( .D(n13818), .SI(\mem3[169][29] ), .SE(test_se), 
        .CLK(n1788), .Q(\mem3[169][30] ), .QN(n28338) );
  SDFFX1 \mem3_reg[169][29]  ( .D(n13817), .SI(\mem3[169][28] ), .SE(test_se), 
        .CLK(n1788), .Q(\mem3[169][29] ), .QN(n28339) );
  SDFFX1 \mem3_reg[169][28]  ( .D(n13816), .SI(\mem3[169][27] ), .SE(test_se), 
        .CLK(n1789), .Q(\mem3[169][28] ), .QN(n28340) );
  SDFFX1 \mem3_reg[169][27]  ( .D(n13815), .SI(\mem3[169][26] ), .SE(test_se), 
        .CLK(n1789), .Q(\mem3[169][27] ), .QN(n28341) );
  SDFFX1 \mem3_reg[169][26]  ( .D(n13814), .SI(\mem3[169][25] ), .SE(test_se), 
        .CLK(n1789), .Q(\mem3[169][26] ), .QN(n28342) );
  SDFFX1 \mem3_reg[169][25]  ( .D(n13813), .SI(\mem3[169][24] ), .SE(test_se), 
        .CLK(n1789), .Q(\mem3[169][25] ), .QN(n28343) );
  SDFFX1 \mem3_reg[169][24]  ( .D(n13812), .SI(\mem3[168][31] ), .SE(test_se), 
        .CLK(n1789), .Q(\mem3[169][24] ), .QN(n28344) );
  SDFFX1 \mem3_reg[168][31]  ( .D(n13811), .SI(\mem3[168][30] ), .SE(test_se), 
        .CLK(n1789), .Q(\mem3[168][31] ), .QN(n28345) );
  SDFFX1 \mem3_reg[168][30]  ( .D(n13810), .SI(\mem3[168][29] ), .SE(test_se), 
        .CLK(n1789), .Q(\mem3[168][30] ), .QN(n28346) );
  SDFFX1 \mem3_reg[168][29]  ( .D(n13809), .SI(\mem3[168][28] ), .SE(test_se), 
        .CLK(n1789), .Q(\mem3[168][29] ), .QN(n28347) );
  SDFFX1 \mem3_reg[168][28]  ( .D(n13808), .SI(\mem3[168][27] ), .SE(test_se), 
        .CLK(n1789), .Q(\mem3[168][28] ), .QN(n28348) );
  SDFFX1 \mem3_reg[168][27]  ( .D(n13807), .SI(\mem3[168][26] ), .SE(test_se), 
        .CLK(n1789), .Q(\mem3[168][27] ), .QN(n28349) );
  SDFFX1 \mem3_reg[168][26]  ( .D(n13806), .SI(\mem3[168][25] ), .SE(test_se), 
        .CLK(n1789), .Q(\mem3[168][26] ), .QN(n28350) );
  SDFFX1 \mem3_reg[168][25]  ( .D(n13805), .SI(\mem3[168][24] ), .SE(test_se), 
        .CLK(n1789), .Q(\mem3[168][25] ), .QN(n28351) );
  SDFFX1 \mem3_reg[168][24]  ( .D(n13804), .SI(\mem3[167][31] ), .SE(test_se), 
        .CLK(n1790), .Q(\mem3[168][24] ), .QN(n28352) );
  SDFFX1 \mem3_reg[167][31]  ( .D(n13803), .SI(\mem3[167][30] ), .SE(test_se), 
        .CLK(n1790), .Q(\mem3[167][31] ), .QN(n28353) );
  SDFFX1 \mem3_reg[167][30]  ( .D(n13802), .SI(\mem3[167][29] ), .SE(test_se), 
        .CLK(n1790), .Q(\mem3[167][30] ), .QN(n28354) );
  SDFFX1 \mem3_reg[167][29]  ( .D(n13801), .SI(\mem3[167][28] ), .SE(test_se), 
        .CLK(n1790), .Q(\mem3[167][29] ), .QN(n28355) );
  SDFFX1 \mem3_reg[167][28]  ( .D(n13800), .SI(\mem3[167][27] ), .SE(test_se), 
        .CLK(n1790), .Q(\mem3[167][28] ), .QN(n28356) );
  SDFFX1 \mem3_reg[167][27]  ( .D(n13799), .SI(\mem3[167][26] ), .SE(test_se), 
        .CLK(n1790), .Q(\mem3[167][27] ), .QN(n28357) );
  SDFFX1 \mem3_reg[167][26]  ( .D(n13798), .SI(\mem3[167][25] ), .SE(test_se), 
        .CLK(n1790), .Q(\mem3[167][26] ), .QN(n28358) );
  SDFFX1 \mem3_reg[167][25]  ( .D(n13797), .SI(\mem3[167][24] ), .SE(test_se), 
        .CLK(n1790), .Q(\mem3[167][25] ), .QN(n28359) );
  SDFFX1 \mem3_reg[167][24]  ( .D(n13796), .SI(\mem3[166][31] ), .SE(test_se), 
        .CLK(n1790), .Q(\mem3[167][24] ), .QN(n28360) );
  SDFFX1 \mem3_reg[166][31]  ( .D(n13795), .SI(\mem3[166][30] ), .SE(test_se), 
        .CLK(n1790), .Q(\mem3[166][31] ), .QN(n28361) );
  SDFFX1 \mem3_reg[166][30]  ( .D(n13794), .SI(\mem3[166][29] ), .SE(test_se), 
        .CLK(n1790), .Q(\mem3[166][30] ), .QN(n28362) );
  SDFFX1 \mem3_reg[166][29]  ( .D(n13793), .SI(\mem3[166][28] ), .SE(test_se), 
        .CLK(n1790), .Q(\mem3[166][29] ), .QN(n28363) );
  SDFFX1 \mem3_reg[166][28]  ( .D(n13792), .SI(\mem3[166][27] ), .SE(test_se), 
        .CLK(n1791), .Q(\mem3[166][28] ), .QN(n28364) );
  SDFFX1 \mem3_reg[166][27]  ( .D(n13791), .SI(\mem3[166][26] ), .SE(test_se), 
        .CLK(n1791), .Q(\mem3[166][27] ), .QN(n28365) );
  SDFFX1 \mem3_reg[166][26]  ( .D(n13790), .SI(\mem3[166][25] ), .SE(test_se), 
        .CLK(n1791), .Q(\mem3[166][26] ), .QN(n28366) );
  SDFFX1 \mem3_reg[166][25]  ( .D(n13789), .SI(\mem3[166][24] ), .SE(test_se), 
        .CLK(n1791), .Q(\mem3[166][25] ), .QN(n28367) );
  SDFFX1 \mem3_reg[166][24]  ( .D(n13788), .SI(\mem3[165][31] ), .SE(test_se), 
        .CLK(n1791), .Q(\mem3[166][24] ), .QN(n28368) );
  SDFFX1 \mem3_reg[165][31]  ( .D(n13787), .SI(\mem3[165][30] ), .SE(test_se), 
        .CLK(n1791), .Q(\mem3[165][31] ), .QN(n28369) );
  SDFFX1 \mem3_reg[165][30]  ( .D(n13786), .SI(\mem3[165][29] ), .SE(test_se), 
        .CLK(n1791), .Q(\mem3[165][30] ), .QN(n28370) );
  SDFFX1 \mem3_reg[165][29]  ( .D(n13785), .SI(\mem3[165][28] ), .SE(test_se), 
        .CLK(n1791), .Q(\mem3[165][29] ), .QN(n28371) );
  SDFFX1 \mem3_reg[165][28]  ( .D(n13784), .SI(\mem3[165][27] ), .SE(test_se), 
        .CLK(n1791), .Q(\mem3[165][28] ), .QN(n28372) );
  SDFFX1 \mem3_reg[165][27]  ( .D(n13783), .SI(\mem3[165][26] ), .SE(test_se), 
        .CLK(n1791), .Q(\mem3[165][27] ), .QN(n28373) );
  SDFFX1 \mem3_reg[165][26]  ( .D(n13782), .SI(\mem3[165][25] ), .SE(test_se), 
        .CLK(n1791), .Q(\mem3[165][26] ), .QN(n28374) );
  SDFFX1 \mem3_reg[165][25]  ( .D(n13781), .SI(\mem3[165][24] ), .SE(test_se), 
        .CLK(n1791), .Q(\mem3[165][25] ), .QN(n28375) );
  SDFFX1 \mem3_reg[165][24]  ( .D(n13780), .SI(\mem3[164][31] ), .SE(test_se), 
        .CLK(n1792), .Q(\mem3[165][24] ), .QN(n28376) );
  SDFFX1 \mem3_reg[164][31]  ( .D(n13779), .SI(\mem3[164][30] ), .SE(test_se), 
        .CLK(n1792), .Q(\mem3[164][31] ), .QN(n28377) );
  SDFFX1 \mem3_reg[164][30]  ( .D(n13778), .SI(\mem3[164][29] ), .SE(test_se), 
        .CLK(n1792), .Q(\mem3[164][30] ), .QN(n28378) );
  SDFFX1 \mem3_reg[164][29]  ( .D(n13777), .SI(\mem3[164][28] ), .SE(test_se), 
        .CLK(n1792), .Q(\mem3[164][29] ), .QN(n28379) );
  SDFFX1 \mem3_reg[164][28]  ( .D(n13776), .SI(\mem3[164][27] ), .SE(test_se), 
        .CLK(n1792), .Q(\mem3[164][28] ), .QN(n28380) );
  SDFFX1 \mem3_reg[164][27]  ( .D(n13775), .SI(\mem3[164][26] ), .SE(test_se), 
        .CLK(n1792), .Q(\mem3[164][27] ), .QN(n28381) );
  SDFFX1 \mem3_reg[164][26]  ( .D(n13774), .SI(\mem3[164][25] ), .SE(test_se), 
        .CLK(n1792), .Q(\mem3[164][26] ), .QN(n28382) );
  SDFFX1 \mem3_reg[164][25]  ( .D(n13773), .SI(\mem3[164][24] ), .SE(test_se), 
        .CLK(n1792), .Q(\mem3[164][25] ), .QN(n28383) );
  SDFFX1 \mem3_reg[164][24]  ( .D(n13772), .SI(\mem3[163][31] ), .SE(test_se), 
        .CLK(n1792), .Q(\mem3[164][24] ), .QN(n28384) );
  SDFFX1 \mem3_reg[163][31]  ( .D(n13771), .SI(\mem3[163][30] ), .SE(test_se), 
        .CLK(n1792), .Q(\mem3[163][31] ), .QN(n28385) );
  SDFFX1 \mem3_reg[163][30]  ( .D(n13770), .SI(\mem3[163][29] ), .SE(test_se), 
        .CLK(n1792), .Q(\mem3[163][30] ), .QN(n28386) );
  SDFFX1 \mem3_reg[163][29]  ( .D(n13769), .SI(\mem3[163][28] ), .SE(test_se), 
        .CLK(n1792), .Q(\mem3[163][29] ), .QN(n28387) );
  SDFFX1 \mem3_reg[163][28]  ( .D(n13768), .SI(\mem3[163][27] ), .SE(test_se), 
        .CLK(n1793), .Q(\mem3[163][28] ), .QN(n28388) );
  SDFFX1 \mem3_reg[163][27]  ( .D(n13767), .SI(\mem3[163][26] ), .SE(test_se), 
        .CLK(n1793), .Q(\mem3[163][27] ), .QN(n28389) );
  SDFFX1 \mem3_reg[163][26]  ( .D(n13766), .SI(\mem3[163][25] ), .SE(test_se), 
        .CLK(n1793), .Q(\mem3[163][26] ), .QN(n28390) );
  SDFFX1 \mem3_reg[163][25]  ( .D(n13765), .SI(\mem3[163][24] ), .SE(test_se), 
        .CLK(n1793), .Q(\mem3[163][25] ), .QN(n28391) );
  SDFFX1 \mem3_reg[163][24]  ( .D(n13764), .SI(\mem3[162][31] ), .SE(test_se), 
        .CLK(n1793), .Q(\mem3[163][24] ), .QN(n28392) );
  SDFFX1 \mem3_reg[162][31]  ( .D(n13763), .SI(\mem3[162][30] ), .SE(test_se), 
        .CLK(n1793), .Q(\mem3[162][31] ), .QN(n28393) );
  SDFFX1 \mem3_reg[162][30]  ( .D(n13762), .SI(\mem3[162][29] ), .SE(test_se), 
        .CLK(n1793), .Q(\mem3[162][30] ), .QN(n28394) );
  SDFFX1 \mem3_reg[162][29]  ( .D(n13761), .SI(\mem3[162][28] ), .SE(test_se), 
        .CLK(n1793), .Q(\mem3[162][29] ), .QN(n28395) );
  SDFFX1 \mem3_reg[162][28]  ( .D(n13760), .SI(\mem3[162][27] ), .SE(test_se), 
        .CLK(n1793), .Q(\mem3[162][28] ), .QN(n28396) );
  SDFFX1 \mem3_reg[162][27]  ( .D(n13759), .SI(\mem3[162][26] ), .SE(test_se), 
        .CLK(n1793), .Q(\mem3[162][27] ), .QN(n28397) );
  SDFFX1 \mem3_reg[162][26]  ( .D(n13758), .SI(\mem3[162][25] ), .SE(test_se), 
        .CLK(n1793), .Q(\mem3[162][26] ), .QN(n28398) );
  SDFFX1 \mem3_reg[162][25]  ( .D(n13757), .SI(\mem3[162][24] ), .SE(test_se), 
        .CLK(n1793), .Q(\mem3[162][25] ), .QN(n28399) );
  SDFFX1 \mem3_reg[162][24]  ( .D(n13756), .SI(\mem3[161][31] ), .SE(test_se), 
        .CLK(n1794), .Q(\mem3[162][24] ), .QN(n28400) );
  SDFFX1 \mem3_reg[161][31]  ( .D(n13755), .SI(\mem3[161][30] ), .SE(test_se), 
        .CLK(n1794), .Q(\mem3[161][31] ), .QN(n28401) );
  SDFFX1 \mem3_reg[161][30]  ( .D(n13754), .SI(\mem3[161][29] ), .SE(test_se), 
        .CLK(n1794), .Q(\mem3[161][30] ), .QN(n28402) );
  SDFFX1 \mem3_reg[161][29]  ( .D(n13753), .SI(\mem3[161][28] ), .SE(test_se), 
        .CLK(n1794), .Q(\mem3[161][29] ), .QN(n28403) );
  SDFFX1 \mem3_reg[161][28]  ( .D(n13752), .SI(\mem3[161][27] ), .SE(test_se), 
        .CLK(n1794), .Q(\mem3[161][28] ), .QN(n28404) );
  SDFFX1 \mem3_reg[161][27]  ( .D(n13751), .SI(\mem3[161][26] ), .SE(test_se), 
        .CLK(n1794), .Q(\mem3[161][27] ), .QN(n28405) );
  SDFFX1 \mem3_reg[161][26]  ( .D(n13750), .SI(\mem3[161][25] ), .SE(test_se), 
        .CLK(n1794), .Q(\mem3[161][26] ), .QN(n28406) );
  SDFFX1 \mem3_reg[161][25]  ( .D(n13749), .SI(\mem3[161][24] ), .SE(test_se), 
        .CLK(n1794), .Q(\mem3[161][25] ), .QN(n28407) );
  SDFFX1 \mem3_reg[161][24]  ( .D(n13748), .SI(\mem3[160][31] ), .SE(test_se), 
        .CLK(n1794), .Q(\mem3[161][24] ), .QN(n28408) );
  SDFFX1 \mem3_reg[160][31]  ( .D(n13747), .SI(\mem3[160][30] ), .SE(test_se), 
        .CLK(n1794), .Q(\mem3[160][31] ), .QN(n28409) );
  SDFFX1 \mem3_reg[160][30]  ( .D(n13746), .SI(\mem3[160][29] ), .SE(test_se), 
        .CLK(n1794), .Q(\mem3[160][30] ), .QN(n28410) );
  SDFFX1 \mem3_reg[160][29]  ( .D(n13745), .SI(\mem3[160][28] ), .SE(test_se), 
        .CLK(n1794), .Q(\mem3[160][29] ), .QN(n28411) );
  SDFFX1 \mem3_reg[160][28]  ( .D(n13744), .SI(\mem3[160][27] ), .SE(test_se), 
        .CLK(n1795), .Q(\mem3[160][28] ), .QN(n28412) );
  SDFFX1 \mem3_reg[160][27]  ( .D(n13743), .SI(\mem3[160][26] ), .SE(test_se), 
        .CLK(n1795), .Q(\mem3[160][27] ), .QN(n28413) );
  SDFFX1 \mem3_reg[160][26]  ( .D(n13742), .SI(\mem3[160][25] ), .SE(test_se), 
        .CLK(n1795), .Q(\mem3[160][26] ), .QN(n28414) );
  SDFFX1 \mem3_reg[160][25]  ( .D(n13741), .SI(\mem3[160][24] ), .SE(test_se), 
        .CLK(n1795), .Q(\mem3[160][25] ), .QN(n28415) );
  SDFFX1 \mem3_reg[160][24]  ( .D(n13740), .SI(\mem3[159][31] ), .SE(test_se), 
        .CLK(n1795), .Q(\mem3[160][24] ), .QN(n28416) );
  SDFFX1 \mem3_reg[159][31]  ( .D(n13739), .SI(\mem3[159][30] ), .SE(test_se), 
        .CLK(n1795), .Q(\mem3[159][31] ), .QN(n28417) );
  SDFFX1 \mem3_reg[159][30]  ( .D(n13738), .SI(\mem3[159][29] ), .SE(test_se), 
        .CLK(n1795), .Q(\mem3[159][30] ), .QN(n28418) );
  SDFFX1 \mem3_reg[159][29]  ( .D(n13737), .SI(\mem3[159][28] ), .SE(test_se), 
        .CLK(n1795), .Q(\mem3[159][29] ), .QN(n28419) );
  SDFFX1 \mem3_reg[159][28]  ( .D(n13736), .SI(\mem3[159][27] ), .SE(test_se), 
        .CLK(n1795), .Q(\mem3[159][28] ), .QN(n28420) );
  SDFFX1 \mem3_reg[159][27]  ( .D(n13735), .SI(\mem3[159][26] ), .SE(test_se), 
        .CLK(n1795), .Q(\mem3[159][27] ), .QN(n28421) );
  SDFFX1 \mem3_reg[159][26]  ( .D(n13734), .SI(\mem3[159][25] ), .SE(test_se), 
        .CLK(n1795), .Q(\mem3[159][26] ), .QN(n28422) );
  SDFFX1 \mem3_reg[159][25]  ( .D(n13733), .SI(\mem3[159][24] ), .SE(test_se), 
        .CLK(n1795), .Q(\mem3[159][25] ), .QN(n28423) );
  SDFFX1 \mem3_reg[159][24]  ( .D(n13732), .SI(\mem3[158][31] ), .SE(test_se), 
        .CLK(n1796), .Q(\mem3[159][24] ), .QN(n28424) );
  SDFFX1 \mem3_reg[158][31]  ( .D(n13731), .SI(\mem3[158][30] ), .SE(test_se), 
        .CLK(n1796), .Q(\mem3[158][31] ), .QN(n28425) );
  SDFFX1 \mem3_reg[158][30]  ( .D(n13730), .SI(\mem3[158][29] ), .SE(test_se), 
        .CLK(n1796), .Q(\mem3[158][30] ), .QN(n28426) );
  SDFFX1 \mem3_reg[158][29]  ( .D(n13729), .SI(\mem3[158][28] ), .SE(test_se), 
        .CLK(n1796), .Q(\mem3[158][29] ), .QN(n28427) );
  SDFFX1 \mem3_reg[158][28]  ( .D(n13728), .SI(\mem3[158][27] ), .SE(test_se), 
        .CLK(n1796), .Q(\mem3[158][28] ), .QN(n28428) );
  SDFFX1 \mem3_reg[158][27]  ( .D(n13727), .SI(\mem3[158][26] ), .SE(test_se), 
        .CLK(n1796), .Q(\mem3[158][27] ), .QN(n28429) );
  SDFFX1 \mem3_reg[158][26]  ( .D(n13726), .SI(\mem3[158][25] ), .SE(test_se), 
        .CLK(n1796), .Q(\mem3[158][26] ), .QN(n28430) );
  SDFFX1 \mem3_reg[158][25]  ( .D(n13725), .SI(\mem3[158][24] ), .SE(test_se), 
        .CLK(n1796), .Q(\mem3[158][25] ), .QN(n28431) );
  SDFFX1 \mem3_reg[158][24]  ( .D(n13724), .SI(\mem3[157][31] ), .SE(test_se), 
        .CLK(n1796), .Q(\mem3[158][24] ), .QN(n28432) );
  SDFFX1 \mem3_reg[157][31]  ( .D(n13723), .SI(\mem3[157][30] ), .SE(test_se), 
        .CLK(n1796), .Q(\mem3[157][31] ), .QN(n28433) );
  SDFFX1 \mem3_reg[157][30]  ( .D(n13722), .SI(\mem3[157][29] ), .SE(test_se), 
        .CLK(n1796), .Q(\mem3[157][30] ), .QN(n28434) );
  SDFFX1 \mem3_reg[157][29]  ( .D(n13721), .SI(\mem3[157][28] ), .SE(test_se), 
        .CLK(n1796), .Q(\mem3[157][29] ), .QN(n28435) );
  SDFFX1 \mem3_reg[157][28]  ( .D(n13720), .SI(\mem3[157][27] ), .SE(test_se), 
        .CLK(n1797), .Q(\mem3[157][28] ), .QN(n28436) );
  SDFFX1 \mem3_reg[157][27]  ( .D(n13719), .SI(\mem3[157][26] ), .SE(test_se), 
        .CLK(n1797), .Q(\mem3[157][27] ), .QN(n28437) );
  SDFFX1 \mem3_reg[157][26]  ( .D(n13718), .SI(\mem3[157][25] ), .SE(test_se), 
        .CLK(n1797), .Q(\mem3[157][26] ), .QN(n28438) );
  SDFFX1 \mem3_reg[157][25]  ( .D(n13717), .SI(\mem3[157][24] ), .SE(test_se), 
        .CLK(n1797), .Q(\mem3[157][25] ), .QN(n28439) );
  SDFFX1 \mem3_reg[157][24]  ( .D(n13716), .SI(\mem3[156][31] ), .SE(test_se), 
        .CLK(n1797), .Q(\mem3[157][24] ), .QN(n28440) );
  SDFFX1 \mem3_reg[156][31]  ( .D(n13715), .SI(\mem3[156][30] ), .SE(test_se), 
        .CLK(n1797), .Q(\mem3[156][31] ), .QN(n28441) );
  SDFFX1 \mem3_reg[156][30]  ( .D(n13714), .SI(\mem3[156][29] ), .SE(test_se), 
        .CLK(n1797), .Q(\mem3[156][30] ), .QN(n28442) );
  SDFFX1 \mem3_reg[156][29]  ( .D(n13713), .SI(\mem3[156][28] ), .SE(test_se), 
        .CLK(n1797), .Q(\mem3[156][29] ), .QN(n28443) );
  SDFFX1 \mem3_reg[156][28]  ( .D(n13712), .SI(\mem3[156][27] ), .SE(test_se), 
        .CLK(n1797), .Q(\mem3[156][28] ), .QN(n28444) );
  SDFFX1 \mem3_reg[156][27]  ( .D(n13711), .SI(\mem3[156][26] ), .SE(test_se), 
        .CLK(n1797), .Q(\mem3[156][27] ), .QN(n28445) );
  SDFFX1 \mem3_reg[156][26]  ( .D(n13710), .SI(\mem3[156][25] ), .SE(test_se), 
        .CLK(n1797), .Q(\mem3[156][26] ), .QN(n28446) );
  SDFFX1 \mem3_reg[156][25]  ( .D(n13709), .SI(\mem3[156][24] ), .SE(test_se), 
        .CLK(n1797), .Q(\mem3[156][25] ), .QN(n28447) );
  SDFFX1 \mem3_reg[156][24]  ( .D(n13708), .SI(\mem3[155][31] ), .SE(test_se), 
        .CLK(n1798), .Q(\mem3[156][24] ), .QN(n28448) );
  SDFFX1 \mem3_reg[155][31]  ( .D(n13707), .SI(\mem3[155][30] ), .SE(test_se), 
        .CLK(n1798), .Q(\mem3[155][31] ), .QN(n28449) );
  SDFFX1 \mem3_reg[155][30]  ( .D(n13706), .SI(\mem3[155][29] ), .SE(test_se), 
        .CLK(n1798), .Q(\mem3[155][30] ), .QN(n28450) );
  SDFFX1 \mem3_reg[155][29]  ( .D(n13705), .SI(\mem3[155][28] ), .SE(test_se), 
        .CLK(n1798), .Q(\mem3[155][29] ), .QN(n28451) );
  SDFFX1 \mem3_reg[155][28]  ( .D(n13704), .SI(\mem3[155][27] ), .SE(test_se), 
        .CLK(n1798), .Q(\mem3[155][28] ), .QN(n28452) );
  SDFFX1 \mem3_reg[155][27]  ( .D(n13703), .SI(\mem3[155][26] ), .SE(test_se), 
        .CLK(n1798), .Q(\mem3[155][27] ), .QN(n28453) );
  SDFFX1 \mem3_reg[155][26]  ( .D(n13702), .SI(\mem3[155][25] ), .SE(test_se), 
        .CLK(n1798), .Q(\mem3[155][26] ), .QN(n28454) );
  SDFFX1 \mem3_reg[155][25]  ( .D(n13701), .SI(\mem3[155][24] ), .SE(test_se), 
        .CLK(n1798), .Q(\mem3[155][25] ), .QN(n28455) );
  SDFFX1 \mem3_reg[155][24]  ( .D(n13700), .SI(\mem3[154][31] ), .SE(test_se), 
        .CLK(n1798), .Q(\mem3[155][24] ), .QN(n28456) );
  SDFFX1 \mem3_reg[154][31]  ( .D(n13699), .SI(\mem3[154][30] ), .SE(test_se), 
        .CLK(n1798), .Q(\mem3[154][31] ), .QN(n28457) );
  SDFFX1 \mem3_reg[154][30]  ( .D(n13698), .SI(\mem3[154][29] ), .SE(test_se), 
        .CLK(n1798), .Q(\mem3[154][30] ), .QN(n28458) );
  SDFFX1 \mem3_reg[154][29]  ( .D(n13697), .SI(\mem3[154][28] ), .SE(test_se), 
        .CLK(n1798), .Q(\mem3[154][29] ), .QN(n28459) );
  SDFFX1 \mem3_reg[154][28]  ( .D(n13696), .SI(\mem3[154][27] ), .SE(test_se), 
        .CLK(n1799), .Q(\mem3[154][28] ), .QN(n28460) );
  SDFFX1 \mem3_reg[154][27]  ( .D(n13695), .SI(\mem3[154][26] ), .SE(test_se), 
        .CLK(n1799), .Q(\mem3[154][27] ), .QN(n28461) );
  SDFFX1 \mem3_reg[154][26]  ( .D(n13694), .SI(\mem3[154][25] ), .SE(test_se), 
        .CLK(n1799), .Q(\mem3[154][26] ), .QN(n28462) );
  SDFFX1 \mem3_reg[154][25]  ( .D(n13693), .SI(\mem3[154][24] ), .SE(test_se), 
        .CLK(n1799), .Q(\mem3[154][25] ), .QN(n28463) );
  SDFFX1 \mem3_reg[154][24]  ( .D(n13692), .SI(\mem3[153][31] ), .SE(test_se), 
        .CLK(n1799), .Q(\mem3[154][24] ), .QN(n28464) );
  SDFFX1 \mem3_reg[153][31]  ( .D(n13691), .SI(\mem3[153][30] ), .SE(test_se), 
        .CLK(n1799), .Q(\mem3[153][31] ), .QN(n28465) );
  SDFFX1 \mem3_reg[153][30]  ( .D(n13690), .SI(\mem3[153][29] ), .SE(test_se), 
        .CLK(n1799), .Q(\mem3[153][30] ), .QN(n28466) );
  SDFFX1 \mem3_reg[153][29]  ( .D(n13689), .SI(\mem3[153][28] ), .SE(test_se), 
        .CLK(n1799), .Q(\mem3[153][29] ), .QN(n28467) );
  SDFFX1 \mem3_reg[153][28]  ( .D(n13688), .SI(\mem3[153][27] ), .SE(test_se), 
        .CLK(n1799), .Q(\mem3[153][28] ), .QN(n28468) );
  SDFFX1 \mem3_reg[153][27]  ( .D(n13687), .SI(\mem3[153][26] ), .SE(test_se), 
        .CLK(n1799), .Q(\mem3[153][27] ), .QN(n28469) );
  SDFFX1 \mem3_reg[153][26]  ( .D(n13686), .SI(\mem3[153][25] ), .SE(test_se), 
        .CLK(n1799), .Q(\mem3[153][26] ), .QN(n28470) );
  SDFFX1 \mem3_reg[153][25]  ( .D(n13685), .SI(\mem3[153][24] ), .SE(test_se), 
        .CLK(n1799), .Q(\mem3[153][25] ), .QN(n28471) );
  SDFFX1 \mem3_reg[153][24]  ( .D(n13684), .SI(\mem3[152][31] ), .SE(test_se), 
        .CLK(n1800), .Q(\mem3[153][24] ), .QN(n28472) );
  SDFFX1 \mem3_reg[152][31]  ( .D(n13683), .SI(\mem3[152][30] ), .SE(test_se), 
        .CLK(n1800), .Q(\mem3[152][31] ), .QN(n28473) );
  SDFFX1 \mem3_reg[152][30]  ( .D(n13682), .SI(\mem3[152][29] ), .SE(test_se), 
        .CLK(n1800), .Q(\mem3[152][30] ), .QN(n28474) );
  SDFFX1 \mem3_reg[152][29]  ( .D(n13681), .SI(\mem3[152][28] ), .SE(test_se), 
        .CLK(n1800), .Q(\mem3[152][29] ), .QN(n28475) );
  SDFFX1 \mem3_reg[152][28]  ( .D(n13680), .SI(\mem3[152][27] ), .SE(test_se), 
        .CLK(n1800), .Q(\mem3[152][28] ), .QN(n28476) );
  SDFFX1 \mem3_reg[152][27]  ( .D(n13679), .SI(\mem3[152][26] ), .SE(test_se), 
        .CLK(n1800), .Q(\mem3[152][27] ), .QN(n28477) );
  SDFFX1 \mem3_reg[152][26]  ( .D(n13678), .SI(\mem3[152][25] ), .SE(test_se), 
        .CLK(n1800), .Q(\mem3[152][26] ), .QN(n28478) );
  SDFFX1 \mem3_reg[152][25]  ( .D(n13677), .SI(\mem3[152][24] ), .SE(test_se), 
        .CLK(n1800), .Q(\mem3[152][25] ), .QN(n28479) );
  SDFFX1 \mem3_reg[152][24]  ( .D(n13676), .SI(\mem3[151][31] ), .SE(test_se), 
        .CLK(n1800), .Q(\mem3[152][24] ), .QN(n28480) );
  SDFFX1 \mem3_reg[151][31]  ( .D(n13675), .SI(\mem3[151][30] ), .SE(test_se), 
        .CLK(n1800), .Q(\mem3[151][31] ), .QN(n28481) );
  SDFFX1 \mem3_reg[151][30]  ( .D(n13674), .SI(\mem3[151][29] ), .SE(test_se), 
        .CLK(n1800), .Q(\mem3[151][30] ), .QN(n28482) );
  SDFFX1 \mem3_reg[151][29]  ( .D(n13673), .SI(\mem3[151][28] ), .SE(test_se), 
        .CLK(n1800), .Q(\mem3[151][29] ), .QN(n28483) );
  SDFFX1 \mem3_reg[151][28]  ( .D(n13672), .SI(\mem3[151][27] ), .SE(test_se), 
        .CLK(n1801), .Q(\mem3[151][28] ), .QN(n28484) );
  SDFFX1 \mem3_reg[151][27]  ( .D(n13671), .SI(\mem3[151][26] ), .SE(test_se), 
        .CLK(n1801), .Q(\mem3[151][27] ), .QN(n28485) );
  SDFFX1 \mem3_reg[151][26]  ( .D(n13670), .SI(\mem3[151][25] ), .SE(test_se), 
        .CLK(n1801), .Q(\mem3[151][26] ), .QN(n28486) );
  SDFFX1 \mem3_reg[151][25]  ( .D(n13669), .SI(\mem3[151][24] ), .SE(test_se), 
        .CLK(n1801), .Q(\mem3[151][25] ), .QN(n28487) );
  SDFFX1 \mem3_reg[151][24]  ( .D(n13668), .SI(\mem3[150][31] ), .SE(test_se), 
        .CLK(n1801), .Q(\mem3[151][24] ), .QN(n28488) );
  SDFFX1 \mem3_reg[150][31]  ( .D(n13667), .SI(\mem3[150][30] ), .SE(test_se), 
        .CLK(n1801), .Q(\mem3[150][31] ), .QN(n28489) );
  SDFFX1 \mem3_reg[150][30]  ( .D(n13666), .SI(\mem3[150][29] ), .SE(test_se), 
        .CLK(n1801), .Q(\mem3[150][30] ), .QN(n28490) );
  SDFFX1 \mem3_reg[150][29]  ( .D(n13665), .SI(\mem3[150][28] ), .SE(test_se), 
        .CLK(n1801), .Q(\mem3[150][29] ), .QN(n28491) );
  SDFFX1 \mem3_reg[150][28]  ( .D(n13664), .SI(\mem3[150][27] ), .SE(test_se), 
        .CLK(n1801), .Q(\mem3[150][28] ), .QN(n28492) );
  SDFFX1 \mem3_reg[150][27]  ( .D(n13663), .SI(\mem3[150][26] ), .SE(test_se), 
        .CLK(n1801), .Q(\mem3[150][27] ), .QN(n28493) );
  SDFFX1 \mem3_reg[150][26]  ( .D(n13662), .SI(\mem3[150][25] ), .SE(test_se), 
        .CLK(n1801), .Q(\mem3[150][26] ), .QN(n28494) );
  SDFFX1 \mem3_reg[150][25]  ( .D(n13661), .SI(\mem3[150][24] ), .SE(test_se), 
        .CLK(n1801), .Q(\mem3[150][25] ), .QN(n28495) );
  SDFFX1 \mem3_reg[150][24]  ( .D(n13660), .SI(\mem3[149][31] ), .SE(test_se), 
        .CLK(n1802), .Q(\mem3[150][24] ), .QN(n28496) );
  SDFFX1 \mem3_reg[149][31]  ( .D(n13659), .SI(\mem3[149][30] ), .SE(test_se), 
        .CLK(n1802), .Q(\mem3[149][31] ), .QN(n28497) );
  SDFFX1 \mem3_reg[149][30]  ( .D(n13658), .SI(\mem3[149][29] ), .SE(test_se), 
        .CLK(n1802), .Q(\mem3[149][30] ), .QN(n28498) );
  SDFFX1 \mem3_reg[149][29]  ( .D(n13657), .SI(\mem3[149][28] ), .SE(test_se), 
        .CLK(n1802), .Q(\mem3[149][29] ), .QN(n28499) );
  SDFFX1 \mem3_reg[149][28]  ( .D(n13656), .SI(\mem3[149][27] ), .SE(test_se), 
        .CLK(n1802), .Q(\mem3[149][28] ), .QN(n28500) );
  SDFFX1 \mem3_reg[149][27]  ( .D(n13655), .SI(\mem3[149][26] ), .SE(test_se), 
        .CLK(n1802), .Q(\mem3[149][27] ), .QN(n28501) );
  SDFFX1 \mem3_reg[149][26]  ( .D(n13654), .SI(\mem3[149][25] ), .SE(test_se), 
        .CLK(n1802), .Q(\mem3[149][26] ), .QN(n28502) );
  SDFFX1 \mem3_reg[149][25]  ( .D(n13653), .SI(\mem3[149][24] ), .SE(test_se), 
        .CLK(n1802), .Q(\mem3[149][25] ), .QN(n28503) );
  SDFFX1 \mem3_reg[149][24]  ( .D(n13652), .SI(\mem3[148][31] ), .SE(test_se), 
        .CLK(n1802), .Q(\mem3[149][24] ), .QN(n28504) );
  SDFFX1 \mem3_reg[148][31]  ( .D(n13651), .SI(\mem3[148][30] ), .SE(test_se), 
        .CLK(n1802), .Q(\mem3[148][31] ), .QN(n28505) );
  SDFFX1 \mem3_reg[148][30]  ( .D(n13650), .SI(\mem3[148][29] ), .SE(test_se), 
        .CLK(n1802), .Q(\mem3[148][30] ), .QN(n28506) );
  SDFFX1 \mem3_reg[148][29]  ( .D(n13649), .SI(\mem3[148][28] ), .SE(test_se), 
        .CLK(n1802), .Q(\mem3[148][29] ), .QN(n28507) );
  SDFFX1 \mem3_reg[148][28]  ( .D(n13648), .SI(\mem3[148][27] ), .SE(test_se), 
        .CLK(n1803), .Q(\mem3[148][28] ), .QN(n28508) );
  SDFFX1 \mem3_reg[148][27]  ( .D(n13647), .SI(\mem3[148][26] ), .SE(test_se), 
        .CLK(n1803), .Q(\mem3[148][27] ), .QN(n28509) );
  SDFFX1 \mem3_reg[148][26]  ( .D(n13646), .SI(\mem3[148][25] ), .SE(test_se), 
        .CLK(n1803), .Q(\mem3[148][26] ), .QN(n28510) );
  SDFFX1 \mem3_reg[148][25]  ( .D(n13645), .SI(\mem3[148][24] ), .SE(test_se), 
        .CLK(n1803), .Q(\mem3[148][25] ), .QN(n28511) );
  SDFFX1 \mem3_reg[148][24]  ( .D(n13644), .SI(\mem3[147][31] ), .SE(test_se), 
        .CLK(n1803), .Q(\mem3[148][24] ), .QN(n28512) );
  SDFFX1 \mem3_reg[147][31]  ( .D(n13643), .SI(\mem3[147][30] ), .SE(test_se), 
        .CLK(n1803), .Q(\mem3[147][31] ), .QN(n28513) );
  SDFFX1 \mem3_reg[147][30]  ( .D(n13642), .SI(\mem3[147][29] ), .SE(test_se), 
        .CLK(n1803), .Q(\mem3[147][30] ), .QN(n28514) );
  SDFFX1 \mem3_reg[147][29]  ( .D(n13641), .SI(\mem3[147][28] ), .SE(test_se), 
        .CLK(n1803), .Q(\mem3[147][29] ), .QN(n28515) );
  SDFFX1 \mem3_reg[147][28]  ( .D(n13640), .SI(\mem3[147][27] ), .SE(test_se), 
        .CLK(n1803), .Q(\mem3[147][28] ), .QN(n28516) );
  SDFFX1 \mem3_reg[147][27]  ( .D(n13639), .SI(\mem3[147][26] ), .SE(test_se), 
        .CLK(n1803), .Q(\mem3[147][27] ), .QN(n28517) );
  SDFFX1 \mem3_reg[147][26]  ( .D(n13638), .SI(\mem3[147][25] ), .SE(test_se), 
        .CLK(n1803), .Q(\mem3[147][26] ), .QN(n28518) );
  SDFFX1 \mem3_reg[147][25]  ( .D(n13637), .SI(\mem3[147][24] ), .SE(test_se), 
        .CLK(n1803), .Q(\mem3[147][25] ), .QN(n28519) );
  SDFFX1 \mem3_reg[147][24]  ( .D(n13636), .SI(\mem3[146][31] ), .SE(test_se), 
        .CLK(n1804), .Q(\mem3[147][24] ), .QN(n28520) );
  SDFFX1 \mem3_reg[146][31]  ( .D(n13635), .SI(\mem3[146][30] ), .SE(test_se), 
        .CLK(n1804), .Q(\mem3[146][31] ), .QN(n28521) );
  SDFFX1 \mem3_reg[146][30]  ( .D(n13634), .SI(\mem3[146][29] ), .SE(test_se), 
        .CLK(n1804), .Q(\mem3[146][30] ), .QN(n28522) );
  SDFFX1 \mem3_reg[146][29]  ( .D(n13633), .SI(\mem3[146][28] ), .SE(test_se), 
        .CLK(n1804), .Q(\mem3[146][29] ), .QN(n28523) );
  SDFFX1 \mem3_reg[146][28]  ( .D(n13632), .SI(\mem3[146][27] ), .SE(test_se), 
        .CLK(n1804), .Q(\mem3[146][28] ), .QN(n28524) );
  SDFFX1 \mem3_reg[146][27]  ( .D(n13631), .SI(\mem3[146][26] ), .SE(test_se), 
        .CLK(n1804), .Q(\mem3[146][27] ), .QN(n28525) );
  SDFFX1 \mem3_reg[146][26]  ( .D(n13630), .SI(\mem3[146][25] ), .SE(test_se), 
        .CLK(n1804), .Q(\mem3[146][26] ), .QN(n28526) );
  SDFFX1 \mem3_reg[146][25]  ( .D(n13629), .SI(\mem3[146][24] ), .SE(test_se), 
        .CLK(n1804), .Q(\mem3[146][25] ), .QN(n28527) );
  SDFFX1 \mem3_reg[146][24]  ( .D(n13628), .SI(\mem3[145][31] ), .SE(test_se), 
        .CLK(n1804), .Q(\mem3[146][24] ), .QN(n28528) );
  SDFFX1 \mem3_reg[145][31]  ( .D(n13627), .SI(\mem3[145][30] ), .SE(test_se), 
        .CLK(n1804), .Q(\mem3[145][31] ), .QN(n28529) );
  SDFFX1 \mem3_reg[145][30]  ( .D(n13626), .SI(\mem3[145][29] ), .SE(test_se), 
        .CLK(n1804), .Q(\mem3[145][30] ), .QN(n28530) );
  SDFFX1 \mem3_reg[145][29]  ( .D(n13625), .SI(\mem3[145][28] ), .SE(test_se), 
        .CLK(n1804), .Q(\mem3[145][29] ), .QN(n28531) );
  SDFFX1 \mem3_reg[145][28]  ( .D(n13624), .SI(\mem3[145][27] ), .SE(test_se), 
        .CLK(n1805), .Q(\mem3[145][28] ), .QN(n28532) );
  SDFFX1 \mem3_reg[145][27]  ( .D(n13623), .SI(\mem3[145][26] ), .SE(test_se), 
        .CLK(n1805), .Q(\mem3[145][27] ), .QN(n28533) );
  SDFFX1 \mem3_reg[145][26]  ( .D(n13622), .SI(\mem3[145][25] ), .SE(test_se), 
        .CLK(n1805), .Q(\mem3[145][26] ), .QN(n28534) );
  SDFFX1 \mem3_reg[145][25]  ( .D(n13621), .SI(\mem3[145][24] ), .SE(test_se), 
        .CLK(n1805), .Q(\mem3[145][25] ), .QN(n28535) );
  SDFFX1 \mem3_reg[145][24]  ( .D(n13620), .SI(\mem3[144][31] ), .SE(test_se), 
        .CLK(n1805), .Q(\mem3[145][24] ), .QN(n28536) );
  SDFFX1 \mem3_reg[144][31]  ( .D(n13619), .SI(\mem3[144][30] ), .SE(test_se), 
        .CLK(n1805), .Q(\mem3[144][31] ), .QN(n28537) );
  SDFFX1 \mem3_reg[144][30]  ( .D(n13618), .SI(\mem3[144][29] ), .SE(test_se), 
        .CLK(n1805), .Q(\mem3[144][30] ), .QN(n28538) );
  SDFFX1 \mem3_reg[144][29]  ( .D(n13617), .SI(\mem3[144][28] ), .SE(test_se), 
        .CLK(n1805), .Q(\mem3[144][29] ), .QN(n28539) );
  SDFFX1 \mem3_reg[144][28]  ( .D(n13616), .SI(\mem3[144][27] ), .SE(test_se), 
        .CLK(n1805), .Q(\mem3[144][28] ), .QN(n28540) );
  SDFFX1 \mem3_reg[144][27]  ( .D(n13615), .SI(\mem3[144][26] ), .SE(test_se), 
        .CLK(n1805), .Q(\mem3[144][27] ), .QN(n28541) );
  SDFFX1 \mem3_reg[144][26]  ( .D(n13614), .SI(\mem3[144][25] ), .SE(test_se), 
        .CLK(n1805), .Q(\mem3[144][26] ), .QN(n28542) );
  SDFFX1 \mem3_reg[144][25]  ( .D(n13613), .SI(\mem3[144][24] ), .SE(test_se), 
        .CLK(n1805), .Q(\mem3[144][25] ), .QN(n28543) );
  SDFFX1 \mem3_reg[144][24]  ( .D(n13612), .SI(\mem3[143][31] ), .SE(test_se), 
        .CLK(n1806), .Q(\mem3[144][24] ), .QN(n28544) );
  SDFFX1 \mem3_reg[143][31]  ( .D(n13611), .SI(\mem3[143][30] ), .SE(test_se), 
        .CLK(n1806), .Q(\mem3[143][31] ), .QN(n28545) );
  SDFFX1 \mem3_reg[143][30]  ( .D(n13610), .SI(\mem3[143][29] ), .SE(test_se), 
        .CLK(n1806), .Q(\mem3[143][30] ), .QN(n28546) );
  SDFFX1 \mem3_reg[143][29]  ( .D(n13609), .SI(\mem3[143][28] ), .SE(test_se), 
        .CLK(n1806), .Q(\mem3[143][29] ), .QN(n28547) );
  SDFFX1 \mem3_reg[143][28]  ( .D(n13608), .SI(\mem3[143][27] ), .SE(test_se), 
        .CLK(n1806), .Q(\mem3[143][28] ), .QN(n28548) );
  SDFFX1 \mem3_reg[143][27]  ( .D(n13607), .SI(\mem3[143][26] ), .SE(test_se), 
        .CLK(n1806), .Q(\mem3[143][27] ), .QN(n28549) );
  SDFFX1 \mem3_reg[143][26]  ( .D(n13606), .SI(\mem3[143][25] ), .SE(test_se), 
        .CLK(n1806), .Q(\mem3[143][26] ), .QN(n28550) );
  SDFFX1 \mem3_reg[143][25]  ( .D(n13605), .SI(\mem3[143][24] ), .SE(test_se), 
        .CLK(n1806), .Q(\mem3[143][25] ), .QN(n28551) );
  SDFFX1 \mem3_reg[143][24]  ( .D(n13604), .SI(\mem3[142][31] ), .SE(test_se), 
        .CLK(n1806), .Q(\mem3[143][24] ), .QN(n28552) );
  SDFFX1 \mem3_reg[142][31]  ( .D(n13603), .SI(\mem3[142][30] ), .SE(test_se), 
        .CLK(n1806), .Q(\mem3[142][31] ), .QN(n28553) );
  SDFFX1 \mem3_reg[142][30]  ( .D(n13602), .SI(\mem3[142][29] ), .SE(test_se), 
        .CLK(n1806), .Q(\mem3[142][30] ), .QN(n28554) );
  SDFFX1 \mem3_reg[142][29]  ( .D(n13601), .SI(\mem3[142][28] ), .SE(test_se), 
        .CLK(n1806), .Q(\mem3[142][29] ), .QN(n28555) );
  SDFFX1 \mem3_reg[142][28]  ( .D(n13600), .SI(\mem3[142][27] ), .SE(test_se), 
        .CLK(n1807), .Q(\mem3[142][28] ), .QN(n28556) );
  SDFFX1 \mem3_reg[142][27]  ( .D(n13599), .SI(\mem3[142][26] ), .SE(test_se), 
        .CLK(n1807), .Q(\mem3[142][27] ), .QN(n28557) );
  SDFFX1 \mem3_reg[142][26]  ( .D(n13598), .SI(\mem3[142][25] ), .SE(test_se), 
        .CLK(n1807), .Q(\mem3[142][26] ), .QN(n28558) );
  SDFFX1 \mem3_reg[142][25]  ( .D(n13597), .SI(\mem3[142][24] ), .SE(test_se), 
        .CLK(n1807), .Q(\mem3[142][25] ), .QN(n28559) );
  SDFFX1 \mem3_reg[142][24]  ( .D(n13596), .SI(\mem3[141][31] ), .SE(test_se), 
        .CLK(n1807), .Q(\mem3[142][24] ), .QN(n28560) );
  SDFFX1 \mem3_reg[141][31]  ( .D(n13595), .SI(\mem3[141][30] ), .SE(test_se), 
        .CLK(n1807), .Q(\mem3[141][31] ), .QN(n28561) );
  SDFFX1 \mem3_reg[141][30]  ( .D(n13594), .SI(\mem3[141][29] ), .SE(test_se), 
        .CLK(n1807), .Q(\mem3[141][30] ), .QN(n28562) );
  SDFFX1 \mem3_reg[141][29]  ( .D(n13593), .SI(\mem3[141][28] ), .SE(test_se), 
        .CLK(n1807), .Q(\mem3[141][29] ), .QN(n28563) );
  SDFFX1 \mem3_reg[141][28]  ( .D(n13592), .SI(\mem3[141][27] ), .SE(test_se), 
        .CLK(n1807), .Q(\mem3[141][28] ), .QN(n28564) );
  SDFFX1 \mem3_reg[141][27]  ( .D(n13591), .SI(\mem3[141][26] ), .SE(test_se), 
        .CLK(n1807), .Q(\mem3[141][27] ), .QN(n28565) );
  SDFFX1 \mem3_reg[141][26]  ( .D(n13590), .SI(\mem3[141][25] ), .SE(test_se), 
        .CLK(n1807), .Q(\mem3[141][26] ), .QN(n28566) );
  SDFFX1 \mem3_reg[141][25]  ( .D(n13589), .SI(\mem3[141][24] ), .SE(test_se), 
        .CLK(n1807), .Q(\mem3[141][25] ), .QN(n28567) );
  SDFFX1 \mem3_reg[141][24]  ( .D(n13588), .SI(\mem3[140][31] ), .SE(test_se), 
        .CLK(n1808), .Q(\mem3[141][24] ), .QN(n28568) );
  SDFFX1 \mem3_reg[140][31]  ( .D(n13587), .SI(\mem3[140][30] ), .SE(test_se), 
        .CLK(n1808), .Q(\mem3[140][31] ), .QN(n28569) );
  SDFFX1 \mem3_reg[140][30]  ( .D(n13586), .SI(\mem3[140][29] ), .SE(test_se), 
        .CLK(n1808), .Q(\mem3[140][30] ), .QN(n28570) );
  SDFFX1 \mem3_reg[140][29]  ( .D(n13585), .SI(\mem3[140][28] ), .SE(test_se), 
        .CLK(n1808), .Q(\mem3[140][29] ), .QN(n28571) );
  SDFFX1 \mem3_reg[140][28]  ( .D(n13584), .SI(\mem3[140][27] ), .SE(test_se), 
        .CLK(n1808), .Q(\mem3[140][28] ), .QN(n28572) );
  SDFFX1 \mem3_reg[140][27]  ( .D(n13583), .SI(\mem3[140][26] ), .SE(test_se), 
        .CLK(n1808), .Q(\mem3[140][27] ), .QN(n28573) );
  SDFFX1 \mem3_reg[140][26]  ( .D(n13582), .SI(\mem3[140][25] ), .SE(test_se), 
        .CLK(n1808), .Q(\mem3[140][26] ), .QN(n28574) );
  SDFFX1 \mem3_reg[140][25]  ( .D(n13581), .SI(\mem3[140][24] ), .SE(test_se), 
        .CLK(n1808), .Q(\mem3[140][25] ), .QN(n28575) );
  SDFFX1 \mem3_reg[140][24]  ( .D(n13580), .SI(\mem3[139][31] ), .SE(test_se), 
        .CLK(n1808), .Q(\mem3[140][24] ), .QN(n28576) );
  SDFFX1 \mem3_reg[139][31]  ( .D(n13579), .SI(\mem3[139][30] ), .SE(test_se), 
        .CLK(n1808), .Q(\mem3[139][31] ), .QN(n28577) );
  SDFFX1 \mem3_reg[139][30]  ( .D(n13578), .SI(\mem3[139][29] ), .SE(test_se), 
        .CLK(n1808), .Q(\mem3[139][30] ), .QN(n28578) );
  SDFFX1 \mem3_reg[139][29]  ( .D(n13577), .SI(\mem3[139][28] ), .SE(test_se), 
        .CLK(n1808), .Q(\mem3[139][29] ), .QN(n28579) );
  SDFFX1 \mem3_reg[139][28]  ( .D(n13576), .SI(\mem3[139][27] ), .SE(test_se), 
        .CLK(n1809), .Q(\mem3[139][28] ), .QN(n28580) );
  SDFFX1 \mem3_reg[139][27]  ( .D(n13575), .SI(\mem3[139][26] ), .SE(test_se), 
        .CLK(n1809), .Q(\mem3[139][27] ), .QN(n28581) );
  SDFFX1 \mem3_reg[139][26]  ( .D(n13574), .SI(\mem3[139][25] ), .SE(test_se), 
        .CLK(n1809), .Q(\mem3[139][26] ), .QN(n28582) );
  SDFFX1 \mem3_reg[139][25]  ( .D(n13573), .SI(\mem3[139][24] ), .SE(test_se), 
        .CLK(n1809), .Q(\mem3[139][25] ), .QN(n28583) );
  SDFFX1 \mem3_reg[139][24]  ( .D(n13572), .SI(\mem3[138][31] ), .SE(test_se), 
        .CLK(n1809), .Q(\mem3[139][24] ), .QN(n28584) );
  SDFFX1 \mem3_reg[138][31]  ( .D(n13571), .SI(\mem3[138][30] ), .SE(test_se), 
        .CLK(n1809), .Q(\mem3[138][31] ), .QN(n28585) );
  SDFFX1 \mem3_reg[138][30]  ( .D(n13570), .SI(\mem3[138][29] ), .SE(test_se), 
        .CLK(n1809), .Q(\mem3[138][30] ), .QN(n28586) );
  SDFFX1 \mem3_reg[138][29]  ( .D(n13569), .SI(\mem3[138][28] ), .SE(test_se), 
        .CLK(n1809), .Q(\mem3[138][29] ), .QN(n28587) );
  SDFFX1 \mem3_reg[138][28]  ( .D(n13568), .SI(\mem3[138][27] ), .SE(test_se), 
        .CLK(n1809), .Q(\mem3[138][28] ), .QN(n28588) );
  SDFFX1 \mem3_reg[138][27]  ( .D(n13567), .SI(\mem3[138][26] ), .SE(test_se), 
        .CLK(n1809), .Q(\mem3[138][27] ), .QN(n28589) );
  SDFFX1 \mem3_reg[138][26]  ( .D(n13566), .SI(\mem3[138][25] ), .SE(test_se), 
        .CLK(n1809), .Q(\mem3[138][26] ), .QN(n28590) );
  SDFFX1 \mem3_reg[138][25]  ( .D(n13565), .SI(\mem3[138][24] ), .SE(test_se), 
        .CLK(n1809), .Q(\mem3[138][25] ), .QN(n28591) );
  SDFFX1 \mem3_reg[138][24]  ( .D(n13564), .SI(\mem3[137][31] ), .SE(test_se), 
        .CLK(n1810), .Q(\mem3[138][24] ), .QN(n28592) );
  SDFFX1 \mem3_reg[137][31]  ( .D(n13563), .SI(\mem3[137][30] ), .SE(test_se), 
        .CLK(n1810), .Q(\mem3[137][31] ), .QN(n28593) );
  SDFFX1 \mem3_reg[137][30]  ( .D(n13562), .SI(\mem3[137][29] ), .SE(test_se), 
        .CLK(n1810), .Q(\mem3[137][30] ), .QN(n28594) );
  SDFFX1 \mem3_reg[137][29]  ( .D(n13561), .SI(\mem3[137][28] ), .SE(test_se), 
        .CLK(n1810), .Q(\mem3[137][29] ), .QN(n28595) );
  SDFFX1 \mem3_reg[137][28]  ( .D(n13560), .SI(\mem3[137][27] ), .SE(test_se), 
        .CLK(n1810), .Q(\mem3[137][28] ), .QN(n28596) );
  SDFFX1 \mem3_reg[137][27]  ( .D(n13559), .SI(\mem3[137][26] ), .SE(test_se), 
        .CLK(n1810), .Q(\mem3[137][27] ), .QN(n28597) );
  SDFFX1 \mem3_reg[137][26]  ( .D(n13558), .SI(\mem3[137][25] ), .SE(test_se), 
        .CLK(n1810), .Q(\mem3[137][26] ), .QN(n28598) );
  SDFFX1 \mem3_reg[137][25]  ( .D(n13557), .SI(\mem3[137][24] ), .SE(test_se), 
        .CLK(n1810), .Q(\mem3[137][25] ), .QN(n28599) );
  SDFFX1 \mem3_reg[137][24]  ( .D(n13556), .SI(\mem3[136][31] ), .SE(test_se), 
        .CLK(n1810), .Q(\mem3[137][24] ), .QN(n28600) );
  SDFFX1 \mem3_reg[136][31]  ( .D(n13555), .SI(\mem3[136][30] ), .SE(test_se), 
        .CLK(n1810), .Q(\mem3[136][31] ), .QN(n28601) );
  SDFFX1 \mem3_reg[136][30]  ( .D(n13554), .SI(\mem3[136][29] ), .SE(test_se), 
        .CLK(n1810), .Q(\mem3[136][30] ), .QN(n28602) );
  SDFFX1 \mem3_reg[136][29]  ( .D(n13553), .SI(\mem3[136][28] ), .SE(test_se), 
        .CLK(n1810), .Q(\mem3[136][29] ), .QN(n28603) );
  SDFFX1 \mem3_reg[136][28]  ( .D(n13552), .SI(\mem3[136][27] ), .SE(test_se), 
        .CLK(n1811), .Q(\mem3[136][28] ), .QN(n28604) );
  SDFFX1 \mem3_reg[136][27]  ( .D(n13551), .SI(\mem3[136][26] ), .SE(test_se), 
        .CLK(n1811), .Q(\mem3[136][27] ), .QN(n28605) );
  SDFFX1 \mem3_reg[136][26]  ( .D(n13550), .SI(\mem3[136][25] ), .SE(test_se), 
        .CLK(n1811), .Q(\mem3[136][26] ), .QN(n28606) );
  SDFFX1 \mem3_reg[136][25]  ( .D(n13549), .SI(\mem3[136][24] ), .SE(test_se), 
        .CLK(n1811), .Q(\mem3[136][25] ), .QN(n28607) );
  SDFFX1 \mem3_reg[136][24]  ( .D(n13548), .SI(\mem3[135][31] ), .SE(test_se), 
        .CLK(n1811), .Q(\mem3[136][24] ), .QN(n28608) );
  SDFFX1 \mem3_reg[135][31]  ( .D(n13547), .SI(\mem3[135][30] ), .SE(test_se), 
        .CLK(n1811), .Q(\mem3[135][31] ), .QN(n28609) );
  SDFFX1 \mem3_reg[135][30]  ( .D(n13546), .SI(\mem3[135][29] ), .SE(test_se), 
        .CLK(n1811), .Q(\mem3[135][30] ), .QN(n28610) );
  SDFFX1 \mem3_reg[135][29]  ( .D(n13545), .SI(\mem3[135][28] ), .SE(test_se), 
        .CLK(n1811), .Q(\mem3[135][29] ), .QN(n28611) );
  SDFFX1 \mem3_reg[135][28]  ( .D(n13544), .SI(\mem3[135][27] ), .SE(test_se), 
        .CLK(n1811), .Q(\mem3[135][28] ), .QN(n28612) );
  SDFFX1 \mem3_reg[135][27]  ( .D(n13543), .SI(\mem3[135][26] ), .SE(test_se), 
        .CLK(n1811), .Q(\mem3[135][27] ), .QN(n28613) );
  SDFFX1 \mem3_reg[135][26]  ( .D(n13542), .SI(\mem3[135][25] ), .SE(test_se), 
        .CLK(n1811), .Q(\mem3[135][26] ), .QN(n28614) );
  SDFFX1 \mem3_reg[135][25]  ( .D(n13541), .SI(\mem3[135][24] ), .SE(test_se), 
        .CLK(n1811), .Q(\mem3[135][25] ), .QN(n28615) );
  SDFFX1 \mem3_reg[135][24]  ( .D(n13540), .SI(\mem3[134][31] ), .SE(test_se), 
        .CLK(n1812), .Q(\mem3[135][24] ), .QN(n28616) );
  SDFFX1 \mem3_reg[134][31]  ( .D(n13539), .SI(\mem3[134][30] ), .SE(test_se), 
        .CLK(n1812), .Q(\mem3[134][31] ), .QN(n28617) );
  SDFFX1 \mem3_reg[134][30]  ( .D(n13538), .SI(\mem3[134][29] ), .SE(test_se), 
        .CLK(n1812), .Q(\mem3[134][30] ), .QN(n28618) );
  SDFFX1 \mem3_reg[134][29]  ( .D(n13537), .SI(\mem3[134][28] ), .SE(test_se), 
        .CLK(n1812), .Q(\mem3[134][29] ), .QN(n28619) );
  SDFFX1 \mem3_reg[134][28]  ( .D(n13536), .SI(\mem3[134][27] ), .SE(test_se), 
        .CLK(n1812), .Q(\mem3[134][28] ), .QN(n28620) );
  SDFFX1 \mem3_reg[134][27]  ( .D(n13535), .SI(\mem3[134][26] ), .SE(test_se), 
        .CLK(n1812), .Q(\mem3[134][27] ), .QN(n28621) );
  SDFFX1 \mem3_reg[134][26]  ( .D(n13534), .SI(\mem3[134][25] ), .SE(test_se), 
        .CLK(n1812), .Q(\mem3[134][26] ), .QN(n28622) );
  SDFFX1 \mem3_reg[134][25]  ( .D(n13533), .SI(\mem3[134][24] ), .SE(test_se), 
        .CLK(n1812), .Q(\mem3[134][25] ), .QN(n28623) );
  SDFFX1 \mem3_reg[134][24]  ( .D(n13532), .SI(\mem3[133][31] ), .SE(test_se), 
        .CLK(n1812), .Q(\mem3[134][24] ), .QN(n28624) );
  SDFFX1 \mem3_reg[133][31]  ( .D(n13531), .SI(\mem3[133][30] ), .SE(test_se), 
        .CLK(n1812), .Q(\mem3[133][31] ), .QN(n28625) );
  SDFFX1 \mem3_reg[133][30]  ( .D(n13530), .SI(\mem3[133][29] ), .SE(test_se), 
        .CLK(n1812), .Q(\mem3[133][30] ), .QN(n28626) );
  SDFFX1 \mem3_reg[133][29]  ( .D(n13529), .SI(\mem3[133][28] ), .SE(test_se), 
        .CLK(n1812), .Q(\mem3[133][29] ), .QN(n28627) );
  SDFFX1 \mem3_reg[133][28]  ( .D(n13528), .SI(\mem3[133][27] ), .SE(test_se), 
        .CLK(n1813), .Q(\mem3[133][28] ), .QN(n28628) );
  SDFFX1 \mem3_reg[133][27]  ( .D(n13527), .SI(\mem3[133][26] ), .SE(test_se), 
        .CLK(n1813), .Q(\mem3[133][27] ), .QN(n28629) );
  SDFFX1 \mem3_reg[133][26]  ( .D(n13526), .SI(\mem3[133][25] ), .SE(test_se), 
        .CLK(n1813), .Q(\mem3[133][26] ), .QN(n28630) );
  SDFFX1 \mem3_reg[133][25]  ( .D(n13525), .SI(\mem3[133][24] ), .SE(test_se), 
        .CLK(n1813), .Q(\mem3[133][25] ), .QN(n28631) );
  SDFFX1 \mem3_reg[133][24]  ( .D(n13524), .SI(\mem3[132][31] ), .SE(test_se), 
        .CLK(n1813), .Q(\mem3[133][24] ), .QN(n28632) );
  SDFFX1 \mem3_reg[132][31]  ( .D(n13523), .SI(\mem3[132][30] ), .SE(test_se), 
        .CLK(n1813), .Q(\mem3[132][31] ), .QN(n28633) );
  SDFFX1 \mem3_reg[132][30]  ( .D(n13522), .SI(\mem3[132][29] ), .SE(test_se), 
        .CLK(n1813), .Q(\mem3[132][30] ), .QN(n28634) );
  SDFFX1 \mem3_reg[132][29]  ( .D(n13521), .SI(\mem3[132][28] ), .SE(test_se), 
        .CLK(n1813), .Q(\mem3[132][29] ), .QN(n28635) );
  SDFFX1 \mem3_reg[132][28]  ( .D(n13520), .SI(\mem3[132][27] ), .SE(test_se), 
        .CLK(n1813), .Q(\mem3[132][28] ), .QN(n28636) );
  SDFFX1 \mem3_reg[132][27]  ( .D(n13519), .SI(\mem3[132][26] ), .SE(test_se), 
        .CLK(n1813), .Q(\mem3[132][27] ), .QN(n28637) );
  SDFFX1 \mem3_reg[132][26]  ( .D(n13518), .SI(\mem3[132][25] ), .SE(test_se), 
        .CLK(n1813), .Q(\mem3[132][26] ), .QN(n28638) );
  SDFFX1 \mem3_reg[132][25]  ( .D(n13517), .SI(\mem3[132][24] ), .SE(test_se), 
        .CLK(n1813), .Q(\mem3[132][25] ), .QN(n28639) );
  SDFFX1 \mem3_reg[132][24]  ( .D(n13516), .SI(\mem3[131][31] ), .SE(test_se), 
        .CLK(n1814), .Q(\mem3[132][24] ), .QN(n28640) );
  SDFFX1 \mem3_reg[131][31]  ( .D(n13515), .SI(\mem3[131][30] ), .SE(test_se), 
        .CLK(n1814), .Q(\mem3[131][31] ), .QN(n28641) );
  SDFFX1 \mem3_reg[131][30]  ( .D(n13514), .SI(\mem3[131][29] ), .SE(test_se), 
        .CLK(n1814), .Q(\mem3[131][30] ), .QN(n28642) );
  SDFFX1 \mem3_reg[131][29]  ( .D(n13513), .SI(\mem3[131][28] ), .SE(test_se), 
        .CLK(n1814), .Q(\mem3[131][29] ), .QN(n28643) );
  SDFFX1 \mem3_reg[131][28]  ( .D(n13512), .SI(\mem3[131][27] ), .SE(test_se), 
        .CLK(n1814), .Q(\mem3[131][28] ), .QN(n28644) );
  SDFFX1 \mem3_reg[131][27]  ( .D(n13511), .SI(\mem3[131][26] ), .SE(test_se), 
        .CLK(n1814), .Q(\mem3[131][27] ), .QN(n28645) );
  SDFFX1 \mem3_reg[131][26]  ( .D(n13510), .SI(\mem3[131][25] ), .SE(test_se), 
        .CLK(n1814), .Q(\mem3[131][26] ), .QN(n28646) );
  SDFFX1 \mem3_reg[131][25]  ( .D(n13509), .SI(\mem3[131][24] ), .SE(test_se), 
        .CLK(n1814), .Q(\mem3[131][25] ), .QN(n28647) );
  SDFFX1 \mem3_reg[131][24]  ( .D(n13508), .SI(\mem3[130][31] ), .SE(test_se), 
        .CLK(n1814), .Q(\mem3[131][24] ), .QN(n28648) );
  SDFFX1 \mem3_reg[130][31]  ( .D(n13507), .SI(\mem3[130][30] ), .SE(test_se), 
        .CLK(n1814), .Q(\mem3[130][31] ), .QN(n28649) );
  SDFFX1 \mem3_reg[130][30]  ( .D(n13506), .SI(\mem3[130][29] ), .SE(test_se), 
        .CLK(n1814), .Q(\mem3[130][30] ), .QN(n28650) );
  SDFFX1 \mem3_reg[130][29]  ( .D(n13505), .SI(\mem3[130][28] ), .SE(test_se), 
        .CLK(n1814), .Q(\mem3[130][29] ), .QN(n28651) );
  SDFFX1 \mem3_reg[130][28]  ( .D(n13504), .SI(\mem3[130][27] ), .SE(test_se), 
        .CLK(n1815), .Q(\mem3[130][28] ), .QN(n28652) );
  SDFFX1 \mem3_reg[130][27]  ( .D(n13503), .SI(\mem3[130][26] ), .SE(test_se), 
        .CLK(n1815), .Q(\mem3[130][27] ), .QN(n28653) );
  SDFFX1 \mem3_reg[130][26]  ( .D(n13502), .SI(\mem3[130][25] ), .SE(test_se), 
        .CLK(n1815), .Q(\mem3[130][26] ), .QN(n28654) );
  SDFFX1 \mem3_reg[130][25]  ( .D(n13501), .SI(\mem3[130][24] ), .SE(test_se), 
        .CLK(n1815), .Q(\mem3[130][25] ), .QN(n28655) );
  SDFFX1 \mem3_reg[130][24]  ( .D(n13500), .SI(\mem3[129][31] ), .SE(test_se), 
        .CLK(n1815), .Q(\mem3[130][24] ), .QN(n28656) );
  SDFFX1 \mem3_reg[129][31]  ( .D(n13499), .SI(\mem3[129][30] ), .SE(test_se), 
        .CLK(n1815), .Q(\mem3[129][31] ), .QN(n28657) );
  SDFFX1 \mem3_reg[129][30]  ( .D(n13498), .SI(\mem3[129][29] ), .SE(test_se), 
        .CLK(n1815), .Q(\mem3[129][30] ), .QN(n28658) );
  SDFFX1 \mem3_reg[129][29]  ( .D(n13497), .SI(\mem3[129][28] ), .SE(test_se), 
        .CLK(n1815), .Q(\mem3[129][29] ), .QN(n28659) );
  SDFFX1 \mem3_reg[129][28]  ( .D(n13496), .SI(\mem3[129][27] ), .SE(test_se), 
        .CLK(n1815), .Q(\mem3[129][28] ), .QN(n28660) );
  SDFFX1 \mem3_reg[129][27]  ( .D(n13495), .SI(\mem3[129][26] ), .SE(test_se), 
        .CLK(n1815), .Q(\mem3[129][27] ), .QN(n28661) );
  SDFFX1 \mem3_reg[129][26]  ( .D(n13494), .SI(\mem3[129][25] ), .SE(test_se), 
        .CLK(n1815), .Q(\mem3[129][26] ), .QN(n28662) );
  SDFFX1 \mem3_reg[129][25]  ( .D(n13493), .SI(\mem3[129][24] ), .SE(test_se), 
        .CLK(n1815), .Q(\mem3[129][25] ), .QN(n28663) );
  SDFFX1 \mem3_reg[129][24]  ( .D(n13492), .SI(\mem3[128][31] ), .SE(test_se), 
        .CLK(n1816), .Q(\mem3[129][24] ), .QN(n28664) );
  SDFFX1 \mem3_reg[128][31]  ( .D(n13491), .SI(\mem3[128][30] ), .SE(test_se), 
        .CLK(n1816), .Q(\mem3[128][31] ), .QN(n28665) );
  SDFFX1 \mem3_reg[128][30]  ( .D(n13490), .SI(\mem3[128][29] ), .SE(test_se), 
        .CLK(n1816), .Q(\mem3[128][30] ), .QN(n28666) );
  SDFFX1 \mem3_reg[128][29]  ( .D(n13489), .SI(\mem3[128][28] ), .SE(test_se), 
        .CLK(n1816), .Q(\mem3[128][29] ), .QN(n28667) );
  SDFFX1 \mem3_reg[128][28]  ( .D(n13488), .SI(\mem3[128][27] ), .SE(test_se), 
        .CLK(n1816), .Q(\mem3[128][28] ), .QN(n28668) );
  SDFFX1 \mem3_reg[128][27]  ( .D(n13487), .SI(\mem3[128][26] ), .SE(test_se), 
        .CLK(n1816), .Q(\mem3[128][27] ), .QN(n28669) );
  SDFFX1 \mem3_reg[128][26]  ( .D(n13486), .SI(\mem3[128][25] ), .SE(test_se), 
        .CLK(n1816), .Q(\mem3[128][26] ), .QN(n28670) );
  SDFFX1 \mem3_reg[128][25]  ( .D(n13485), .SI(\mem3[128][24] ), .SE(test_se), 
        .CLK(n1816), .Q(\mem3[128][25] ), .QN(n28671) );
  SDFFX1 \mem3_reg[128][24]  ( .D(n13484), .SI(\mem3[127][31] ), .SE(test_se), 
        .CLK(n1816), .Q(\mem3[128][24] ), .QN(n28672) );
  SDFFX1 \mem3_reg[127][31]  ( .D(n13483), .SI(\mem3[127][30] ), .SE(test_se), 
        .CLK(n1816), .Q(\mem3[127][31] ), .QN(n28673) );
  SDFFX1 \mem3_reg[127][30]  ( .D(n13482), .SI(\mem3[127][29] ), .SE(test_se), 
        .CLK(n1816), .Q(\mem3[127][30] ), .QN(n28674) );
  SDFFX1 \mem3_reg[127][29]  ( .D(n13481), .SI(\mem3[127][28] ), .SE(test_se), 
        .CLK(n1816), .Q(\mem3[127][29] ), .QN(n28675) );
  SDFFX1 \mem3_reg[127][28]  ( .D(n13480), .SI(\mem3[127][27] ), .SE(test_se), 
        .CLK(n1817), .Q(\mem3[127][28] ), .QN(n28676) );
  SDFFX1 \mem3_reg[127][27]  ( .D(n13479), .SI(\mem3[127][26] ), .SE(test_se), 
        .CLK(n1817), .Q(\mem3[127][27] ), .QN(n28677) );
  SDFFX1 \mem3_reg[127][26]  ( .D(n13478), .SI(\mem3[127][25] ), .SE(test_se), 
        .CLK(n1817), .Q(\mem3[127][26] ), .QN(n28678) );
  SDFFX1 \mem3_reg[127][25]  ( .D(n13477), .SI(\mem3[127][24] ), .SE(test_se), 
        .CLK(n1817), .Q(\mem3[127][25] ), .QN(n28679) );
  SDFFX1 \mem3_reg[127][24]  ( .D(n13476), .SI(\mem3[126][31] ), .SE(test_se), 
        .CLK(n1817), .Q(\mem3[127][24] ), .QN(n28680) );
  SDFFX1 \mem3_reg[126][31]  ( .D(n13475), .SI(\mem3[126][30] ), .SE(test_se), 
        .CLK(n1817), .Q(\mem3[126][31] ), .QN(n28681) );
  SDFFX1 \mem3_reg[126][30]  ( .D(n13474), .SI(\mem3[126][29] ), .SE(test_se), 
        .CLK(n1817), .Q(\mem3[126][30] ), .QN(n28682) );
  SDFFX1 \mem3_reg[126][29]  ( .D(n13473), .SI(\mem3[126][28] ), .SE(test_se), 
        .CLK(n1817), .Q(\mem3[126][29] ), .QN(n28683) );
  SDFFX1 \mem3_reg[126][28]  ( .D(n13472), .SI(\mem3[126][27] ), .SE(test_se), 
        .CLK(n1817), .Q(\mem3[126][28] ), .QN(n28684) );
  SDFFX1 \mem3_reg[126][27]  ( .D(n13471), .SI(\mem3[126][26] ), .SE(test_se), 
        .CLK(n1817), .Q(\mem3[126][27] ), .QN(n28685) );
  SDFFX1 \mem3_reg[126][26]  ( .D(n13470), .SI(\mem3[126][25] ), .SE(test_se), 
        .CLK(n1817), .Q(\mem3[126][26] ), .QN(n28686) );
  SDFFX1 \mem3_reg[126][25]  ( .D(n13469), .SI(\mem3[126][24] ), .SE(test_se), 
        .CLK(n1817), .Q(\mem3[126][25] ), .QN(n28687) );
  SDFFX1 \mem3_reg[126][24]  ( .D(n13468), .SI(\mem3[125][31] ), .SE(test_se), 
        .CLK(n1818), .Q(\mem3[126][24] ), .QN(n28688) );
  SDFFX1 \mem3_reg[125][31]  ( .D(n13467), .SI(\mem3[125][30] ), .SE(test_se), 
        .CLK(n1818), .Q(\mem3[125][31] ), .QN(n28689) );
  SDFFX1 \mem3_reg[125][30]  ( .D(n13466), .SI(\mem3[125][29] ), .SE(test_se), 
        .CLK(n1818), .Q(\mem3[125][30] ), .QN(n28690) );
  SDFFX1 \mem3_reg[125][29]  ( .D(n13465), .SI(\mem3[125][28] ), .SE(test_se), 
        .CLK(n1818), .Q(\mem3[125][29] ), .QN(n28691) );
  SDFFX1 \mem3_reg[125][28]  ( .D(n13464), .SI(\mem3[125][27] ), .SE(test_se), 
        .CLK(n1818), .Q(\mem3[125][28] ), .QN(n28692) );
  SDFFX1 \mem3_reg[125][27]  ( .D(n13463), .SI(\mem3[125][26] ), .SE(test_se), 
        .CLK(n1818), .Q(\mem3[125][27] ), .QN(n28693) );
  SDFFX1 \mem3_reg[125][26]  ( .D(n13462), .SI(\mem3[125][25] ), .SE(test_se), 
        .CLK(n1818), .Q(\mem3[125][26] ), .QN(n28694) );
  SDFFX1 \mem3_reg[125][25]  ( .D(n13461), .SI(\mem3[125][24] ), .SE(test_se), 
        .CLK(n1818), .Q(\mem3[125][25] ), .QN(n28695) );
  SDFFX1 \mem3_reg[125][24]  ( .D(n13460), .SI(\mem3[124][31] ), .SE(test_se), 
        .CLK(n1818), .Q(\mem3[125][24] ), .QN(n28696) );
  SDFFX1 \mem3_reg[124][31]  ( .D(n13459), .SI(\mem3[124][30] ), .SE(test_se), 
        .CLK(n1818), .Q(\mem3[124][31] ), .QN(n28697) );
  SDFFX1 \mem3_reg[124][30]  ( .D(n13458), .SI(\mem3[124][29] ), .SE(test_se), 
        .CLK(n1818), .Q(\mem3[124][30] ), .QN(n28698) );
  SDFFX1 \mem3_reg[124][29]  ( .D(n13457), .SI(\mem3[124][28] ), .SE(test_se), 
        .CLK(n1818), .Q(\mem3[124][29] ), .QN(n28699) );
  SDFFX1 \mem3_reg[124][28]  ( .D(n13456), .SI(\mem3[124][27] ), .SE(test_se), 
        .CLK(n1819), .Q(\mem3[124][28] ), .QN(n28700) );
  SDFFX1 \mem3_reg[124][27]  ( .D(n13455), .SI(\mem3[124][26] ), .SE(test_se), 
        .CLK(n1819), .Q(\mem3[124][27] ), .QN(n28701) );
  SDFFX1 \mem3_reg[124][26]  ( .D(n13454), .SI(\mem3[124][25] ), .SE(test_se), 
        .CLK(n1819), .Q(\mem3[124][26] ), .QN(n28702) );
  SDFFX1 \mem3_reg[124][25]  ( .D(n13453), .SI(\mem3[124][24] ), .SE(test_se), 
        .CLK(n1819), .Q(\mem3[124][25] ), .QN(n28703) );
  SDFFX1 \mem3_reg[124][24]  ( .D(n13452), .SI(\mem3[123][31] ), .SE(test_se), 
        .CLK(n1819), .Q(\mem3[124][24] ), .QN(n28704) );
  SDFFX1 \mem3_reg[123][31]  ( .D(n13451), .SI(\mem3[123][30] ), .SE(test_se), 
        .CLK(n1819), .Q(\mem3[123][31] ), .QN(n28705) );
  SDFFX1 \mem3_reg[123][30]  ( .D(n13450), .SI(\mem3[123][29] ), .SE(test_se), 
        .CLK(n1819), .Q(\mem3[123][30] ), .QN(n28706) );
  SDFFX1 \mem3_reg[123][29]  ( .D(n13449), .SI(\mem3[123][28] ), .SE(test_se), 
        .CLK(n1819), .Q(\mem3[123][29] ), .QN(n28707) );
  SDFFX1 \mem3_reg[123][28]  ( .D(n13448), .SI(\mem3[123][27] ), .SE(test_se), 
        .CLK(n1819), .Q(\mem3[123][28] ), .QN(n28708) );
  SDFFX1 \mem3_reg[123][27]  ( .D(n13447), .SI(\mem3[123][26] ), .SE(test_se), 
        .CLK(n1819), .Q(\mem3[123][27] ), .QN(n28709) );
  SDFFX1 \mem3_reg[123][26]  ( .D(n13446), .SI(\mem3[123][25] ), .SE(test_se), 
        .CLK(n1819), .Q(\mem3[123][26] ), .QN(n28710) );
  SDFFX1 \mem3_reg[123][25]  ( .D(n13445), .SI(\mem3[123][24] ), .SE(test_se), 
        .CLK(n1819), .Q(\mem3[123][25] ), .QN(n28711) );
  SDFFX1 \mem3_reg[123][24]  ( .D(n13444), .SI(\mem3[122][31] ), .SE(test_se), 
        .CLK(n1820), .Q(\mem3[123][24] ), .QN(n28712) );
  SDFFX1 \mem3_reg[122][31]  ( .D(n13443), .SI(\mem3[122][30] ), .SE(test_se), 
        .CLK(n1820), .Q(\mem3[122][31] ), .QN(n28713) );
  SDFFX1 \mem3_reg[122][30]  ( .D(n13442), .SI(\mem3[122][29] ), .SE(test_se), 
        .CLK(n1820), .Q(\mem3[122][30] ), .QN(n28714) );
  SDFFX1 \mem3_reg[122][29]  ( .D(n13441), .SI(\mem3[122][28] ), .SE(test_se), 
        .CLK(n1820), .Q(\mem3[122][29] ), .QN(n28715) );
  SDFFX1 \mem3_reg[122][28]  ( .D(n13440), .SI(\mem3[122][27] ), .SE(test_se), 
        .CLK(n1820), .Q(\mem3[122][28] ), .QN(n28716) );
  SDFFX1 \mem3_reg[122][27]  ( .D(n13439), .SI(\mem3[122][26] ), .SE(test_se), 
        .CLK(n1820), .Q(\mem3[122][27] ), .QN(n28717) );
  SDFFX1 \mem3_reg[122][26]  ( .D(n13438), .SI(\mem3[122][25] ), .SE(test_se), 
        .CLK(n1820), .Q(\mem3[122][26] ), .QN(n28718) );
  SDFFX1 \mem3_reg[122][25]  ( .D(n13437), .SI(\mem3[122][24] ), .SE(test_se), 
        .CLK(n1820), .Q(\mem3[122][25] ), .QN(n28719) );
  SDFFX1 \mem3_reg[122][24]  ( .D(n13436), .SI(\mem3[121][31] ), .SE(test_se), 
        .CLK(n1820), .Q(\mem3[122][24] ), .QN(n28720) );
  SDFFX1 \mem3_reg[121][31]  ( .D(n13435), .SI(\mem3[121][30] ), .SE(test_se), 
        .CLK(n1820), .Q(\mem3[121][31] ), .QN(n28721) );
  SDFFX1 \mem3_reg[121][30]  ( .D(n13434), .SI(\mem3[121][29] ), .SE(test_se), 
        .CLK(n1820), .Q(\mem3[121][30] ), .QN(n28722) );
  SDFFX1 \mem3_reg[121][29]  ( .D(n13433), .SI(\mem3[121][28] ), .SE(test_se), 
        .CLK(n1820), .Q(\mem3[121][29] ), .QN(n28723) );
  SDFFX1 \mem3_reg[121][28]  ( .D(n13432), .SI(\mem3[121][27] ), .SE(test_se), 
        .CLK(n1821), .Q(\mem3[121][28] ), .QN(n28724) );
  SDFFX1 \mem3_reg[121][27]  ( .D(n13431), .SI(\mem3[121][26] ), .SE(test_se), 
        .CLK(n1821), .Q(\mem3[121][27] ), .QN(n28725) );
  SDFFX1 \mem3_reg[121][26]  ( .D(n13430), .SI(\mem3[121][25] ), .SE(test_se), 
        .CLK(n1821), .Q(\mem3[121][26] ), .QN(n28726) );
  SDFFX1 \mem3_reg[121][25]  ( .D(n13429), .SI(\mem3[121][24] ), .SE(test_se), 
        .CLK(n1821), .Q(\mem3[121][25] ), .QN(n28727) );
  SDFFX1 \mem3_reg[121][24]  ( .D(n13428), .SI(\mem3[120][31] ), .SE(test_se), 
        .CLK(n1821), .Q(\mem3[121][24] ), .QN(n28728) );
  SDFFX1 \mem3_reg[120][31]  ( .D(n13427), .SI(\mem3[120][30] ), .SE(test_se), 
        .CLK(n1821), .Q(\mem3[120][31] ), .QN(n28729) );
  SDFFX1 \mem3_reg[120][30]  ( .D(n13426), .SI(\mem3[120][29] ), .SE(test_se), 
        .CLK(n1821), .Q(\mem3[120][30] ), .QN(n28730) );
  SDFFX1 \mem3_reg[120][29]  ( .D(n13425), .SI(\mem3[120][28] ), .SE(test_se), 
        .CLK(n1821), .Q(\mem3[120][29] ), .QN(n28731) );
  SDFFX1 \mem3_reg[120][28]  ( .D(n13424), .SI(\mem3[120][27] ), .SE(test_se), 
        .CLK(n1821), .Q(\mem3[120][28] ), .QN(n28732) );
  SDFFX1 \mem3_reg[120][27]  ( .D(n13423), .SI(\mem3[120][26] ), .SE(test_se), 
        .CLK(n1821), .Q(\mem3[120][27] ), .QN(n28733) );
  SDFFX1 \mem3_reg[120][26]  ( .D(n13422), .SI(\mem3[120][25] ), .SE(test_se), 
        .CLK(n1821), .Q(\mem3[120][26] ), .QN(n28734) );
  SDFFX1 \mem3_reg[120][25]  ( .D(n13421), .SI(\mem3[120][24] ), .SE(test_se), 
        .CLK(n1821), .Q(\mem3[120][25] ), .QN(n28735) );
  SDFFX1 \mem3_reg[120][24]  ( .D(n13420), .SI(\mem3[119][31] ), .SE(test_se), 
        .CLK(n1822), .Q(\mem3[120][24] ), .QN(n28736) );
  SDFFX1 \mem3_reg[119][31]  ( .D(n13419), .SI(\mem3[119][30] ), .SE(test_se), 
        .CLK(n1822), .Q(\mem3[119][31] ), .QN(n28737) );
  SDFFX1 \mem3_reg[119][30]  ( .D(n13418), .SI(\mem3[119][29] ), .SE(test_se), 
        .CLK(n1822), .Q(\mem3[119][30] ), .QN(n28738) );
  SDFFX1 \mem3_reg[119][29]  ( .D(n13417), .SI(\mem3[119][28] ), .SE(test_se), 
        .CLK(n1822), .Q(\mem3[119][29] ), .QN(n28739) );
  SDFFX1 \mem3_reg[119][28]  ( .D(n13416), .SI(\mem3[119][27] ), .SE(test_se), 
        .CLK(n1822), .Q(\mem3[119][28] ), .QN(n28740) );
  SDFFX1 \mem3_reg[119][27]  ( .D(n13415), .SI(\mem3[119][26] ), .SE(test_se), 
        .CLK(n1822), .Q(\mem3[119][27] ), .QN(n28741) );
  SDFFX1 \mem3_reg[119][26]  ( .D(n13414), .SI(\mem3[119][25] ), .SE(test_se), 
        .CLK(n1822), .Q(\mem3[119][26] ), .QN(n28742) );
  SDFFX1 \mem3_reg[119][25]  ( .D(n13413), .SI(\mem3[119][24] ), .SE(test_se), 
        .CLK(n1822), .Q(\mem3[119][25] ), .QN(n28743) );
  SDFFX1 \mem3_reg[119][24]  ( .D(n13412), .SI(\mem3[118][31] ), .SE(test_se), 
        .CLK(n1822), .Q(\mem3[119][24] ), .QN(n28744) );
  SDFFX1 \mem3_reg[118][31]  ( .D(n13411), .SI(\mem3[118][30] ), .SE(test_se), 
        .CLK(n1822), .Q(\mem3[118][31] ), .QN(n28745) );
  SDFFX1 \mem3_reg[118][30]  ( .D(n13410), .SI(\mem3[118][29] ), .SE(test_se), 
        .CLK(n1822), .Q(\mem3[118][30] ), .QN(n28746) );
  SDFFX1 \mem3_reg[118][29]  ( .D(n13409), .SI(\mem3[118][28] ), .SE(test_se), 
        .CLK(n1822), .Q(\mem3[118][29] ), .QN(n28747) );
  SDFFX1 \mem3_reg[118][28]  ( .D(n13408), .SI(\mem3[118][27] ), .SE(test_se), 
        .CLK(n1823), .Q(\mem3[118][28] ), .QN(n28748) );
  SDFFX1 \mem3_reg[118][27]  ( .D(n13407), .SI(\mem3[118][26] ), .SE(test_se), 
        .CLK(n1823), .Q(\mem3[118][27] ), .QN(n28749) );
  SDFFX1 \mem3_reg[118][26]  ( .D(n13406), .SI(\mem3[118][25] ), .SE(test_se), 
        .CLK(n1823), .Q(\mem3[118][26] ), .QN(n28750) );
  SDFFX1 \mem3_reg[118][25]  ( .D(n13405), .SI(\mem3[118][24] ), .SE(test_se), 
        .CLK(n1823), .Q(\mem3[118][25] ), .QN(n28751) );
  SDFFX1 \mem3_reg[118][24]  ( .D(n13404), .SI(\mem3[117][31] ), .SE(test_se), 
        .CLK(n1823), .Q(\mem3[118][24] ), .QN(n28752) );
  SDFFX1 \mem3_reg[117][31]  ( .D(n13403), .SI(\mem3[117][30] ), .SE(test_se), 
        .CLK(n1823), .Q(\mem3[117][31] ), .QN(n28753) );
  SDFFX1 \mem3_reg[117][30]  ( .D(n13402), .SI(\mem3[117][29] ), .SE(test_se), 
        .CLK(n1823), .Q(\mem3[117][30] ), .QN(n28754) );
  SDFFX1 \mem3_reg[117][29]  ( .D(n13401), .SI(\mem3[117][28] ), .SE(test_se), 
        .CLK(n1823), .Q(\mem3[117][29] ), .QN(n28755) );
  SDFFX1 \mem3_reg[117][28]  ( .D(n13400), .SI(\mem3[117][27] ), .SE(test_se), 
        .CLK(n1823), .Q(\mem3[117][28] ), .QN(n28756) );
  SDFFX1 \mem3_reg[117][27]  ( .D(n13399), .SI(\mem3[117][26] ), .SE(test_se), 
        .CLK(n1823), .Q(\mem3[117][27] ), .QN(n28757) );
  SDFFX1 \mem3_reg[117][26]  ( .D(n13398), .SI(\mem3[117][25] ), .SE(test_se), 
        .CLK(n1823), .Q(\mem3[117][26] ), .QN(n28758) );
  SDFFX1 \mem3_reg[117][25]  ( .D(n13397), .SI(\mem3[117][24] ), .SE(test_se), 
        .CLK(n1823), .Q(\mem3[117][25] ), .QN(n28759) );
  SDFFX1 \mem3_reg[117][24]  ( .D(n13396), .SI(\mem3[116][31] ), .SE(test_se), 
        .CLK(n1824), .Q(\mem3[117][24] ), .QN(n28760) );
  SDFFX1 \mem3_reg[116][31]  ( .D(n13395), .SI(\mem3[116][30] ), .SE(test_se), 
        .CLK(n1824), .Q(\mem3[116][31] ), .QN(n28761) );
  SDFFX1 \mem3_reg[116][30]  ( .D(n13394), .SI(\mem3[116][29] ), .SE(test_se), 
        .CLK(n1824), .Q(\mem3[116][30] ), .QN(n28762) );
  SDFFX1 \mem3_reg[116][29]  ( .D(n13393), .SI(\mem3[116][28] ), .SE(test_se), 
        .CLK(n1824), .Q(\mem3[116][29] ), .QN(n28763) );
  SDFFX1 \mem3_reg[116][28]  ( .D(n13392), .SI(\mem3[116][27] ), .SE(test_se), 
        .CLK(n1824), .Q(\mem3[116][28] ), .QN(n28764) );
  SDFFX1 \mem3_reg[116][27]  ( .D(n13391), .SI(\mem3[116][26] ), .SE(test_se), 
        .CLK(n1824), .Q(\mem3[116][27] ), .QN(n28765) );
  SDFFX1 \mem3_reg[116][26]  ( .D(n13390), .SI(\mem3[116][25] ), .SE(test_se), 
        .CLK(n1824), .Q(\mem3[116][26] ), .QN(n28766) );
  SDFFX1 \mem3_reg[116][25]  ( .D(n13389), .SI(\mem3[116][24] ), .SE(test_se), 
        .CLK(n1824), .Q(\mem3[116][25] ), .QN(n28767) );
  SDFFX1 \mem3_reg[116][24]  ( .D(n13388), .SI(\mem3[115][31] ), .SE(test_se), 
        .CLK(n1824), .Q(\mem3[116][24] ), .QN(n28768) );
  SDFFX1 \mem3_reg[115][31]  ( .D(n13387), .SI(\mem3[115][30] ), .SE(test_se), 
        .CLK(n1824), .Q(\mem3[115][31] ), .QN(n28769) );
  SDFFX1 \mem3_reg[115][30]  ( .D(n13386), .SI(\mem3[115][29] ), .SE(test_se), 
        .CLK(n1824), .Q(\mem3[115][30] ), .QN(n28770) );
  SDFFX1 \mem3_reg[115][29]  ( .D(n13385), .SI(\mem3[115][28] ), .SE(test_se), 
        .CLK(n1824), .Q(\mem3[115][29] ), .QN(n28771) );
  SDFFX1 \mem3_reg[115][28]  ( .D(n13384), .SI(\mem3[115][27] ), .SE(test_se), 
        .CLK(n1825), .Q(\mem3[115][28] ), .QN(n28772) );
  SDFFX1 \mem3_reg[115][27]  ( .D(n13383), .SI(\mem3[115][26] ), .SE(test_se), 
        .CLK(n1825), .Q(\mem3[115][27] ), .QN(n28773) );
  SDFFX1 \mem3_reg[115][26]  ( .D(n13382), .SI(\mem3[115][25] ), .SE(test_se), 
        .CLK(n1825), .Q(\mem3[115][26] ), .QN(n28774) );
  SDFFX1 \mem3_reg[115][25]  ( .D(n13381), .SI(\mem3[115][24] ), .SE(test_se), 
        .CLK(n1825), .Q(\mem3[115][25] ), .QN(n28775) );
  SDFFX1 \mem3_reg[115][24]  ( .D(n13380), .SI(\mem3[114][31] ), .SE(test_se), 
        .CLK(n1825), .Q(\mem3[115][24] ), .QN(n28776) );
  SDFFX1 \mem3_reg[114][31]  ( .D(n13379), .SI(\mem3[114][30] ), .SE(test_se), 
        .CLK(n1825), .Q(\mem3[114][31] ), .QN(n28777) );
  SDFFX1 \mem3_reg[114][30]  ( .D(n13378), .SI(\mem3[114][29] ), .SE(test_se), 
        .CLK(n1825), .Q(\mem3[114][30] ), .QN(n28778) );
  SDFFX1 \mem3_reg[114][29]  ( .D(n13377), .SI(\mem3[114][28] ), .SE(test_se), 
        .CLK(n1825), .Q(\mem3[114][29] ), .QN(n28779) );
  SDFFX1 \mem3_reg[114][28]  ( .D(n13376), .SI(\mem3[114][27] ), .SE(test_se), 
        .CLK(n1825), .Q(\mem3[114][28] ), .QN(n28780) );
  SDFFX1 \mem3_reg[114][27]  ( .D(n13375), .SI(\mem3[114][26] ), .SE(test_se), 
        .CLK(n1825), .Q(\mem3[114][27] ), .QN(n28781) );
  SDFFX1 \mem3_reg[114][26]  ( .D(n13374), .SI(\mem3[114][25] ), .SE(test_se), 
        .CLK(n1825), .Q(\mem3[114][26] ), .QN(n28782) );
  SDFFX1 \mem3_reg[114][25]  ( .D(n13373), .SI(\mem3[114][24] ), .SE(test_se), 
        .CLK(n1825), .Q(\mem3[114][25] ), .QN(n28783) );
  SDFFX1 \mem3_reg[114][24]  ( .D(n13372), .SI(\mem3[113][31] ), .SE(test_se), 
        .CLK(n1826), .Q(\mem3[114][24] ), .QN(n28784) );
  SDFFX1 \mem3_reg[113][31]  ( .D(n13371), .SI(\mem3[113][30] ), .SE(test_se), 
        .CLK(n1826), .Q(\mem3[113][31] ), .QN(n28785) );
  SDFFX1 \mem3_reg[113][30]  ( .D(n13370), .SI(\mem3[113][29] ), .SE(test_se), 
        .CLK(n1826), .Q(\mem3[113][30] ), .QN(n28786) );
  SDFFX1 \mem3_reg[113][29]  ( .D(n13369), .SI(\mem3[113][28] ), .SE(test_se), 
        .CLK(n1826), .Q(\mem3[113][29] ), .QN(n28787) );
  SDFFX1 \mem3_reg[113][28]  ( .D(n13368), .SI(\mem3[113][27] ), .SE(test_se), 
        .CLK(n1826), .Q(\mem3[113][28] ), .QN(n28788) );
  SDFFX1 \mem3_reg[113][27]  ( .D(n13367), .SI(\mem3[113][26] ), .SE(test_se), 
        .CLK(n1826), .Q(\mem3[113][27] ), .QN(n28789) );
  SDFFX1 \mem3_reg[113][26]  ( .D(n13366), .SI(\mem3[113][25] ), .SE(test_se), 
        .CLK(n1826), .Q(\mem3[113][26] ), .QN(n28790) );
  SDFFX1 \mem3_reg[113][25]  ( .D(n13365), .SI(\mem3[113][24] ), .SE(test_se), 
        .CLK(n1826), .Q(\mem3[113][25] ), .QN(n28791) );
  SDFFX1 \mem3_reg[113][24]  ( .D(n13364), .SI(\mem3[112][31] ), .SE(test_se), 
        .CLK(n1826), .Q(\mem3[113][24] ), .QN(n28792) );
  SDFFX1 \mem3_reg[112][31]  ( .D(n13363), .SI(\mem3[112][30] ), .SE(test_se), 
        .CLK(n1826), .Q(\mem3[112][31] ), .QN(n28793) );
  SDFFX1 \mem3_reg[112][30]  ( .D(n13362), .SI(\mem3[112][29] ), .SE(test_se), 
        .CLK(n1826), .Q(\mem3[112][30] ), .QN(n28794) );
  SDFFX1 \mem3_reg[112][29]  ( .D(n13361), .SI(\mem3[112][28] ), .SE(test_se), 
        .CLK(n1826), .Q(\mem3[112][29] ), .QN(n28795) );
  SDFFX1 \mem3_reg[112][28]  ( .D(n13360), .SI(\mem3[112][27] ), .SE(test_se), 
        .CLK(n1827), .Q(\mem3[112][28] ), .QN(n28796) );
  SDFFX1 \mem3_reg[112][27]  ( .D(n13359), .SI(\mem3[112][26] ), .SE(test_se), 
        .CLK(n1827), .Q(\mem3[112][27] ), .QN(n28797) );
  SDFFX1 \mem3_reg[112][26]  ( .D(n13358), .SI(\mem3[112][25] ), .SE(test_se), 
        .CLK(n1827), .Q(\mem3[112][26] ), .QN(n28798) );
  SDFFX1 \mem3_reg[112][25]  ( .D(n13357), .SI(\mem3[112][24] ), .SE(test_se), 
        .CLK(n1827), .Q(\mem3[112][25] ), .QN(n28799) );
  SDFFX1 \mem3_reg[112][24]  ( .D(n13356), .SI(\mem3[111][31] ), .SE(test_se), 
        .CLK(n1827), .Q(\mem3[112][24] ), .QN(n28800) );
  SDFFX1 \mem3_reg[111][31]  ( .D(n13355), .SI(\mem3[111][30] ), .SE(test_se), 
        .CLK(n1827), .Q(\mem3[111][31] ), .QN(n28801) );
  SDFFX1 \mem3_reg[111][30]  ( .D(n13354), .SI(\mem3[111][29] ), .SE(test_se), 
        .CLK(n1827), .Q(\mem3[111][30] ), .QN(n28802) );
  SDFFX1 \mem3_reg[111][29]  ( .D(n13353), .SI(\mem3[111][28] ), .SE(test_se), 
        .CLK(n1827), .Q(\mem3[111][29] ), .QN(n28803) );
  SDFFX1 \mem3_reg[111][28]  ( .D(n13352), .SI(\mem3[111][27] ), .SE(test_se), 
        .CLK(n1827), .Q(\mem3[111][28] ), .QN(n28804) );
  SDFFX1 \mem3_reg[111][27]  ( .D(n13351), .SI(\mem3[111][26] ), .SE(test_se), 
        .CLK(n1827), .Q(\mem3[111][27] ), .QN(n28805) );
  SDFFX1 \mem3_reg[111][26]  ( .D(n13350), .SI(\mem3[111][25] ), .SE(test_se), 
        .CLK(n1827), .Q(\mem3[111][26] ), .QN(n28806) );
  SDFFX1 \mem3_reg[111][25]  ( .D(n13349), .SI(\mem3[111][24] ), .SE(test_se), 
        .CLK(n1827), .Q(\mem3[111][25] ), .QN(n28807) );
  SDFFX1 \mem3_reg[111][24]  ( .D(n13348), .SI(\mem3[110][31] ), .SE(test_se), 
        .CLK(n1828), .Q(\mem3[111][24] ), .QN(n28808) );
  SDFFX1 \mem3_reg[110][31]  ( .D(n13347), .SI(\mem3[110][30] ), .SE(test_se), 
        .CLK(n1828), .Q(\mem3[110][31] ), .QN(n28809) );
  SDFFX1 \mem3_reg[110][30]  ( .D(n13346), .SI(\mem3[110][29] ), .SE(test_se), 
        .CLK(n1828), .Q(\mem3[110][30] ), .QN(n28810) );
  SDFFX1 \mem3_reg[110][29]  ( .D(n13345), .SI(\mem3[110][28] ), .SE(test_se), 
        .CLK(n1828), .Q(\mem3[110][29] ), .QN(n28811) );
  SDFFX1 \mem3_reg[110][28]  ( .D(n13344), .SI(\mem3[110][27] ), .SE(test_se), 
        .CLK(n1828), .Q(\mem3[110][28] ), .QN(n28812) );
  SDFFX1 \mem3_reg[110][27]  ( .D(n13343), .SI(\mem3[110][26] ), .SE(test_se), 
        .CLK(n1828), .Q(\mem3[110][27] ), .QN(n28813) );
  SDFFX1 \mem3_reg[110][26]  ( .D(n13342), .SI(\mem3[110][25] ), .SE(test_se), 
        .CLK(n1828), .Q(\mem3[110][26] ), .QN(n28814) );
  SDFFX1 \mem3_reg[110][25]  ( .D(n13341), .SI(\mem3[110][24] ), .SE(test_se), 
        .CLK(n1828), .Q(\mem3[110][25] ), .QN(n28815) );
  SDFFX1 \mem3_reg[110][24]  ( .D(n13340), .SI(\mem3[109][31] ), .SE(test_se), 
        .CLK(n1828), .Q(\mem3[110][24] ), .QN(n28816) );
  SDFFX1 \mem3_reg[109][31]  ( .D(n13339), .SI(\mem3[109][30] ), .SE(test_se), 
        .CLK(n1828), .Q(\mem3[109][31] ), .QN(n28817) );
  SDFFX1 \mem3_reg[109][30]  ( .D(n13338), .SI(\mem3[109][29] ), .SE(test_se), 
        .CLK(n1828), .Q(\mem3[109][30] ), .QN(n28818) );
  SDFFX1 \mem3_reg[109][29]  ( .D(n13337), .SI(\mem3[109][28] ), .SE(test_se), 
        .CLK(n1828), .Q(\mem3[109][29] ), .QN(n28819) );
  SDFFX1 \mem3_reg[109][28]  ( .D(n13336), .SI(\mem3[109][27] ), .SE(test_se), 
        .CLK(n1829), .Q(\mem3[109][28] ), .QN(n28820) );
  SDFFX1 \mem3_reg[109][27]  ( .D(n13335), .SI(\mem3[109][26] ), .SE(test_se), 
        .CLK(n1829), .Q(\mem3[109][27] ), .QN(n28821) );
  SDFFX1 \mem3_reg[109][26]  ( .D(n13334), .SI(\mem3[109][25] ), .SE(test_se), 
        .CLK(n1829), .Q(\mem3[109][26] ), .QN(n28822) );
  SDFFX1 \mem3_reg[109][25]  ( .D(n13333), .SI(\mem3[109][24] ), .SE(test_se), 
        .CLK(n1829), .Q(\mem3[109][25] ), .QN(n28823) );
  SDFFX1 \mem3_reg[109][24]  ( .D(n13332), .SI(\mem3[108][31] ), .SE(test_se), 
        .CLK(n1829), .Q(\mem3[109][24] ), .QN(n28824) );
  SDFFX1 \mem3_reg[108][31]  ( .D(n13331), .SI(\mem3[108][30] ), .SE(test_se), 
        .CLK(n1829), .Q(\mem3[108][31] ), .QN(n28825) );
  SDFFX1 \mem3_reg[108][30]  ( .D(n13330), .SI(\mem3[108][29] ), .SE(test_se), 
        .CLK(n1829), .Q(\mem3[108][30] ), .QN(n28826) );
  SDFFX1 \mem3_reg[108][29]  ( .D(n13329), .SI(\mem3[108][28] ), .SE(test_se), 
        .CLK(n1829), .Q(\mem3[108][29] ), .QN(n28827) );
  SDFFX1 \mem3_reg[108][28]  ( .D(n13328), .SI(\mem3[108][27] ), .SE(test_se), 
        .CLK(n1829), .Q(\mem3[108][28] ), .QN(n28828) );
  SDFFX1 \mem3_reg[108][27]  ( .D(n13327), .SI(\mem3[108][26] ), .SE(test_se), 
        .CLK(n1829), .Q(\mem3[108][27] ), .QN(n28829) );
  SDFFX1 \mem3_reg[108][26]  ( .D(n13326), .SI(\mem3[108][25] ), .SE(test_se), 
        .CLK(n1829), .Q(\mem3[108][26] ), .QN(n28830) );
  SDFFX1 \mem3_reg[108][25]  ( .D(n13325), .SI(\mem3[108][24] ), .SE(test_se), 
        .CLK(n1829), .Q(\mem3[108][25] ), .QN(n28831) );
  SDFFX1 \mem3_reg[108][24]  ( .D(n13324), .SI(\mem3[107][31] ), .SE(test_se), 
        .CLK(n1830), .Q(\mem3[108][24] ), .QN(n28832) );
  SDFFX1 \mem3_reg[107][31]  ( .D(n13323), .SI(\mem3[107][30] ), .SE(test_se), 
        .CLK(n1830), .Q(\mem3[107][31] ), .QN(n28833) );
  SDFFX1 \mem3_reg[107][30]  ( .D(n13322), .SI(\mem3[107][29] ), .SE(test_se), 
        .CLK(n1830), .Q(\mem3[107][30] ), .QN(n28834) );
  SDFFX1 \mem3_reg[107][29]  ( .D(n13321), .SI(\mem3[107][28] ), .SE(test_se), 
        .CLK(n1830), .Q(\mem3[107][29] ), .QN(n28835) );
  SDFFX1 \mem3_reg[107][28]  ( .D(n13320), .SI(\mem3[107][27] ), .SE(test_se), 
        .CLK(n1830), .Q(\mem3[107][28] ), .QN(n28836) );
  SDFFX1 \mem3_reg[107][27]  ( .D(n13319), .SI(\mem3[107][26] ), .SE(test_se), 
        .CLK(n1830), .Q(\mem3[107][27] ), .QN(n28837) );
  SDFFX1 \mem3_reg[107][26]  ( .D(n13318), .SI(\mem3[107][25] ), .SE(test_se), 
        .CLK(n1830), .Q(\mem3[107][26] ), .QN(n28838) );
  SDFFX1 \mem3_reg[107][25]  ( .D(n13317), .SI(\mem3[107][24] ), .SE(test_se), 
        .CLK(n1830), .Q(\mem3[107][25] ), .QN(n28839) );
  SDFFX1 \mem3_reg[107][24]  ( .D(n13316), .SI(\mem3[106][31] ), .SE(test_se), 
        .CLK(n1830), .Q(\mem3[107][24] ), .QN(n28840) );
  SDFFX1 \mem3_reg[106][31]  ( .D(n13315), .SI(\mem3[106][30] ), .SE(test_se), 
        .CLK(n1830), .Q(\mem3[106][31] ), .QN(n28841) );
  SDFFX1 \mem3_reg[106][30]  ( .D(n13314), .SI(\mem3[106][29] ), .SE(test_se), 
        .CLK(n1830), .Q(\mem3[106][30] ), .QN(n28842) );
  SDFFX1 \mem3_reg[106][29]  ( .D(n13313), .SI(\mem3[106][28] ), .SE(test_se), 
        .CLK(n1830), .Q(\mem3[106][29] ), .QN(n28843) );
  SDFFX1 \mem3_reg[106][28]  ( .D(n13312), .SI(\mem3[106][27] ), .SE(test_se), 
        .CLK(n1831), .Q(\mem3[106][28] ), .QN(n28844) );
  SDFFX1 \mem3_reg[106][27]  ( .D(n13311), .SI(\mem3[106][26] ), .SE(test_se), 
        .CLK(n1831), .Q(\mem3[106][27] ), .QN(n28845) );
  SDFFX1 \mem3_reg[106][26]  ( .D(n13310), .SI(\mem3[106][25] ), .SE(test_se), 
        .CLK(n1831), .Q(\mem3[106][26] ), .QN(n28846) );
  SDFFX1 \mem3_reg[106][25]  ( .D(n13309), .SI(\mem3[106][24] ), .SE(test_se), 
        .CLK(n1831), .Q(\mem3[106][25] ), .QN(n28847) );
  SDFFX1 \mem3_reg[106][24]  ( .D(n13308), .SI(\mem3[105][31] ), .SE(test_se), 
        .CLK(n1831), .Q(\mem3[106][24] ), .QN(n28848) );
  SDFFX1 \mem3_reg[105][31]  ( .D(n13307), .SI(\mem3[105][30] ), .SE(test_se), 
        .CLK(n1831), .Q(\mem3[105][31] ), .QN(n28849) );
  SDFFX1 \mem3_reg[105][30]  ( .D(n13306), .SI(\mem3[105][29] ), .SE(test_se), 
        .CLK(n1831), .Q(\mem3[105][30] ), .QN(n28850) );
  SDFFX1 \mem3_reg[105][29]  ( .D(n13305), .SI(\mem3[105][28] ), .SE(test_se), 
        .CLK(n1831), .Q(\mem3[105][29] ), .QN(n28851) );
  SDFFX1 \mem3_reg[105][28]  ( .D(n13304), .SI(\mem3[105][27] ), .SE(test_se), 
        .CLK(n1831), .Q(\mem3[105][28] ), .QN(n28852) );
  SDFFX1 \mem3_reg[105][27]  ( .D(n13303), .SI(\mem3[105][26] ), .SE(test_se), 
        .CLK(n1831), .Q(\mem3[105][27] ), .QN(n28853) );
  SDFFX1 \mem3_reg[105][26]  ( .D(n13302), .SI(\mem3[105][25] ), .SE(test_se), 
        .CLK(n1831), .Q(\mem3[105][26] ), .QN(n28854) );
  SDFFX1 \mem3_reg[105][25]  ( .D(n13301), .SI(\mem3[105][24] ), .SE(test_se), 
        .CLK(n1831), .Q(\mem3[105][25] ), .QN(n28855) );
  SDFFX1 \mem3_reg[105][24]  ( .D(n13300), .SI(\mem3[104][31] ), .SE(test_se), 
        .CLK(n1832), .Q(\mem3[105][24] ), .QN(n28856) );
  SDFFX1 \mem3_reg[104][31]  ( .D(n13299), .SI(\mem3[104][30] ), .SE(test_se), 
        .CLK(n1832), .Q(\mem3[104][31] ), .QN(n28857) );
  SDFFX1 \mem3_reg[104][30]  ( .D(n13298), .SI(\mem3[104][29] ), .SE(test_se), 
        .CLK(n1832), .Q(\mem3[104][30] ), .QN(n28858) );
  SDFFX1 \mem3_reg[104][29]  ( .D(n13297), .SI(\mem3[104][28] ), .SE(test_se), 
        .CLK(n1832), .Q(\mem3[104][29] ), .QN(n28859) );
  SDFFX1 \mem3_reg[104][28]  ( .D(n13296), .SI(\mem3[104][27] ), .SE(test_se), 
        .CLK(n1832), .Q(\mem3[104][28] ), .QN(n28860) );
  SDFFX1 \mem3_reg[104][27]  ( .D(n13295), .SI(\mem3[104][26] ), .SE(test_se), 
        .CLK(n1832), .Q(\mem3[104][27] ), .QN(n28861) );
  SDFFX1 \mem3_reg[104][26]  ( .D(n13294), .SI(\mem3[104][25] ), .SE(test_se), 
        .CLK(n1832), .Q(\mem3[104][26] ), .QN(n28862) );
  SDFFX1 \mem3_reg[104][25]  ( .D(n13293), .SI(\mem3[104][24] ), .SE(test_se), 
        .CLK(n1832), .Q(\mem3[104][25] ), .QN(n28863) );
  SDFFX1 \mem3_reg[104][24]  ( .D(n13292), .SI(\mem3[103][31] ), .SE(test_se), 
        .CLK(n1832), .Q(\mem3[104][24] ), .QN(n28864) );
  SDFFX1 \mem3_reg[103][31]  ( .D(n13291), .SI(\mem3[103][30] ), .SE(test_se), 
        .CLK(n1832), .Q(\mem3[103][31] ), .QN(n28865) );
  SDFFX1 \mem3_reg[103][30]  ( .D(n13290), .SI(\mem3[103][29] ), .SE(test_se), 
        .CLK(n1832), .Q(\mem3[103][30] ), .QN(n28866) );
  SDFFX1 \mem3_reg[103][29]  ( .D(n13289), .SI(\mem3[103][28] ), .SE(test_se), 
        .CLK(n1832), .Q(\mem3[103][29] ), .QN(n28867) );
  SDFFX1 \mem3_reg[103][28]  ( .D(n13288), .SI(\mem3[103][27] ), .SE(test_se), 
        .CLK(n1833), .Q(\mem3[103][28] ), .QN(n28868) );
  SDFFX1 \mem3_reg[103][27]  ( .D(n13287), .SI(\mem3[103][26] ), .SE(test_se), 
        .CLK(n1833), .Q(\mem3[103][27] ), .QN(n28869) );
  SDFFX1 \mem3_reg[103][26]  ( .D(n13286), .SI(\mem3[103][25] ), .SE(test_se), 
        .CLK(n1833), .Q(\mem3[103][26] ), .QN(n28870) );
  SDFFX1 \mem3_reg[103][25]  ( .D(n13285), .SI(\mem3[103][24] ), .SE(test_se), 
        .CLK(n1833), .Q(\mem3[103][25] ), .QN(n28871) );
  SDFFX1 \mem3_reg[103][24]  ( .D(n13284), .SI(\mem3[102][31] ), .SE(test_se), 
        .CLK(n1833), .Q(\mem3[103][24] ), .QN(n28872) );
  SDFFX1 \mem3_reg[102][31]  ( .D(n13283), .SI(\mem3[102][30] ), .SE(test_se), 
        .CLK(n1833), .Q(\mem3[102][31] ), .QN(n28873) );
  SDFFX1 \mem3_reg[102][30]  ( .D(n13282), .SI(\mem3[102][29] ), .SE(test_se), 
        .CLK(n1833), .Q(\mem3[102][30] ), .QN(n28874) );
  SDFFX1 \mem3_reg[102][29]  ( .D(n13281), .SI(\mem3[102][28] ), .SE(test_se), 
        .CLK(n1833), .Q(\mem3[102][29] ), .QN(n28875) );
  SDFFX1 \mem3_reg[102][28]  ( .D(n13280), .SI(\mem3[102][27] ), .SE(test_se), 
        .CLK(n1833), .Q(\mem3[102][28] ), .QN(n28876) );
  SDFFX1 \mem3_reg[102][27]  ( .D(n13279), .SI(\mem3[102][26] ), .SE(test_se), 
        .CLK(n1833), .Q(\mem3[102][27] ), .QN(n28877) );
  SDFFX1 \mem3_reg[102][26]  ( .D(n13278), .SI(\mem3[102][25] ), .SE(test_se), 
        .CLK(n1833), .Q(\mem3[102][26] ), .QN(n28878) );
  SDFFX1 \mem3_reg[102][25]  ( .D(n13277), .SI(\mem3[102][24] ), .SE(test_se), 
        .CLK(n1833), .Q(\mem3[102][25] ), .QN(n28879) );
  SDFFX1 \mem3_reg[102][24]  ( .D(n13276), .SI(\mem3[101][31] ), .SE(test_se), 
        .CLK(n1834), .Q(\mem3[102][24] ), .QN(n28880) );
  SDFFX1 \mem3_reg[101][31]  ( .D(n13275), .SI(\mem3[101][30] ), .SE(test_se), 
        .CLK(n1834), .Q(\mem3[101][31] ), .QN(n28881) );
  SDFFX1 \mem3_reg[101][30]  ( .D(n13274), .SI(\mem3[101][29] ), .SE(test_se), 
        .CLK(n1834), .Q(\mem3[101][30] ), .QN(n28882) );
  SDFFX1 \mem3_reg[101][29]  ( .D(n13273), .SI(\mem3[101][28] ), .SE(test_se), 
        .CLK(n1834), .Q(\mem3[101][29] ), .QN(n28883) );
  SDFFX1 \mem3_reg[101][28]  ( .D(n13272), .SI(\mem3[101][27] ), .SE(test_se), 
        .CLK(n1834), .Q(\mem3[101][28] ), .QN(n28884) );
  SDFFX1 \mem3_reg[101][27]  ( .D(n13271), .SI(\mem3[101][26] ), .SE(test_se), 
        .CLK(n1834), .Q(\mem3[101][27] ), .QN(n28885) );
  SDFFX1 \mem3_reg[101][26]  ( .D(n13270), .SI(\mem3[101][25] ), .SE(test_se), 
        .CLK(n1834), .Q(\mem3[101][26] ), .QN(n28886) );
  SDFFX1 \mem3_reg[101][25]  ( .D(n13269), .SI(\mem3[101][24] ), .SE(test_se), 
        .CLK(n1834), .Q(\mem3[101][25] ), .QN(n28887) );
  SDFFX1 \mem3_reg[101][24]  ( .D(n13268), .SI(\mem3[100][31] ), .SE(test_se), 
        .CLK(n1834), .Q(\mem3[101][24] ), .QN(n28888) );
  SDFFX1 \mem3_reg[100][31]  ( .D(n13267), .SI(\mem3[100][30] ), .SE(test_se), 
        .CLK(n1834), .Q(\mem3[100][31] ), .QN(n28889) );
  SDFFX1 \mem3_reg[100][30]  ( .D(n13266), .SI(\mem3[100][29] ), .SE(test_se), 
        .CLK(n1834), .Q(\mem3[100][30] ), .QN(n28890) );
  SDFFX1 \mem3_reg[100][29]  ( .D(n13265), .SI(\mem3[100][28] ), .SE(test_se), 
        .CLK(n1834), .Q(\mem3[100][29] ), .QN(n28891) );
  SDFFX1 \mem3_reg[100][28]  ( .D(n13264), .SI(\mem3[100][27] ), .SE(test_se), 
        .CLK(n1835), .Q(\mem3[100][28] ), .QN(n28892) );
  SDFFX1 \mem3_reg[100][27]  ( .D(n13263), .SI(\mem3[100][26] ), .SE(test_se), 
        .CLK(n1835), .Q(\mem3[100][27] ), .QN(n28893) );
  SDFFX1 \mem3_reg[100][26]  ( .D(n13262), .SI(\mem3[100][25] ), .SE(test_se), 
        .CLK(n1835), .Q(\mem3[100][26] ), .QN(n28894) );
  SDFFX1 \mem3_reg[100][25]  ( .D(n13261), .SI(\mem3[100][24] ), .SE(test_se), 
        .CLK(n1835), .Q(\mem3[100][25] ), .QN(n28895) );
  SDFFX1 \mem3_reg[100][24]  ( .D(n13260), .SI(\mem3[99][31] ), .SE(test_se), 
        .CLK(n1835), .Q(\mem3[100][24] ), .QN(n28896) );
  SDFFX1 \mem3_reg[99][31]  ( .D(n13259), .SI(\mem3[99][30] ), .SE(test_se), 
        .CLK(n1835), .Q(\mem3[99][31] ), .QN(n28897) );
  SDFFX1 \mem3_reg[99][30]  ( .D(n13258), .SI(\mem3[99][29] ), .SE(test_se), 
        .CLK(n1835), .Q(\mem3[99][30] ), .QN(n28898) );
  SDFFX1 \mem3_reg[99][29]  ( .D(n13257), .SI(\mem3[99][28] ), .SE(test_se), 
        .CLK(n1835), .Q(\mem3[99][29] ), .QN(n28899) );
  SDFFX1 \mem3_reg[99][28]  ( .D(n13256), .SI(\mem3[99][27] ), .SE(test_se), 
        .CLK(n1835), .Q(\mem3[99][28] ), .QN(n28900) );
  SDFFX1 \mem3_reg[99][27]  ( .D(n13255), .SI(\mem3[99][26] ), .SE(test_se), 
        .CLK(n1835), .Q(\mem3[99][27] ), .QN(n28901) );
  SDFFX1 \mem3_reg[99][26]  ( .D(n13254), .SI(\mem3[99][25] ), .SE(test_se), 
        .CLK(n1835), .Q(\mem3[99][26] ), .QN(n28902) );
  SDFFX1 \mem3_reg[99][25]  ( .D(n13253), .SI(\mem3[99][24] ), .SE(test_se), 
        .CLK(n1835), .Q(\mem3[99][25] ), .QN(n28903) );
  SDFFX1 \mem3_reg[99][24]  ( .D(n13252), .SI(\mem3[98][31] ), .SE(test_se), 
        .CLK(n1836), .Q(\mem3[99][24] ), .QN(n28904) );
  SDFFX1 \mem3_reg[98][31]  ( .D(n13251), .SI(\mem3[98][30] ), .SE(test_se), 
        .CLK(n1836), .Q(\mem3[98][31] ), .QN(n28905) );
  SDFFX1 \mem3_reg[98][30]  ( .D(n13250), .SI(\mem3[98][29] ), .SE(test_se), 
        .CLK(n1836), .Q(\mem3[98][30] ), .QN(n28906) );
  SDFFX1 \mem3_reg[98][29]  ( .D(n13249), .SI(\mem3[98][28] ), .SE(test_se), 
        .CLK(n1836), .Q(\mem3[98][29] ), .QN(n28907) );
  SDFFX1 \mem3_reg[98][28]  ( .D(n13248), .SI(\mem3[98][27] ), .SE(test_se), 
        .CLK(n1836), .Q(\mem3[98][28] ), .QN(n28908) );
  SDFFX1 \mem3_reg[98][27]  ( .D(n13247), .SI(\mem3[98][26] ), .SE(test_se), 
        .CLK(n1836), .Q(\mem3[98][27] ), .QN(n28909) );
  SDFFX1 \mem3_reg[98][26]  ( .D(n13246), .SI(\mem3[98][25] ), .SE(test_se), 
        .CLK(n1836), .Q(\mem3[98][26] ), .QN(n28910) );
  SDFFX1 \mem3_reg[98][25]  ( .D(n13245), .SI(\mem3[98][24] ), .SE(test_se), 
        .CLK(n1836), .Q(\mem3[98][25] ), .QN(n28911) );
  SDFFX1 \mem3_reg[98][24]  ( .D(n13244), .SI(\mem3[97][31] ), .SE(test_se), 
        .CLK(n1836), .Q(\mem3[98][24] ), .QN(n28912) );
  SDFFX1 \mem3_reg[97][31]  ( .D(n13243), .SI(\mem3[97][30] ), .SE(test_se), 
        .CLK(n1836), .Q(\mem3[97][31] ), .QN(n28913) );
  SDFFX1 \mem3_reg[97][30]  ( .D(n13242), .SI(\mem3[97][29] ), .SE(test_se), 
        .CLK(n1836), .Q(\mem3[97][30] ), .QN(n28914) );
  SDFFX1 \mem3_reg[97][29]  ( .D(n13241), .SI(\mem3[97][28] ), .SE(test_se), 
        .CLK(n1836), .Q(\mem3[97][29] ), .QN(n28915) );
  SDFFX1 \mem3_reg[97][28]  ( .D(n13240), .SI(\mem3[97][27] ), .SE(test_se), 
        .CLK(n1837), .Q(\mem3[97][28] ), .QN(n28916) );
  SDFFX1 \mem3_reg[97][27]  ( .D(n13239), .SI(\mem3[97][26] ), .SE(test_se), 
        .CLK(n1837), .Q(\mem3[97][27] ), .QN(n28917) );
  SDFFX1 \mem3_reg[97][26]  ( .D(n13238), .SI(\mem3[97][25] ), .SE(test_se), 
        .CLK(n1837), .Q(\mem3[97][26] ), .QN(n28918) );
  SDFFX1 \mem3_reg[97][25]  ( .D(n13237), .SI(\mem3[97][24] ), .SE(test_se), 
        .CLK(n1837), .Q(\mem3[97][25] ), .QN(n28919) );
  SDFFX1 \mem3_reg[97][24]  ( .D(n13236), .SI(\mem3[96][31] ), .SE(test_se), 
        .CLK(n1837), .Q(\mem3[97][24] ), .QN(n28920) );
  SDFFX1 \mem3_reg[96][31]  ( .D(n13235), .SI(\mem3[96][30] ), .SE(test_se), 
        .CLK(n1837), .Q(\mem3[96][31] ), .QN(n28921) );
  SDFFX1 \mem3_reg[96][30]  ( .D(n13234), .SI(\mem3[96][29] ), .SE(test_se), 
        .CLK(n1837), .Q(\mem3[96][30] ), .QN(n28922) );
  SDFFX1 \mem3_reg[96][29]  ( .D(n13233), .SI(\mem3[96][28] ), .SE(test_se), 
        .CLK(n1837), .Q(\mem3[96][29] ), .QN(n28923) );
  SDFFX1 \mem3_reg[96][28]  ( .D(n13232), .SI(\mem3[96][27] ), .SE(test_se), 
        .CLK(n1837), .Q(\mem3[96][28] ), .QN(n28924) );
  SDFFX1 \mem3_reg[96][27]  ( .D(n13231), .SI(\mem3[96][26] ), .SE(test_se), 
        .CLK(n1837), .Q(\mem3[96][27] ), .QN(n28925) );
  SDFFX1 \mem3_reg[96][26]  ( .D(n13230), .SI(\mem3[96][25] ), .SE(test_se), 
        .CLK(n1837), .Q(\mem3[96][26] ), .QN(n28926) );
  SDFFX1 \mem3_reg[96][25]  ( .D(n13229), .SI(\mem3[96][24] ), .SE(test_se), 
        .CLK(n1837), .Q(\mem3[96][25] ), .QN(n28927) );
  SDFFX1 \mem3_reg[96][24]  ( .D(n13228), .SI(\mem3[95][31] ), .SE(test_se), 
        .CLK(n1838), .Q(\mem3[96][24] ), .QN(n28928) );
  SDFFX1 \mem3_reg[95][31]  ( .D(n13227), .SI(\mem3[95][30] ), .SE(test_se), 
        .CLK(n1838), .Q(\mem3[95][31] ), .QN(n28929) );
  SDFFX1 \mem3_reg[95][30]  ( .D(n13226), .SI(\mem3[95][29] ), .SE(test_se), 
        .CLK(n1838), .Q(\mem3[95][30] ), .QN(n28930) );
  SDFFX1 \mem3_reg[95][29]  ( .D(n13225), .SI(\mem3[95][28] ), .SE(test_se), 
        .CLK(n1838), .Q(\mem3[95][29] ), .QN(n28931) );
  SDFFX1 \mem3_reg[95][28]  ( .D(n13224), .SI(\mem3[95][27] ), .SE(test_se), 
        .CLK(n1838), .Q(\mem3[95][28] ), .QN(n28932) );
  SDFFX1 \mem3_reg[95][27]  ( .D(n13223), .SI(\mem3[95][26] ), .SE(test_se), 
        .CLK(n1838), .Q(\mem3[95][27] ), .QN(n28933) );
  SDFFX1 \mem3_reg[95][26]  ( .D(n13222), .SI(\mem3[95][25] ), .SE(test_se), 
        .CLK(n1838), .Q(\mem3[95][26] ), .QN(n28934) );
  SDFFX1 \mem3_reg[95][25]  ( .D(n13221), .SI(\mem3[95][24] ), .SE(test_se), 
        .CLK(n1838), .Q(\mem3[95][25] ), .QN(n28935) );
  SDFFX1 \mem3_reg[95][24]  ( .D(n13220), .SI(\mem3[94][31] ), .SE(test_se), 
        .CLK(n1838), .Q(\mem3[95][24] ), .QN(n28936) );
  SDFFX1 \mem3_reg[94][31]  ( .D(n13219), .SI(\mem3[94][30] ), .SE(test_se), 
        .CLK(n1838), .Q(\mem3[94][31] ), .QN(n28937) );
  SDFFX1 \mem3_reg[94][30]  ( .D(n13218), .SI(\mem3[94][29] ), .SE(test_se), 
        .CLK(n1838), .Q(\mem3[94][30] ), .QN(n28938) );
  SDFFX1 \mem3_reg[94][29]  ( .D(n13217), .SI(\mem3[94][28] ), .SE(test_se), 
        .CLK(n1838), .Q(\mem3[94][29] ), .QN(n28939) );
  SDFFX1 \mem3_reg[94][28]  ( .D(n13216), .SI(\mem3[94][27] ), .SE(test_se), 
        .CLK(n1839), .Q(\mem3[94][28] ), .QN(n28940) );
  SDFFX1 \mem3_reg[94][27]  ( .D(n13215), .SI(\mem3[94][26] ), .SE(test_se), 
        .CLK(n1839), .Q(\mem3[94][27] ), .QN(n28941) );
  SDFFX1 \mem3_reg[94][26]  ( .D(n13214), .SI(\mem3[94][25] ), .SE(test_se), 
        .CLK(n1839), .Q(\mem3[94][26] ), .QN(n28942) );
  SDFFX1 \mem3_reg[94][25]  ( .D(n13213), .SI(\mem3[94][24] ), .SE(test_se), 
        .CLK(n1839), .Q(\mem3[94][25] ), .QN(n28943) );
  SDFFX1 \mem3_reg[94][24]  ( .D(n13212), .SI(\mem3[93][31] ), .SE(test_se), 
        .CLK(n1839), .Q(\mem3[94][24] ), .QN(n28944) );
  SDFFX1 \mem3_reg[93][31]  ( .D(n13211), .SI(\mem3[93][30] ), .SE(test_se), 
        .CLK(n1839), .Q(\mem3[93][31] ), .QN(n28945) );
  SDFFX1 \mem3_reg[93][30]  ( .D(n13210), .SI(\mem3[93][29] ), .SE(test_se), 
        .CLK(n1839), .Q(\mem3[93][30] ), .QN(n28946) );
  SDFFX1 \mem3_reg[93][29]  ( .D(n13209), .SI(\mem3[93][28] ), .SE(test_se), 
        .CLK(n1839), .Q(\mem3[93][29] ), .QN(n28947) );
  SDFFX1 \mem3_reg[93][28]  ( .D(n13208), .SI(\mem3[93][27] ), .SE(test_se), 
        .CLK(n1839), .Q(\mem3[93][28] ), .QN(n28948) );
  SDFFX1 \mem3_reg[93][27]  ( .D(n13207), .SI(\mem3[93][26] ), .SE(test_se), 
        .CLK(n1839), .Q(\mem3[93][27] ), .QN(n28949) );
  SDFFX1 \mem3_reg[93][26]  ( .D(n13206), .SI(\mem3[93][25] ), .SE(test_se), 
        .CLK(n1839), .Q(\mem3[93][26] ), .QN(n28950) );
  SDFFX1 \mem3_reg[93][25]  ( .D(n13205), .SI(\mem3[93][24] ), .SE(test_se), 
        .CLK(n1839), .Q(\mem3[93][25] ), .QN(n28951) );
  SDFFX1 \mem3_reg[93][24]  ( .D(n13204), .SI(\mem3[92][31] ), .SE(test_se), 
        .CLK(n1840), .Q(\mem3[93][24] ), .QN(n28952) );
  SDFFX1 \mem3_reg[92][31]  ( .D(n13203), .SI(\mem3[92][30] ), .SE(test_se), 
        .CLK(n1840), .Q(\mem3[92][31] ), .QN(n28953) );
  SDFFX1 \mem3_reg[92][30]  ( .D(n13202), .SI(\mem3[92][29] ), .SE(test_se), 
        .CLK(n1840), .Q(\mem3[92][30] ), .QN(n28954) );
  SDFFX1 \mem3_reg[92][29]  ( .D(n13201), .SI(\mem3[92][28] ), .SE(test_se), 
        .CLK(n1840), .Q(\mem3[92][29] ), .QN(n28955) );
  SDFFX1 \mem3_reg[92][28]  ( .D(n13200), .SI(\mem3[92][27] ), .SE(test_se), 
        .CLK(n1840), .Q(\mem3[92][28] ), .QN(n28956) );
  SDFFX1 \mem3_reg[92][27]  ( .D(n13199), .SI(\mem3[92][26] ), .SE(test_se), 
        .CLK(n1840), .Q(\mem3[92][27] ), .QN(n28957) );
  SDFFX1 \mem3_reg[92][26]  ( .D(n13198), .SI(\mem3[92][25] ), .SE(test_se), 
        .CLK(n1840), .Q(\mem3[92][26] ), .QN(n28958) );
  SDFFX1 \mem3_reg[92][25]  ( .D(n13197), .SI(\mem3[92][24] ), .SE(test_se), 
        .CLK(n1840), .Q(\mem3[92][25] ), .QN(n28959) );
  SDFFX1 \mem3_reg[92][24]  ( .D(n13196), .SI(\mem3[91][31] ), .SE(test_se), 
        .CLK(n1840), .Q(\mem3[92][24] ), .QN(n28960) );
  SDFFX1 \mem3_reg[91][31]  ( .D(n13195), .SI(\mem3[91][30] ), .SE(test_se), 
        .CLK(n2047), .Q(\mem3[91][31] ), .QN(n28961) );
  SDFFX1 \mem3_reg[91][30]  ( .D(n13194), .SI(\mem3[91][29] ), .SE(test_se), 
        .CLK(n2047), .Q(\mem3[91][30] ), .QN(n28962) );
  SDFFX1 \mem3_reg[91][29]  ( .D(n13193), .SI(\mem3[91][28] ), .SE(test_se), 
        .CLK(n2048), .Q(\mem3[91][29] ), .QN(n28963) );
  SDFFX1 \mem3_reg[91][28]  ( .D(n13192), .SI(\mem3[91][27] ), .SE(test_se), 
        .CLK(n2048), .Q(\mem3[91][28] ), .QN(n28964) );
  SDFFX1 \mem3_reg[91][27]  ( .D(n13191), .SI(\mem3[91][26] ), .SE(test_se), 
        .CLK(n2048), .Q(\mem3[91][27] ), .QN(n28965) );
  SDFFX1 \mem3_reg[91][26]  ( .D(n13190), .SI(\mem3[91][25] ), .SE(test_se), 
        .CLK(n2048), .Q(\mem3[91][26] ), .QN(n28966) );
  SDFFX1 \mem3_reg[91][25]  ( .D(n13189), .SI(\mem3[91][24] ), .SE(test_se), 
        .CLK(n2048), .Q(\mem3[91][25] ), .QN(n28967) );
  SDFFX1 \mem3_reg[91][24]  ( .D(n13188), .SI(\mem3[90][31] ), .SE(test_se), 
        .CLK(n2048), .Q(\mem3[91][24] ), .QN(n28968) );
  SDFFX1 \mem3_reg[90][31]  ( .D(n13187), .SI(\mem3[90][30] ), .SE(test_se), 
        .CLK(n2048), .Q(\mem3[90][31] ), .QN(n28969) );
  SDFFX1 \mem3_reg[90][30]  ( .D(n13186), .SI(\mem3[90][29] ), .SE(test_se), 
        .CLK(n2048), .Q(\mem3[90][30] ), .QN(n28970) );
  SDFFX1 \mem3_reg[90][29]  ( .D(n13185), .SI(\mem3[90][28] ), .SE(test_se), 
        .CLK(n2048), .Q(\mem3[90][29] ), .QN(n28971) );
  SDFFX1 \mem3_reg[90][28]  ( .D(n13184), .SI(\mem3[90][27] ), .SE(test_se), 
        .CLK(n2048), .Q(\mem3[90][28] ), .QN(n28972) );
  SDFFX1 \mem3_reg[90][27]  ( .D(n13183), .SI(\mem3[90][26] ), .SE(test_se), 
        .CLK(n2048), .Q(\mem3[90][27] ), .QN(n28973) );
  SDFFX1 \mem3_reg[90][26]  ( .D(n13182), .SI(\mem3[90][25] ), .SE(test_se), 
        .CLK(n2048), .Q(\mem3[90][26] ), .QN(n28974) );
  SDFFX1 \mem3_reg[90][25]  ( .D(n13181), .SI(\mem3[90][24] ), .SE(test_se), 
        .CLK(n2049), .Q(\mem3[90][25] ), .QN(n28975) );
  SDFFX1 \mem3_reg[90][24]  ( .D(n13180), .SI(\mem3[89][31] ), .SE(test_se), 
        .CLK(n2049), .Q(\mem3[90][24] ), .QN(n28976) );
  SDFFX1 \mem3_reg[89][31]  ( .D(n13179), .SI(\mem3[89][30] ), .SE(test_se), 
        .CLK(n2049), .Q(\mem3[89][31] ), .QN(n28977) );
  SDFFX1 \mem3_reg[89][30]  ( .D(n13178), .SI(\mem3[89][29] ), .SE(test_se), 
        .CLK(n2049), .Q(\mem3[89][30] ), .QN(n28978) );
  SDFFX1 \mem3_reg[89][29]  ( .D(n13177), .SI(\mem3[89][28] ), .SE(test_se), 
        .CLK(n2049), .Q(\mem3[89][29] ), .QN(n28979) );
  SDFFX1 \mem3_reg[89][28]  ( .D(n13176), .SI(\mem3[89][27] ), .SE(test_se), 
        .CLK(n2049), .Q(\mem3[89][28] ), .QN(n28980) );
  SDFFX1 \mem3_reg[89][27]  ( .D(n13175), .SI(\mem3[89][26] ), .SE(test_se), 
        .CLK(n2049), .Q(\mem3[89][27] ), .QN(n28981) );
  SDFFX1 \mem3_reg[89][26]  ( .D(n13174), .SI(\mem3[89][25] ), .SE(test_se), 
        .CLK(n2049), .Q(\mem3[89][26] ), .QN(n28982) );
  SDFFX1 \mem3_reg[89][25]  ( .D(n13173), .SI(\mem3[89][24] ), .SE(test_se), 
        .CLK(n2049), .Q(\mem3[89][25] ), .QN(n28983) );
  SDFFX1 \mem3_reg[89][24]  ( .D(n13172), .SI(\mem3[88][31] ), .SE(test_se), 
        .CLK(n2049), .Q(\mem3[89][24] ), .QN(n28984) );
  SDFFX1 \mem3_reg[88][31]  ( .D(n13171), .SI(\mem3[88][30] ), .SE(test_se), 
        .CLK(n2049), .Q(\mem3[88][31] ), .QN(n28985) );
  SDFFX1 \mem3_reg[88][30]  ( .D(n13170), .SI(\mem3[88][29] ), .SE(test_se), 
        .CLK(n2049), .Q(\mem3[88][30] ), .QN(n28986) );
  SDFFX1 \mem3_reg[88][29]  ( .D(n13169), .SI(\mem3[88][28] ), .SE(test_se), 
        .CLK(n2050), .Q(\mem3[88][29] ), .QN(n28987) );
  SDFFX1 \mem3_reg[88][28]  ( .D(n13168), .SI(\mem3[88][27] ), .SE(test_se), 
        .CLK(n2050), .Q(\mem3[88][28] ), .QN(n28988) );
  SDFFX1 \mem3_reg[88][27]  ( .D(n13167), .SI(\mem3[88][26] ), .SE(test_se), 
        .CLK(n2050), .Q(\mem3[88][27] ), .QN(n28989) );
  SDFFX1 \mem3_reg[88][26]  ( .D(n13166), .SI(\mem3[88][25] ), .SE(test_se), 
        .CLK(n2050), .Q(\mem3[88][26] ), .QN(n28990) );
  SDFFX1 \mem3_reg[88][25]  ( .D(n13165), .SI(\mem3[88][24] ), .SE(test_se), 
        .CLK(n2050), .Q(\mem3[88][25] ), .QN(n28991) );
  SDFFX1 \mem3_reg[88][24]  ( .D(n13164), .SI(\mem3[87][31] ), .SE(test_se), 
        .CLK(n2050), .Q(\mem3[88][24] ), .QN(n28992) );
  SDFFX1 \mem3_reg[87][31]  ( .D(n13163), .SI(\mem3[87][30] ), .SE(test_se), 
        .CLK(n2058), .Q(\mem3[87][31] ), .QN(n28993) );
  SDFFX1 \mem3_reg[87][30]  ( .D(n13162), .SI(\mem3[87][29] ), .SE(test_se), 
        .CLK(n2058), .Q(\mem3[87][30] ), .QN(n28994) );
  SDFFX1 \mem3_reg[87][29]  ( .D(n13161), .SI(\mem3[87][28] ), .SE(test_se), 
        .CLK(n2058), .Q(\mem3[87][29] ), .QN(n28995) );
  SDFFX1 \mem3_reg[87][28]  ( .D(n13160), .SI(\mem3[87][27] ), .SE(test_se), 
        .CLK(n2058), .Q(\mem3[87][28] ), .QN(n28996) );
  SDFFX1 \mem3_reg[87][27]  ( .D(n13159), .SI(\mem3[87][26] ), .SE(test_se), 
        .CLK(n2058), .Q(\mem3[87][27] ), .QN(n28997) );
  SDFFX1 \mem3_reg[87][26]  ( .D(n13158), .SI(\mem3[87][25] ), .SE(test_se), 
        .CLK(n2058), .Q(\mem3[87][26] ), .QN(n28998) );
  SDFFX1 \mem3_reg[87][25]  ( .D(n13157), .SI(\mem3[87][24] ), .SE(test_se), 
        .CLK(n2059), .Q(\mem3[87][25] ), .QN(n28999) );
  SDFFX1 \mem3_reg[87][24]  ( .D(n13156), .SI(\mem3[86][31] ), .SE(test_se), 
        .CLK(n2059), .Q(\mem3[87][24] ), .QN(n29000) );
  SDFFX1 \mem3_reg[86][31]  ( .D(n13155), .SI(\mem3[86][30] ), .SE(test_se), 
        .CLK(n2059), .Q(\mem3[86][31] ), .QN(n29001) );
  SDFFX1 \mem3_reg[86][30]  ( .D(n13154), .SI(\mem3[86][29] ), .SE(test_se), 
        .CLK(n2059), .Q(\mem3[86][30] ), .QN(n29002) );
  SDFFX1 \mem3_reg[86][29]  ( .D(n13153), .SI(\mem3[86][28] ), .SE(test_se), 
        .CLK(n2059), .Q(\mem3[86][29] ), .QN(n29003) );
  SDFFX1 \mem3_reg[86][28]  ( .D(n13152), .SI(\mem3[86][27] ), .SE(test_se), 
        .CLK(n2059), .Q(\mem3[86][28] ), .QN(n29004) );
  SDFFX1 \mem3_reg[86][27]  ( .D(n13151), .SI(\mem3[86][26] ), .SE(test_se), 
        .CLK(n2059), .Q(\mem3[86][27] ), .QN(n29005) );
  SDFFX1 \mem3_reg[86][26]  ( .D(n13150), .SI(\mem3[86][25] ), .SE(test_se), 
        .CLK(n2059), .Q(\mem3[86][26] ), .QN(n29006) );
  SDFFX1 \mem3_reg[86][25]  ( .D(n13149), .SI(\mem3[86][24] ), .SE(test_se), 
        .CLK(n2059), .Q(\mem3[86][25] ), .QN(n29007) );
  SDFFX1 \mem3_reg[86][24]  ( .D(n13148), .SI(\mem3[85][31] ), .SE(test_se), 
        .CLK(n2059), .Q(\mem3[86][24] ), .QN(n29008) );
  SDFFX1 \mem3_reg[85][31]  ( .D(n13147), .SI(\mem3[85][30] ), .SE(test_se), 
        .CLK(n2059), .Q(\mem3[85][31] ), .QN(n29009) );
  SDFFX1 \mem3_reg[85][30]  ( .D(n13146), .SI(\mem3[85][29] ), .SE(test_se), 
        .CLK(n2059), .Q(\mem3[85][30] ), .QN(n29010) );
  SDFFX1 \mem3_reg[85][29]  ( .D(n13145), .SI(\mem3[85][28] ), .SE(test_se), 
        .CLK(n2060), .Q(\mem3[85][29] ), .QN(n29011) );
  SDFFX1 \mem3_reg[85][28]  ( .D(n13144), .SI(\mem3[85][27] ), .SE(test_se), 
        .CLK(n2060), .Q(\mem3[85][28] ), .QN(n29012) );
  SDFFX1 \mem3_reg[85][27]  ( .D(n13143), .SI(\mem3[85][26] ), .SE(test_se), 
        .CLK(n2060), .Q(\mem3[85][27] ), .QN(n29013) );
  SDFFX1 \mem3_reg[85][26]  ( .D(n13142), .SI(\mem3[85][25] ), .SE(test_se), 
        .CLK(n2060), .Q(\mem3[85][26] ), .QN(n29014) );
  SDFFX1 \mem3_reg[85][25]  ( .D(n13141), .SI(\mem3[85][24] ), .SE(test_se), 
        .CLK(n2060), .Q(\mem3[85][25] ), .QN(n29015) );
  SDFFX1 \mem3_reg[85][24]  ( .D(n13140), .SI(\mem3[84][31] ), .SE(test_se), 
        .CLK(n2060), .Q(\mem3[85][24] ), .QN(n29016) );
  SDFFX1 \mem3_reg[84][31]  ( .D(n13139), .SI(\mem3[84][30] ), .SE(test_se), 
        .CLK(n2060), .Q(\mem3[84][31] ), .QN(n29017) );
  SDFFX1 \mem3_reg[84][30]  ( .D(n13138), .SI(\mem3[84][29] ), .SE(test_se), 
        .CLK(n2060), .Q(\mem3[84][30] ), .QN(n29018) );
  SDFFX1 \mem3_reg[84][29]  ( .D(n13137), .SI(\mem3[84][28] ), .SE(test_se), 
        .CLK(n2060), .Q(\mem3[84][29] ), .QN(n29019) );
  SDFFX1 \mem3_reg[84][28]  ( .D(n13136), .SI(\mem3[84][27] ), .SE(test_se), 
        .CLK(n2060), .Q(\mem3[84][28] ), .QN(n29020) );
  SDFFX1 \mem3_reg[84][27]  ( .D(n13135), .SI(\mem3[84][26] ), .SE(test_se), 
        .CLK(n2060), .Q(\mem3[84][27] ), .QN(n29021) );
  SDFFX1 \mem3_reg[84][26]  ( .D(n13134), .SI(\mem3[84][25] ), .SE(test_se), 
        .CLK(n2060), .Q(\mem3[84][26] ), .QN(n29022) );
  SDFFX1 \mem3_reg[84][25]  ( .D(n13133), .SI(\mem3[84][24] ), .SE(test_se), 
        .CLK(n2061), .Q(\mem3[84][25] ), .QN(n29023) );
  SDFFX1 \mem3_reg[84][24]  ( .D(n13132), .SI(\mem3[83][31] ), .SE(test_se), 
        .CLK(n2061), .Q(\mem3[84][24] ), .QN(n29024) );
  SDFFX1 \mem3_reg[83][31]  ( .D(n13131), .SI(\mem3[83][30] ), .SE(test_se), 
        .CLK(n2066), .Q(\mem3[83][31] ), .QN(n29025) );
  SDFFX1 \mem3_reg[83][30]  ( .D(n13130), .SI(\mem3[83][29] ), .SE(test_se), 
        .CLK(n2066), .Q(\mem3[83][30] ), .QN(n29026) );
  SDFFX1 \mem3_reg[83][29]  ( .D(n13129), .SI(\mem3[83][28] ), .SE(test_se), 
        .CLK(n2066), .Q(\mem3[83][29] ), .QN(n29027) );
  SDFFX1 \mem3_reg[83][28]  ( .D(n13128), .SI(\mem3[83][27] ), .SE(test_se), 
        .CLK(n2066), .Q(\mem3[83][28] ), .QN(n29028) );
  SDFFX1 \mem3_reg[83][27]  ( .D(n13127), .SI(\mem3[83][26] ), .SE(test_se), 
        .CLK(n2066), .Q(\mem3[83][27] ), .QN(n29029) );
  SDFFX1 \mem3_reg[83][26]  ( .D(n13126), .SI(\mem3[83][25] ), .SE(test_se), 
        .CLK(n2066), .Q(\mem3[83][26] ), .QN(n29030) );
  SDFFX1 \mem3_reg[83][25]  ( .D(n13125), .SI(\mem3[83][24] ), .SE(test_se), 
        .CLK(n2066), .Q(\mem3[83][25] ), .QN(n29031) );
  SDFFX1 \mem3_reg[83][24]  ( .D(n13124), .SI(\mem3[82][31] ), .SE(test_se), 
        .CLK(n2066), .Q(\mem3[83][24] ), .QN(n29032) );
  SDFFX1 \mem3_reg[82][31]  ( .D(n13123), .SI(\mem3[82][30] ), .SE(test_se), 
        .CLK(n2067), .Q(\mem3[82][31] ), .QN(n29033) );
  SDFFX1 \mem3_reg[82][30]  ( .D(n13122), .SI(\mem3[82][29] ), .SE(test_se), 
        .CLK(n2067), .Q(\mem3[82][30] ), .QN(n29034) );
  SDFFX1 \mem3_reg[82][29]  ( .D(n13121), .SI(\mem3[82][28] ), .SE(test_se), 
        .CLK(n2067), .Q(\mem3[82][29] ), .QN(n29035) );
  SDFFX1 \mem3_reg[82][28]  ( .D(n13120), .SI(\mem3[82][27] ), .SE(test_se), 
        .CLK(n2067), .Q(\mem3[82][28] ), .QN(n29036) );
  SDFFX1 \mem3_reg[82][27]  ( .D(n13119), .SI(\mem3[82][26] ), .SE(test_se), 
        .CLK(n2067), .Q(\mem3[82][27] ), .QN(n29037) );
  SDFFX1 \mem3_reg[82][26]  ( .D(n13118), .SI(\mem3[82][25] ), .SE(test_se), 
        .CLK(n2067), .Q(\mem3[82][26] ), .QN(n29038) );
  SDFFX1 \mem3_reg[82][25]  ( .D(n13117), .SI(\mem3[82][24] ), .SE(test_se), 
        .CLK(n2067), .Q(\mem3[82][25] ), .QN(n29039) );
  SDFFX1 \mem3_reg[82][24]  ( .D(n13116), .SI(\mem3[81][31] ), .SE(test_se), 
        .CLK(n2067), .Q(\mem3[82][24] ), .QN(n29040) );
  SDFFX1 \mem3_reg[81][31]  ( .D(n13115), .SI(\mem3[81][30] ), .SE(test_se), 
        .CLK(n2067), .Q(\mem3[81][31] ), .QN(n29041) );
  SDFFX1 \mem3_reg[81][30]  ( .D(n13114), .SI(\mem3[81][29] ), .SE(test_se), 
        .CLK(n2067), .Q(\mem3[81][30] ), .QN(n29042) );
  SDFFX1 \mem3_reg[81][29]  ( .D(n13113), .SI(\mem3[81][28] ), .SE(test_se), 
        .CLK(n2067), .Q(\mem3[81][29] ), .QN(n29043) );
  SDFFX1 \mem3_reg[81][28]  ( .D(n13112), .SI(\mem3[81][27] ), .SE(test_se), 
        .CLK(n2067), .Q(\mem3[81][28] ), .QN(n29044) );
  SDFFX1 \mem3_reg[81][27]  ( .D(n13111), .SI(\mem3[81][26] ), .SE(test_se), 
        .CLK(n2068), .Q(\mem3[81][27] ), .QN(n29045) );
  SDFFX1 \mem3_reg[81][26]  ( .D(n13110), .SI(\mem3[81][25] ), .SE(test_se), 
        .CLK(n2068), .Q(\mem3[81][26] ), .QN(n29046) );
  SDFFX1 \mem3_reg[81][25]  ( .D(n13109), .SI(\mem3[81][24] ), .SE(test_se), 
        .CLK(n2068), .Q(\mem3[81][25] ), .QN(n29047) );
  SDFFX1 \mem3_reg[81][24]  ( .D(n13108), .SI(\mem3[80][31] ), .SE(test_se), 
        .CLK(n2068), .Q(\mem3[81][24] ), .QN(n29048) );
  SDFFX1 \mem3_reg[80][31]  ( .D(n13107), .SI(\mem3[80][30] ), .SE(test_se), 
        .CLK(n2068), .Q(\mem3[80][31] ), .QN(n29049) );
  SDFFX1 \mem3_reg[80][30]  ( .D(n13106), .SI(\mem3[80][29] ), .SE(test_se), 
        .CLK(n2068), .Q(\mem3[80][30] ), .QN(n29050) );
  SDFFX1 \mem3_reg[80][29]  ( .D(n13105), .SI(\mem3[80][28] ), .SE(test_se), 
        .CLK(n2068), .Q(\mem3[80][29] ), .QN(n29051) );
  SDFFX1 \mem3_reg[80][28]  ( .D(n13104), .SI(\mem3[80][27] ), .SE(test_se), 
        .CLK(n2068), .Q(\mem3[80][28] ), .QN(n29052) );
  SDFFX1 \mem3_reg[80][27]  ( .D(n13103), .SI(\mem3[80][26] ), .SE(test_se), 
        .CLK(n2068), .Q(\mem3[80][27] ), .QN(n29053) );
  SDFFX1 \mem3_reg[80][26]  ( .D(n13102), .SI(\mem3[80][25] ), .SE(test_se), 
        .CLK(n2068), .Q(\mem3[80][26] ), .QN(n29054) );
  SDFFX1 \mem3_reg[80][25]  ( .D(n13101), .SI(\mem3[80][24] ), .SE(test_se), 
        .CLK(n2068), .Q(\mem3[80][25] ), .QN(n29055) );
  SDFFX1 \mem3_reg[80][24]  ( .D(n13100), .SI(\mem3[79][31] ), .SE(test_se), 
        .CLK(n2068), .Q(\mem3[80][24] ), .QN(n29056) );
  SDFFX1 \mem3_reg[79][31]  ( .D(n13099), .SI(\mem3[79][30] ), .SE(test_se), 
        .CLK(n2071), .Q(\mem3[79][31] ), .QN(n29057) );
  SDFFX1 \mem3_reg[79][30]  ( .D(n13098), .SI(\mem3[79][29] ), .SE(test_se), 
        .CLK(n2071), .Q(\mem3[79][30] ), .QN(n29058) );
  SDFFX1 \mem3_reg[79][29]  ( .D(n13097), .SI(\mem3[79][28] ), .SE(test_se), 
        .CLK(n2071), .Q(\mem3[79][29] ), .QN(n29059) );
  SDFFX1 \mem3_reg[79][28]  ( .D(n13096), .SI(\mem3[79][27] ), .SE(test_se), 
        .CLK(n2071), .Q(\mem3[79][28] ), .QN(n29060) );
  SDFFX1 \mem3_reg[79][27]  ( .D(n13095), .SI(\mem3[79][26] ), .SE(test_se), 
        .CLK(n2071), .Q(\mem3[79][27] ), .QN(n29061) );
  SDFFX1 \mem3_reg[79][26]  ( .D(n13094), .SI(\mem3[79][25] ), .SE(test_se), 
        .CLK(n2072), .Q(\mem3[79][26] ), .QN(n29062) );
  SDFFX1 \mem3_reg[79][25]  ( .D(n13093), .SI(\mem3[79][24] ), .SE(test_se), 
        .CLK(n2072), .Q(\mem3[79][25] ), .QN(n29063) );
  SDFFX1 \mem3_reg[79][24]  ( .D(n13092), .SI(\mem3[78][31] ), .SE(test_se), 
        .CLK(n2072), .Q(\mem3[79][24] ), .QN(n29064) );
  SDFFX1 \mem3_reg[78][31]  ( .D(n13091), .SI(\mem3[78][30] ), .SE(test_se), 
        .CLK(n2073), .Q(\mem3[78][31] ), .QN(n29065) );
  SDFFX1 \mem3_reg[78][30]  ( .D(n13090), .SI(\mem3[78][29] ), .SE(test_se), 
        .CLK(n2073), .Q(\mem3[78][30] ), .QN(n29066) );
  SDFFX1 \mem3_reg[78][29]  ( .D(n13089), .SI(\mem3[78][28] ), .SE(test_se), 
        .CLK(n2073), .Q(\mem3[78][29] ), .QN(n29067) );
  SDFFX1 \mem3_reg[78][28]  ( .D(n13088), .SI(\mem3[78][27] ), .SE(test_se), 
        .CLK(n2073), .Q(\mem3[78][28] ), .QN(n29068) );
  SDFFX1 \mem3_reg[78][27]  ( .D(n13087), .SI(\mem3[78][26] ), .SE(test_se), 
        .CLK(n2073), .Q(\mem3[78][27] ), .QN(n29069) );
  SDFFX1 \mem3_reg[78][26]  ( .D(n13086), .SI(\mem3[78][25] ), .SE(test_se), 
        .CLK(n2074), .Q(\mem3[78][26] ), .QN(n29070) );
  SDFFX1 \mem3_reg[78][25]  ( .D(n13085), .SI(\mem3[78][24] ), .SE(test_se), 
        .CLK(n2074), .Q(\mem3[78][25] ), .QN(n29071) );
  SDFFX1 \mem3_reg[78][24]  ( .D(n13084), .SI(\mem3[77][31] ), .SE(test_se), 
        .CLK(n2074), .Q(\mem3[78][24] ), .QN(n29072) );
  SDFFX1 \mem3_reg[77][31]  ( .D(n13083), .SI(\mem3[77][30] ), .SE(test_se), 
        .CLK(n2074), .Q(\mem3[77][31] ), .QN(n29073) );
  SDFFX1 \mem3_reg[77][30]  ( .D(n13082), .SI(test_si7), .SE(test_se), .CLK(
        n2074), .Q(\mem3[77][30] ), .QN(n29074) );
  SDFFX1 \mem3_reg[77][29]  ( .D(n13081), .SI(\mem3[77][28] ), .SE(test_se), 
        .CLK(n1840), .Q(\mem3[77][29] ), .QN(n29075) );
  SDFFX1 \mem3_reg[77][28]  ( .D(n13080), .SI(\mem3[77][27] ), .SE(test_se), 
        .CLK(n1840), .Q(\mem3[77][28] ), .QN(n29076) );
  SDFFX1 \mem3_reg[77][27]  ( .D(n13079), .SI(\mem3[77][26] ), .SE(test_se), 
        .CLK(n1840), .Q(\mem3[77][27] ), .QN(n29077) );
  SDFFX1 \mem3_reg[77][26]  ( .D(n13078), .SI(\mem3[77][25] ), .SE(test_se), 
        .CLK(n1841), .Q(\mem3[77][26] ), .QN(n29078) );
  SDFFX1 \mem3_reg[77][25]  ( .D(n13077), .SI(\mem3[77][24] ), .SE(test_se), 
        .CLK(n1841), .Q(\mem3[77][25] ), .QN(n29079) );
  SDFFX1 \mem3_reg[77][24]  ( .D(n13076), .SI(\mem3[76][31] ), .SE(test_se), 
        .CLK(n1841), .Q(\mem3[77][24] ), .QN(n29080) );
  SDFFX1 \mem3_reg[76][31]  ( .D(n13075), .SI(\mem3[76][30] ), .SE(test_se), 
        .CLK(n1841), .Q(\mem3[76][31] ), .QN(n29081) );
  SDFFX1 \mem3_reg[76][30]  ( .D(n13074), .SI(\mem3[76][29] ), .SE(test_se), 
        .CLK(n1841), .Q(\mem3[76][30] ), .QN(n29082) );
  SDFFX1 \mem3_reg[76][29]  ( .D(n13073), .SI(\mem3[76][28] ), .SE(test_se), 
        .CLK(n1841), .Q(\mem3[76][29] ), .QN(n29083) );
  SDFFX1 \mem3_reg[76][28]  ( .D(n13072), .SI(\mem3[76][27] ), .SE(test_se), 
        .CLK(n1841), .Q(\mem3[76][28] ), .QN(n29084) );
  SDFFX1 \mem3_reg[76][27]  ( .D(n13071), .SI(\mem3[76][26] ), .SE(test_se), 
        .CLK(n1841), .Q(\mem3[76][27] ), .QN(n29085) );
  SDFFX1 \mem3_reg[76][26]  ( .D(n13070), .SI(\mem3[76][25] ), .SE(test_se), 
        .CLK(n1841), .Q(\mem3[76][26] ), .QN(n29086) );
  SDFFX1 \mem3_reg[76][25]  ( .D(n13069), .SI(\mem3[76][24] ), .SE(test_se), 
        .CLK(n1841), .Q(\mem3[76][25] ), .QN(n29087) );
  SDFFX1 \mem3_reg[76][24]  ( .D(n13068), .SI(\mem3[75][31] ), .SE(test_se), 
        .CLK(n1841), .Q(\mem3[76][24] ), .QN(n29088) );
  SDFFX1 \mem3_reg[75][31]  ( .D(n13067), .SI(\mem3[75][30] ), .SE(test_se), 
        .CLK(n1841), .Q(\mem3[75][31] ), .QN(n29089) );
  SDFFX1 \mem3_reg[75][30]  ( .D(n13066), .SI(\mem3[75][29] ), .SE(test_se), 
        .CLK(n1842), .Q(\mem3[75][30] ), .QN(n29090) );
  SDFFX1 \mem3_reg[75][29]  ( .D(n13065), .SI(\mem3[75][28] ), .SE(test_se), 
        .CLK(n1842), .Q(\mem3[75][29] ), .QN(n29091) );
  SDFFX1 \mem3_reg[75][28]  ( .D(n13064), .SI(\mem3[75][27] ), .SE(test_se), 
        .CLK(n1842), .Q(\mem3[75][28] ), .QN(n29092) );
  SDFFX1 \mem3_reg[75][27]  ( .D(n13063), .SI(\mem3[75][26] ), .SE(test_se), 
        .CLK(n1842), .Q(\mem3[75][27] ), .QN(n29093) );
  SDFFX1 \mem3_reg[75][26]  ( .D(n13062), .SI(\mem3[75][25] ), .SE(test_se), 
        .CLK(n1842), .Q(\mem3[75][26] ), .QN(n29094) );
  SDFFX1 \mem3_reg[75][25]  ( .D(n13061), .SI(\mem3[75][24] ), .SE(test_se), 
        .CLK(n1842), .Q(\mem3[75][25] ), .QN(n29095) );
  SDFFX1 \mem3_reg[75][24]  ( .D(n13060), .SI(\mem3[74][31] ), .SE(test_se), 
        .CLK(n1842), .Q(\mem3[75][24] ), .QN(n29096) );
  SDFFX1 \mem3_reg[74][31]  ( .D(n13059), .SI(\mem3[74][30] ), .SE(test_se), 
        .CLK(n1842), .Q(\mem3[74][31] ), .QN(n29097) );
  SDFFX1 \mem3_reg[74][30]  ( .D(n13058), .SI(\mem3[74][29] ), .SE(test_se), 
        .CLK(n1842), .Q(\mem3[74][30] ), .QN(n29098) );
  SDFFX1 \mem3_reg[74][29]  ( .D(n13057), .SI(\mem3[74][28] ), .SE(test_se), 
        .CLK(n1842), .Q(\mem3[74][29] ), .QN(n29099) );
  SDFFX1 \mem3_reg[74][28]  ( .D(n13056), .SI(\mem3[74][27] ), .SE(test_se), 
        .CLK(n1842), .Q(\mem3[74][28] ), .QN(n29100) );
  SDFFX1 \mem3_reg[74][27]  ( .D(n13055), .SI(\mem3[74][26] ), .SE(test_se), 
        .CLK(n1842), .Q(\mem3[74][27] ), .QN(n29101) );
  SDFFX1 \mem3_reg[74][26]  ( .D(n13054), .SI(\mem3[74][25] ), .SE(test_se), 
        .CLK(n1843), .Q(\mem3[74][26] ), .QN(n29102) );
  SDFFX1 \mem3_reg[74][25]  ( .D(n13053), .SI(\mem3[74][24] ), .SE(test_se), 
        .CLK(n1843), .Q(\mem3[74][25] ), .QN(n29103) );
  SDFFX1 \mem3_reg[74][24]  ( .D(n13052), .SI(\mem3[73][31] ), .SE(test_se), 
        .CLK(n1843), .Q(\mem3[74][24] ), .QN(n29104) );
  SDFFX1 \mem3_reg[73][31]  ( .D(n13051), .SI(\mem3[73][30] ), .SE(test_se), 
        .CLK(n1843), .Q(\mem3[73][31] ), .QN(n29105) );
  SDFFX1 \mem3_reg[73][30]  ( .D(n13050), .SI(\mem3[73][29] ), .SE(test_se), 
        .CLK(n1843), .Q(\mem3[73][30] ), .QN(n29106) );
  SDFFX1 \mem3_reg[73][29]  ( .D(n13049), .SI(\mem3[73][28] ), .SE(test_se), 
        .CLK(n1843), .Q(\mem3[73][29] ), .QN(n29107) );
  SDFFX1 \mem3_reg[73][28]  ( .D(n13048), .SI(\mem3[73][27] ), .SE(test_se), 
        .CLK(n1843), .Q(\mem3[73][28] ), .QN(n29108) );
  SDFFX1 \mem3_reg[73][27]  ( .D(n13047), .SI(\mem3[73][26] ), .SE(test_se), 
        .CLK(n1843), .Q(\mem3[73][27] ), .QN(n29109) );
  SDFFX1 \mem3_reg[73][26]  ( .D(n13046), .SI(\mem3[73][25] ), .SE(test_se), 
        .CLK(n1843), .Q(\mem3[73][26] ), .QN(n29110) );
  SDFFX1 \mem3_reg[73][25]  ( .D(n13045), .SI(\mem3[73][24] ), .SE(test_se), 
        .CLK(n1843), .Q(\mem3[73][25] ), .QN(n29111) );
  SDFFX1 \mem3_reg[73][24]  ( .D(n13044), .SI(\mem3[72][31] ), .SE(test_se), 
        .CLK(n1843), .Q(\mem3[73][24] ), .QN(n29112) );
  SDFFX1 \mem3_reg[72][31]  ( .D(n13043), .SI(\mem3[72][30] ), .SE(test_se), 
        .CLK(n1843), .Q(\mem3[72][31] ), .QN(n29113) );
  SDFFX1 \mem3_reg[72][30]  ( .D(n13042), .SI(\mem3[72][29] ), .SE(test_se), 
        .CLK(n1844), .Q(\mem3[72][30] ), .QN(n29114) );
  SDFFX1 \mem3_reg[72][29]  ( .D(n13041), .SI(\mem3[72][28] ), .SE(test_se), 
        .CLK(n1844), .Q(\mem3[72][29] ), .QN(n29115) );
  SDFFX1 \mem3_reg[72][28]  ( .D(n13040), .SI(\mem3[72][27] ), .SE(test_se), 
        .CLK(n1844), .Q(\mem3[72][28] ), .QN(n29116) );
  SDFFX1 \mem3_reg[72][27]  ( .D(n13039), .SI(\mem3[72][26] ), .SE(test_se), 
        .CLK(n1844), .Q(\mem3[72][27] ), .QN(n29117) );
  SDFFX1 \mem3_reg[72][26]  ( .D(n13038), .SI(\mem3[72][25] ), .SE(test_se), 
        .CLK(n1844), .Q(\mem3[72][26] ), .QN(n29118) );
  SDFFX1 \mem3_reg[72][25]  ( .D(n13037), .SI(\mem3[72][24] ), .SE(test_se), 
        .CLK(n1844), .Q(\mem3[72][25] ), .QN(n29119) );
  SDFFX1 \mem3_reg[72][24]  ( .D(n13036), .SI(\mem3[71][31] ), .SE(test_se), 
        .CLK(n1844), .Q(\mem3[72][24] ), .QN(n29120) );
  SDFFX1 \mem3_reg[71][31]  ( .D(n13035), .SI(\mem3[71][30] ), .SE(test_se), 
        .CLK(n1844), .Q(\mem3[71][31] ), .QN(n29121) );
  SDFFX1 \mem3_reg[71][30]  ( .D(n13034), .SI(\mem3[71][29] ), .SE(test_se), 
        .CLK(n1844), .Q(\mem3[71][30] ), .QN(n29122) );
  SDFFX1 \mem3_reg[71][29]  ( .D(n13033), .SI(\mem3[71][28] ), .SE(test_se), 
        .CLK(n1844), .Q(\mem3[71][29] ), .QN(n29123) );
  SDFFX1 \mem3_reg[71][28]  ( .D(n13032), .SI(\mem3[71][27] ), .SE(test_se), 
        .CLK(n1844), .Q(\mem3[71][28] ), .QN(n29124) );
  SDFFX1 \mem3_reg[71][27]  ( .D(n13031), .SI(\mem3[71][26] ), .SE(test_se), 
        .CLK(n1844), .Q(\mem3[71][27] ), .QN(n29125) );
  SDFFX1 \mem3_reg[71][26]  ( .D(n13030), .SI(\mem3[71][25] ), .SE(test_se), 
        .CLK(n1845), .Q(\mem3[71][26] ), .QN(n29126) );
  SDFFX1 \mem3_reg[71][25]  ( .D(n13029), .SI(\mem3[71][24] ), .SE(test_se), 
        .CLK(n1845), .Q(\mem3[71][25] ), .QN(n29127) );
  SDFFX1 \mem3_reg[71][24]  ( .D(n13028), .SI(\mem3[70][31] ), .SE(test_se), 
        .CLK(n1845), .Q(\mem3[71][24] ), .QN(n29128) );
  SDFFX1 \mem3_reg[70][31]  ( .D(n13027), .SI(\mem3[70][30] ), .SE(test_se), 
        .CLK(n1845), .Q(\mem3[70][31] ), .QN(n29129) );
  SDFFX1 \mem3_reg[70][30]  ( .D(n13026), .SI(\mem3[70][29] ), .SE(test_se), 
        .CLK(n1845), .Q(\mem3[70][30] ), .QN(n29130) );
  SDFFX1 \mem3_reg[70][29]  ( .D(n13025), .SI(\mem3[70][28] ), .SE(test_se), 
        .CLK(n1845), .Q(\mem3[70][29] ), .QN(n29131) );
  SDFFX1 \mem3_reg[70][28]  ( .D(n13024), .SI(\mem3[70][27] ), .SE(test_se), 
        .CLK(n1845), .Q(\mem3[70][28] ), .QN(n29132) );
  SDFFX1 \mem3_reg[70][27]  ( .D(n13023), .SI(\mem3[70][26] ), .SE(test_se), 
        .CLK(n1845), .Q(\mem3[70][27] ), .QN(n29133) );
  SDFFX1 \mem3_reg[70][26]  ( .D(n13022), .SI(\mem3[70][25] ), .SE(test_se), 
        .CLK(n1845), .Q(\mem3[70][26] ), .QN(n29134) );
  SDFFX1 \mem3_reg[70][25]  ( .D(n13021), .SI(\mem3[70][24] ), .SE(test_se), 
        .CLK(n1845), .Q(\mem3[70][25] ), .QN(n29135) );
  SDFFX1 \mem3_reg[70][24]  ( .D(n13020), .SI(\mem3[69][31] ), .SE(test_se), 
        .CLK(n1845), .Q(\mem3[70][24] ), .QN(n29136) );
  SDFFX1 \mem3_reg[69][31]  ( .D(n13019), .SI(\mem3[69][30] ), .SE(test_se), 
        .CLK(n1845), .Q(\mem3[69][31] ), .QN(n29137) );
  SDFFX1 \mem3_reg[69][30]  ( .D(n13018), .SI(\mem3[69][29] ), .SE(test_se), 
        .CLK(n1846), .Q(\mem3[69][30] ), .QN(n29138) );
  SDFFX1 \mem3_reg[69][29]  ( .D(n13017), .SI(\mem3[69][28] ), .SE(test_se), 
        .CLK(n1846), .Q(\mem3[69][29] ), .QN(n29139) );
  SDFFX1 \mem3_reg[69][28]  ( .D(n13016), .SI(\mem3[69][27] ), .SE(test_se), 
        .CLK(n1846), .Q(\mem3[69][28] ), .QN(n29140) );
  SDFFX1 \mem3_reg[69][27]  ( .D(n13015), .SI(\mem3[69][26] ), .SE(test_se), 
        .CLK(n1846), .Q(\mem3[69][27] ), .QN(n29141) );
  SDFFX1 \mem3_reg[69][26]  ( .D(n13014), .SI(\mem3[69][25] ), .SE(test_se), 
        .CLK(n1846), .Q(\mem3[69][26] ), .QN(n29142) );
  SDFFX1 \mem3_reg[69][25]  ( .D(n13013), .SI(\mem3[69][24] ), .SE(test_se), 
        .CLK(n1846), .Q(\mem3[69][25] ), .QN(n29143) );
  SDFFX1 \mem3_reg[69][24]  ( .D(n13012), .SI(\mem3[68][31] ), .SE(test_se), 
        .CLK(n1846), .Q(\mem3[69][24] ), .QN(n29144) );
  SDFFX1 \mem3_reg[68][31]  ( .D(n13011), .SI(\mem3[68][30] ), .SE(test_se), 
        .CLK(n1846), .Q(\mem3[68][31] ), .QN(n29145) );
  SDFFX1 \mem3_reg[68][30]  ( .D(n13010), .SI(\mem3[68][29] ), .SE(test_se), 
        .CLK(n1846), .Q(\mem3[68][30] ), .QN(n29146) );
  SDFFX1 \mem3_reg[68][29]  ( .D(n13009), .SI(\mem3[68][28] ), .SE(test_se), 
        .CLK(n1846), .Q(\mem3[68][29] ), .QN(n29147) );
  SDFFX1 \mem3_reg[68][28]  ( .D(n13008), .SI(\mem3[68][27] ), .SE(test_se), 
        .CLK(n1846), .Q(\mem3[68][28] ), .QN(n29148) );
  SDFFX1 \mem3_reg[68][27]  ( .D(n13007), .SI(\mem3[68][26] ), .SE(test_se), 
        .CLK(n1846), .Q(\mem3[68][27] ), .QN(n29149) );
  SDFFX1 \mem3_reg[68][26]  ( .D(n13006), .SI(\mem3[68][25] ), .SE(test_se), 
        .CLK(n1847), .Q(\mem3[68][26] ), .QN(n29150) );
  SDFFX1 \mem3_reg[68][25]  ( .D(n13005), .SI(\mem3[68][24] ), .SE(test_se), 
        .CLK(n1847), .Q(\mem3[68][25] ), .QN(n29151) );
  SDFFX1 \mem3_reg[68][24]  ( .D(n13004), .SI(\mem3[67][31] ), .SE(test_se), 
        .CLK(n1847), .Q(\mem3[68][24] ), .QN(n29152) );
  SDFFX1 \mem3_reg[67][31]  ( .D(n13003), .SI(\mem3[67][30] ), .SE(test_se), 
        .CLK(n1847), .Q(\mem3[67][31] ), .QN(n29153) );
  SDFFX1 \mem3_reg[67][30]  ( .D(n13002), .SI(\mem3[67][29] ), .SE(test_se), 
        .CLK(n1847), .Q(\mem3[67][30] ), .QN(n29154) );
  SDFFX1 \mem3_reg[67][29]  ( .D(n13001), .SI(\mem3[67][28] ), .SE(test_se), 
        .CLK(n1847), .Q(\mem3[67][29] ), .QN(n29155) );
  SDFFX1 \mem3_reg[67][28]  ( .D(n13000), .SI(\mem3[67][27] ), .SE(test_se), 
        .CLK(n1847), .Q(\mem3[67][28] ), .QN(n29156) );
  SDFFX1 \mem3_reg[67][27]  ( .D(n12999), .SI(\mem3[67][26] ), .SE(test_se), 
        .CLK(n1847), .Q(\mem3[67][27] ), .QN(n29157) );
  SDFFX1 \mem3_reg[67][26]  ( .D(n12998), .SI(\mem3[67][25] ), .SE(test_se), 
        .CLK(n1847), .Q(\mem3[67][26] ), .QN(n29158) );
  SDFFX1 \mem3_reg[67][25]  ( .D(n12997), .SI(\mem3[67][24] ), .SE(test_se), 
        .CLK(n1847), .Q(\mem3[67][25] ), .QN(n29159) );
  SDFFX1 \mem3_reg[67][24]  ( .D(n12996), .SI(\mem3[66][31] ), .SE(test_se), 
        .CLK(n1847), .Q(\mem3[67][24] ), .QN(n29160) );
  SDFFX1 \mem3_reg[66][31]  ( .D(n12995), .SI(\mem3[66][30] ), .SE(test_se), 
        .CLK(n1847), .Q(\mem3[66][31] ), .QN(n29161) );
  SDFFX1 \mem3_reg[66][30]  ( .D(n12994), .SI(\mem3[66][29] ), .SE(test_se), 
        .CLK(n1848), .Q(\mem3[66][30] ), .QN(n29162) );
  SDFFX1 \mem3_reg[66][29]  ( .D(n12993), .SI(\mem3[66][28] ), .SE(test_se), 
        .CLK(n1848), .Q(\mem3[66][29] ), .QN(n29163) );
  SDFFX1 \mem3_reg[66][28]  ( .D(n12992), .SI(\mem3[66][27] ), .SE(test_se), 
        .CLK(n1848), .Q(\mem3[66][28] ), .QN(n29164) );
  SDFFX1 \mem3_reg[66][27]  ( .D(n12991), .SI(\mem3[66][26] ), .SE(test_se), 
        .CLK(n1848), .Q(\mem3[66][27] ), .QN(n29165) );
  SDFFX1 \mem3_reg[66][26]  ( .D(n12990), .SI(\mem3[66][25] ), .SE(test_se), 
        .CLK(n1848), .Q(\mem3[66][26] ), .QN(n29166) );
  SDFFX1 \mem3_reg[66][25]  ( .D(n12989), .SI(\mem3[66][24] ), .SE(test_se), 
        .CLK(n1848), .Q(\mem3[66][25] ), .QN(n29167) );
  SDFFX1 \mem3_reg[66][24]  ( .D(n12988), .SI(\mem3[65][31] ), .SE(test_se), 
        .CLK(n1848), .Q(\mem3[66][24] ), .QN(n29168) );
  SDFFX1 \mem3_reg[65][31]  ( .D(n12987), .SI(\mem3[65][30] ), .SE(test_se), 
        .CLK(n1848), .Q(\mem3[65][31] ), .QN(n29169) );
  SDFFX1 \mem3_reg[65][30]  ( .D(n12986), .SI(\mem3[65][29] ), .SE(test_se), 
        .CLK(n1848), .Q(\mem3[65][30] ), .QN(n29170) );
  SDFFX1 \mem3_reg[65][29]  ( .D(n12985), .SI(\mem3[65][28] ), .SE(test_se), 
        .CLK(n1848), .Q(\mem3[65][29] ), .QN(n29171) );
  SDFFX1 \mem3_reg[65][28]  ( .D(n12984), .SI(\mem3[65][27] ), .SE(test_se), 
        .CLK(n1848), .Q(\mem3[65][28] ), .QN(n29172) );
  SDFFX1 \mem3_reg[65][27]  ( .D(n12983), .SI(\mem3[65][26] ), .SE(test_se), 
        .CLK(n1848), .Q(\mem3[65][27] ), .QN(n29173) );
  SDFFX1 \mem3_reg[65][26]  ( .D(n12982), .SI(\mem3[65][25] ), .SE(test_se), 
        .CLK(n1849), .Q(\mem3[65][26] ), .QN(n29174) );
  SDFFX1 \mem3_reg[65][25]  ( .D(n12981), .SI(\mem3[65][24] ), .SE(test_se), 
        .CLK(n1849), .Q(\mem3[65][25] ), .QN(n29175) );
  SDFFX1 \mem3_reg[65][24]  ( .D(n12980), .SI(\mem3[64][31] ), .SE(test_se), 
        .CLK(n1849), .Q(\mem3[65][24] ), .QN(n29176) );
  SDFFX1 \mem3_reg[64][31]  ( .D(n12979), .SI(\mem3[64][30] ), .SE(test_se), 
        .CLK(n1849), .Q(\mem3[64][31] ), .QN(n29177) );
  SDFFX1 \mem3_reg[64][30]  ( .D(n12978), .SI(\mem3[64][29] ), .SE(test_se), 
        .CLK(n1849), .Q(\mem3[64][30] ), .QN(n29178) );
  SDFFX1 \mem3_reg[64][29]  ( .D(n12977), .SI(\mem3[64][28] ), .SE(test_se), 
        .CLK(n1849), .Q(\mem3[64][29] ), .QN(n29179) );
  SDFFX1 \mem3_reg[64][28]  ( .D(n12976), .SI(\mem3[64][27] ), .SE(test_se), 
        .CLK(n1849), .Q(\mem3[64][28] ), .QN(n29180) );
  SDFFX1 \mem3_reg[64][27]  ( .D(n12975), .SI(\mem3[64][26] ), .SE(test_se), 
        .CLK(n1849), .Q(\mem3[64][27] ), .QN(n29181) );
  SDFFX1 \mem3_reg[64][26]  ( .D(n12974), .SI(\mem3[64][25] ), .SE(test_se), 
        .CLK(n1849), .Q(\mem3[64][26] ), .QN(n29182) );
  SDFFX1 \mem3_reg[64][25]  ( .D(n12973), .SI(\mem3[64][24] ), .SE(test_se), 
        .CLK(n1849), .Q(\mem3[64][25] ), .QN(n29183) );
  SDFFX1 \mem3_reg[64][24]  ( .D(n12972), .SI(\mem3[63][31] ), .SE(test_se), 
        .CLK(n1849), .Q(\mem3[64][24] ), .QN(n29184) );
  SDFFX1 \mem3_reg[63][31]  ( .D(n12971), .SI(\mem3[63][30] ), .SE(test_se), 
        .CLK(n1849), .Q(\mem3[63][31] ), .QN(n29185) );
  SDFFX1 \mem3_reg[63][30]  ( .D(n12970), .SI(\mem3[63][29] ), .SE(test_se), 
        .CLK(n1850), .Q(\mem3[63][30] ), .QN(n29186) );
  SDFFX1 \mem3_reg[63][29]  ( .D(n12969), .SI(\mem3[63][28] ), .SE(test_se), 
        .CLK(n1850), .Q(\mem3[63][29] ), .QN(n29187) );
  SDFFX1 \mem3_reg[63][28]  ( .D(n12968), .SI(\mem3[63][27] ), .SE(test_se), 
        .CLK(n1850), .Q(\mem3[63][28] ), .QN(n29188) );
  SDFFX1 \mem3_reg[63][27]  ( .D(n12967), .SI(\mem3[63][26] ), .SE(test_se), 
        .CLK(n1850), .Q(\mem3[63][27] ), .QN(n29189) );
  SDFFX1 \mem3_reg[63][26]  ( .D(n12966), .SI(\mem3[63][25] ), .SE(test_se), 
        .CLK(n1850), .Q(\mem3[63][26] ), .QN(n29190) );
  SDFFX1 \mem3_reg[63][25]  ( .D(n12965), .SI(\mem3[63][24] ), .SE(test_se), 
        .CLK(n1850), .Q(\mem3[63][25] ), .QN(n29191) );
  SDFFX1 \mem3_reg[63][24]  ( .D(n12964), .SI(\mem3[62][31] ), .SE(test_se), 
        .CLK(n1850), .Q(\mem3[63][24] ), .QN(n29192) );
  SDFFX1 \mem3_reg[62][31]  ( .D(n12963), .SI(\mem3[62][30] ), .SE(test_se), 
        .CLK(n1850), .Q(\mem3[62][31] ), .QN(n29193) );
  SDFFX1 \mem3_reg[62][30]  ( .D(n12962), .SI(\mem3[62][29] ), .SE(test_se), 
        .CLK(n1850), .Q(\mem3[62][30] ), .QN(n29194) );
  SDFFX1 \mem3_reg[62][29]  ( .D(n12961), .SI(\mem3[62][28] ), .SE(test_se), 
        .CLK(n1850), .Q(\mem3[62][29] ), .QN(n29195) );
  SDFFX1 \mem3_reg[62][28]  ( .D(n12960), .SI(\mem3[62][27] ), .SE(test_se), 
        .CLK(n1850), .Q(\mem3[62][28] ), .QN(n29196) );
  SDFFX1 \mem3_reg[62][27]  ( .D(n12959), .SI(\mem3[62][26] ), .SE(test_se), 
        .CLK(n1850), .Q(\mem3[62][27] ), .QN(n29197) );
  SDFFX1 \mem3_reg[62][26]  ( .D(n12958), .SI(\mem3[62][25] ), .SE(test_se), 
        .CLK(n1851), .Q(\mem3[62][26] ), .QN(n29198) );
  SDFFX1 \mem3_reg[62][25]  ( .D(n12957), .SI(\mem3[62][24] ), .SE(test_se), 
        .CLK(n1851), .Q(\mem3[62][25] ), .QN(n29199) );
  SDFFX1 \mem3_reg[62][24]  ( .D(n12956), .SI(\mem3[61][31] ), .SE(test_se), 
        .CLK(n1851), .Q(\mem3[62][24] ), .QN(n29200) );
  SDFFX1 \mem3_reg[61][31]  ( .D(n12955), .SI(\mem3[61][30] ), .SE(test_se), 
        .CLK(n1851), .Q(\mem3[61][31] ), .QN(n29201) );
  SDFFX1 \mem3_reg[61][30]  ( .D(n12954), .SI(\mem3[61][29] ), .SE(test_se), 
        .CLK(n1851), .Q(\mem3[61][30] ), .QN(n29202) );
  SDFFX1 \mem3_reg[61][29]  ( .D(n12953), .SI(\mem3[61][28] ), .SE(test_se), 
        .CLK(n1851), .Q(\mem3[61][29] ), .QN(n29203) );
  SDFFX1 \mem3_reg[61][28]  ( .D(n12952), .SI(\mem3[61][27] ), .SE(test_se), 
        .CLK(n1851), .Q(\mem3[61][28] ), .QN(n29204) );
  SDFFX1 \mem3_reg[61][27]  ( .D(n12951), .SI(\mem3[61][26] ), .SE(test_se), 
        .CLK(n1851), .Q(\mem3[61][27] ), .QN(n29205) );
  SDFFX1 \mem3_reg[61][26]  ( .D(n12950), .SI(\mem3[61][25] ), .SE(test_se), 
        .CLK(n1851), .Q(\mem3[61][26] ), .QN(n29206) );
  SDFFX1 \mem3_reg[61][25]  ( .D(n12949), .SI(\mem3[61][24] ), .SE(test_se), 
        .CLK(n1851), .Q(\mem3[61][25] ), .QN(n29207) );
  SDFFX1 \mem3_reg[61][24]  ( .D(n12948), .SI(\mem3[60][31] ), .SE(test_se), 
        .CLK(n1851), .Q(\mem3[61][24] ), .QN(n29208) );
  SDFFX1 \mem3_reg[60][31]  ( .D(n12947), .SI(\mem3[60][30] ), .SE(test_se), 
        .CLK(n1851), .Q(\mem3[60][31] ), .QN(n29209) );
  SDFFX1 \mem3_reg[60][30]  ( .D(n12946), .SI(\mem3[60][29] ), .SE(test_se), 
        .CLK(n1852), .Q(\mem3[60][30] ), .QN(n29210) );
  SDFFX1 \mem3_reg[60][29]  ( .D(n12945), .SI(\mem3[60][28] ), .SE(test_se), 
        .CLK(n1852), .Q(\mem3[60][29] ), .QN(n29211) );
  SDFFX1 \mem3_reg[60][28]  ( .D(n12944), .SI(\mem3[60][27] ), .SE(test_se), 
        .CLK(n1852), .Q(\mem3[60][28] ), .QN(n29212) );
  SDFFX1 \mem3_reg[60][27]  ( .D(n12943), .SI(\mem3[60][26] ), .SE(test_se), 
        .CLK(n1852), .Q(\mem3[60][27] ), .QN(n29213) );
  SDFFX1 \mem3_reg[60][26]  ( .D(n12942), .SI(\mem3[60][25] ), .SE(test_se), 
        .CLK(n1852), .Q(\mem3[60][26] ), .QN(n29214) );
  SDFFX1 \mem3_reg[60][25]  ( .D(n12941), .SI(\mem3[60][24] ), .SE(test_se), 
        .CLK(n1852), .Q(\mem3[60][25] ), .QN(n29215) );
  SDFFX1 \mem3_reg[60][24]  ( .D(n12940), .SI(\mem3[59][31] ), .SE(test_se), 
        .CLK(n1852), .Q(\mem3[60][24] ), .QN(n29216) );
  SDFFX1 \mem3_reg[59][31]  ( .D(n12939), .SI(\mem3[59][30] ), .SE(test_se), 
        .CLK(n1852), .Q(\mem3[59][31] ), .QN(n29217) );
  SDFFX1 \mem3_reg[59][30]  ( .D(n12938), .SI(\mem3[59][29] ), .SE(test_se), 
        .CLK(n1852), .Q(\mem3[59][30] ), .QN(n29218) );
  SDFFX1 \mem3_reg[59][29]  ( .D(n12937), .SI(\mem3[59][28] ), .SE(test_se), 
        .CLK(n1852), .Q(\mem3[59][29] ), .QN(n29219) );
  SDFFX1 \mem3_reg[59][28]  ( .D(n12936), .SI(\mem3[59][27] ), .SE(test_se), 
        .CLK(n1852), .Q(\mem3[59][28] ), .QN(n29220) );
  SDFFX1 \mem3_reg[59][27]  ( .D(n12935), .SI(\mem3[59][26] ), .SE(test_se), 
        .CLK(n1852), .Q(\mem3[59][27] ), .QN(n29221) );
  SDFFX1 \mem3_reg[59][26]  ( .D(n12934), .SI(\mem3[59][25] ), .SE(test_se), 
        .CLK(n1853), .Q(\mem3[59][26] ), .QN(n29222) );
  SDFFX1 \mem3_reg[59][25]  ( .D(n12933), .SI(\mem3[59][24] ), .SE(test_se), 
        .CLK(n1853), .Q(\mem3[59][25] ), .QN(n29223) );
  SDFFX1 \mem3_reg[59][24]  ( .D(n12932), .SI(\mem3[58][31] ), .SE(test_se), 
        .CLK(n1853), .Q(\mem3[59][24] ), .QN(n29224) );
  SDFFX1 \mem3_reg[58][31]  ( .D(n12931), .SI(\mem3[58][30] ), .SE(test_se), 
        .CLK(n1853), .Q(\mem3[58][31] ), .QN(n29225) );
  SDFFX1 \mem3_reg[58][30]  ( .D(n12930), .SI(\mem3[58][29] ), .SE(test_se), 
        .CLK(n1853), .Q(\mem3[58][30] ), .QN(n29226) );
  SDFFX1 \mem3_reg[58][29]  ( .D(n12929), .SI(\mem3[58][28] ), .SE(test_se), 
        .CLK(n1853), .Q(\mem3[58][29] ), .QN(n29227) );
  SDFFX1 \mem3_reg[58][28]  ( .D(n12928), .SI(\mem3[58][27] ), .SE(test_se), 
        .CLK(n1853), .Q(\mem3[58][28] ), .QN(n29228) );
  SDFFX1 \mem3_reg[58][27]  ( .D(n12927), .SI(\mem3[58][26] ), .SE(test_se), 
        .CLK(n1853), .Q(\mem3[58][27] ), .QN(n29229) );
  SDFFX1 \mem3_reg[58][26]  ( .D(n12926), .SI(\mem3[58][25] ), .SE(test_se), 
        .CLK(n1853), .Q(\mem3[58][26] ), .QN(n29230) );
  SDFFX1 \mem3_reg[58][25]  ( .D(n12925), .SI(\mem3[58][24] ), .SE(test_se), 
        .CLK(n1853), .Q(\mem3[58][25] ), .QN(n29231) );
  SDFFX1 \mem3_reg[58][24]  ( .D(n12924), .SI(\mem3[57][31] ), .SE(test_se), 
        .CLK(n1853), .Q(\mem3[58][24] ), .QN(n29232) );
  SDFFX1 \mem3_reg[57][31]  ( .D(n12923), .SI(\mem3[57][30] ), .SE(test_se), 
        .CLK(n1853), .Q(\mem3[57][31] ), .QN(n29233) );
  SDFFX1 \mem3_reg[57][30]  ( .D(n12922), .SI(\mem3[57][29] ), .SE(test_se), 
        .CLK(n1854), .Q(\mem3[57][30] ), .QN(n29234) );
  SDFFX1 \mem3_reg[57][29]  ( .D(n12921), .SI(\mem3[57][28] ), .SE(test_se), 
        .CLK(n1854), .Q(\mem3[57][29] ), .QN(n29235) );
  SDFFX1 \mem3_reg[57][28]  ( .D(n12920), .SI(\mem3[57][27] ), .SE(test_se), 
        .CLK(n1854), .Q(\mem3[57][28] ), .QN(n29236) );
  SDFFX1 \mem3_reg[57][27]  ( .D(n12919), .SI(\mem3[57][26] ), .SE(test_se), 
        .CLK(n1854), .Q(\mem3[57][27] ), .QN(n29237) );
  SDFFX1 \mem3_reg[57][26]  ( .D(n12918), .SI(\mem3[57][25] ), .SE(test_se), 
        .CLK(n1854), .Q(\mem3[57][26] ), .QN(n29238) );
  SDFFX1 \mem3_reg[57][25]  ( .D(n12917), .SI(\mem3[57][24] ), .SE(test_se), 
        .CLK(n1854), .Q(\mem3[57][25] ), .QN(n29239) );
  SDFFX1 \mem3_reg[57][24]  ( .D(n12916), .SI(\mem3[56][31] ), .SE(test_se), 
        .CLK(n1854), .Q(\mem3[57][24] ), .QN(n29240) );
  SDFFX1 \mem3_reg[56][31]  ( .D(n12915), .SI(\mem3[56][30] ), .SE(test_se), 
        .CLK(n1854), .Q(\mem3[56][31] ), .QN(n29241) );
  SDFFX1 \mem3_reg[56][30]  ( .D(n12914), .SI(\mem3[56][29] ), .SE(test_se), 
        .CLK(n1854), .Q(\mem3[56][30] ), .QN(n29242) );
  SDFFX1 \mem3_reg[56][29]  ( .D(n12913), .SI(\mem3[56][28] ), .SE(test_se), 
        .CLK(n1854), .Q(\mem3[56][29] ), .QN(n29243) );
  SDFFX1 \mem3_reg[56][28]  ( .D(n12912), .SI(\mem3[56][27] ), .SE(test_se), 
        .CLK(n1854), .Q(\mem3[56][28] ), .QN(n29244) );
  SDFFX1 \mem3_reg[56][27]  ( .D(n12911), .SI(\mem3[56][26] ), .SE(test_se), 
        .CLK(n1854), .Q(\mem3[56][27] ), .QN(n29245) );
  SDFFX1 \mem3_reg[56][26]  ( .D(n12910), .SI(\mem3[56][25] ), .SE(test_se), 
        .CLK(n1855), .Q(\mem3[56][26] ), .QN(n29246) );
  SDFFX1 \mem3_reg[56][25]  ( .D(n12909), .SI(\mem3[56][24] ), .SE(test_se), 
        .CLK(n1855), .Q(\mem3[56][25] ), .QN(n29247) );
  SDFFX1 \mem3_reg[56][24]  ( .D(n12908), .SI(\mem3[55][31] ), .SE(test_se), 
        .CLK(n1855), .Q(\mem3[56][24] ), .QN(n29248) );
  SDFFX1 \mem3_reg[55][31]  ( .D(n12907), .SI(\mem3[55][30] ), .SE(test_se), 
        .CLK(n1855), .Q(\mem3[55][31] ), .QN(n29249) );
  SDFFX1 \mem3_reg[55][30]  ( .D(n12906), .SI(\mem3[55][29] ), .SE(test_se), 
        .CLK(n1855), .Q(\mem3[55][30] ), .QN(n29250) );
  SDFFX1 \mem3_reg[55][29]  ( .D(n12905), .SI(\mem3[55][28] ), .SE(test_se), 
        .CLK(n1855), .Q(\mem3[55][29] ), .QN(n29251) );
  SDFFX1 \mem3_reg[55][28]  ( .D(n12904), .SI(\mem3[55][27] ), .SE(test_se), 
        .CLK(n1855), .Q(\mem3[55][28] ), .QN(n29252) );
  SDFFX1 \mem3_reg[55][27]  ( .D(n12903), .SI(\mem3[55][26] ), .SE(test_se), 
        .CLK(n1855), .Q(\mem3[55][27] ), .QN(n29253) );
  SDFFX1 \mem3_reg[55][26]  ( .D(n12902), .SI(\mem3[55][25] ), .SE(test_se), 
        .CLK(n1855), .Q(\mem3[55][26] ), .QN(n29254) );
  SDFFX1 \mem3_reg[55][25]  ( .D(n12901), .SI(\mem3[55][24] ), .SE(test_se), 
        .CLK(n1855), .Q(\mem3[55][25] ), .QN(n29255) );
  SDFFX1 \mem3_reg[55][24]  ( .D(n12900), .SI(\mem3[54][31] ), .SE(test_se), 
        .CLK(n1855), .Q(\mem3[55][24] ), .QN(n29256) );
  SDFFX1 \mem3_reg[54][31]  ( .D(n12899), .SI(\mem3[54][30] ), .SE(test_se), 
        .CLK(n1855), .Q(\mem3[54][31] ), .QN(n29257) );
  SDFFX1 \mem3_reg[54][30]  ( .D(n12898), .SI(\mem3[54][29] ), .SE(test_se), 
        .CLK(n1856), .Q(\mem3[54][30] ), .QN(n29258) );
  SDFFX1 \mem3_reg[54][29]  ( .D(n12897), .SI(\mem3[54][28] ), .SE(test_se), 
        .CLK(n1856), .Q(\mem3[54][29] ), .QN(n29259) );
  SDFFX1 \mem3_reg[54][28]  ( .D(n12896), .SI(\mem3[54][27] ), .SE(test_se), 
        .CLK(n1856), .Q(\mem3[54][28] ), .QN(n29260) );
  SDFFX1 \mem3_reg[54][27]  ( .D(n12895), .SI(\mem3[54][26] ), .SE(test_se), 
        .CLK(n1856), .Q(\mem3[54][27] ), .QN(n29261) );
  SDFFX1 \mem3_reg[54][26]  ( .D(n12894), .SI(\mem3[54][25] ), .SE(test_se), 
        .CLK(n1856), .Q(\mem3[54][26] ), .QN(n29262) );
  SDFFX1 \mem3_reg[54][25]  ( .D(n12893), .SI(\mem3[54][24] ), .SE(test_se), 
        .CLK(n1856), .Q(\mem3[54][25] ), .QN(n29263) );
  SDFFX1 \mem3_reg[54][24]  ( .D(n12892), .SI(\mem3[53][31] ), .SE(test_se), 
        .CLK(n1856), .Q(\mem3[54][24] ), .QN(n29264) );
  SDFFX1 \mem3_reg[53][31]  ( .D(n12891), .SI(\mem3[53][30] ), .SE(test_se), 
        .CLK(n1856), .Q(\mem3[53][31] ), .QN(n29265) );
  SDFFX1 \mem3_reg[53][30]  ( .D(n12890), .SI(\mem3[53][29] ), .SE(test_se), 
        .CLK(n1856), .Q(\mem3[53][30] ), .QN(n29266) );
  SDFFX1 \mem3_reg[53][29]  ( .D(n12889), .SI(\mem3[53][28] ), .SE(test_se), 
        .CLK(n1856), .Q(\mem3[53][29] ), .QN(n29267) );
  SDFFX1 \mem3_reg[53][28]  ( .D(n12888), .SI(\mem3[53][27] ), .SE(test_se), 
        .CLK(n1856), .Q(\mem3[53][28] ), .QN(n29268) );
  SDFFX1 \mem3_reg[53][27]  ( .D(n12887), .SI(\mem3[53][26] ), .SE(test_se), 
        .CLK(n1856), .Q(\mem3[53][27] ), .QN(n29269) );
  SDFFX1 \mem3_reg[53][26]  ( .D(n12886), .SI(\mem3[53][25] ), .SE(test_se), 
        .CLK(n1857), .Q(\mem3[53][26] ), .QN(n29270) );
  SDFFX1 \mem3_reg[53][25]  ( .D(n12885), .SI(\mem3[53][24] ), .SE(test_se), 
        .CLK(n1857), .Q(\mem3[53][25] ), .QN(n29271) );
  SDFFX1 \mem3_reg[53][24]  ( .D(n12884), .SI(\mem3[52][31] ), .SE(test_se), 
        .CLK(n1857), .Q(\mem3[53][24] ), .QN(n29272) );
  SDFFX1 \mem3_reg[52][31]  ( .D(n12883), .SI(\mem3[52][30] ), .SE(test_se), 
        .CLK(n1857), .Q(\mem3[52][31] ), .QN(n29273) );
  SDFFX1 \mem3_reg[52][30]  ( .D(n12882), .SI(\mem3[52][29] ), .SE(test_se), 
        .CLK(n1857), .Q(\mem3[52][30] ), .QN(n29274) );
  SDFFX1 \mem3_reg[52][29]  ( .D(n12881), .SI(\mem3[52][28] ), .SE(test_se), 
        .CLK(n1857), .Q(\mem3[52][29] ), .QN(n29275) );
  SDFFX1 \mem3_reg[52][28]  ( .D(n12880), .SI(\mem3[52][27] ), .SE(test_se), 
        .CLK(n1857), .Q(\mem3[52][28] ), .QN(n29276) );
  SDFFX1 \mem3_reg[52][27]  ( .D(n12879), .SI(\mem3[52][26] ), .SE(test_se), 
        .CLK(n1857), .Q(\mem3[52][27] ), .QN(n29277) );
  SDFFX1 \mem3_reg[52][26]  ( .D(n12878), .SI(\mem3[52][25] ), .SE(test_se), 
        .CLK(n1857), .Q(\mem3[52][26] ), .QN(n29278) );
  SDFFX1 \mem3_reg[52][25]  ( .D(n12877), .SI(\mem3[52][24] ), .SE(test_se), 
        .CLK(n1857), .Q(\mem3[52][25] ), .QN(n29279) );
  SDFFX1 \mem3_reg[52][24]  ( .D(n12876), .SI(\mem3[51][31] ), .SE(test_se), 
        .CLK(n1857), .Q(\mem3[52][24] ), .QN(n29280) );
  SDFFX1 \mem3_reg[51][31]  ( .D(n12875), .SI(\mem3[51][30] ), .SE(test_se), 
        .CLK(n1857), .Q(\mem3[51][31] ), .QN(n29281) );
  SDFFX1 \mem3_reg[51][30]  ( .D(n12874), .SI(\mem3[51][29] ), .SE(test_se), 
        .CLK(n1858), .Q(\mem3[51][30] ), .QN(n29282) );
  SDFFX1 \mem3_reg[51][29]  ( .D(n12873), .SI(\mem3[51][28] ), .SE(test_se), 
        .CLK(n1858), .Q(\mem3[51][29] ), .QN(n29283) );
  SDFFX1 \mem3_reg[51][28]  ( .D(n12872), .SI(\mem3[51][27] ), .SE(test_se), 
        .CLK(n1858), .Q(\mem3[51][28] ), .QN(n29284) );
  SDFFX1 \mem3_reg[51][27]  ( .D(n12871), .SI(\mem3[51][26] ), .SE(test_se), 
        .CLK(n1858), .Q(\mem3[51][27] ), .QN(n29285) );
  SDFFX1 \mem3_reg[51][26]  ( .D(n12870), .SI(\mem3[51][25] ), .SE(test_se), 
        .CLK(n1858), .Q(\mem3[51][26] ), .QN(n29286) );
  SDFFX1 \mem3_reg[51][25]  ( .D(n12869), .SI(\mem3[51][24] ), .SE(test_se), 
        .CLK(n1858), .Q(\mem3[51][25] ), .QN(n29287) );
  SDFFX1 \mem3_reg[51][24]  ( .D(n12868), .SI(\mem3[50][31] ), .SE(test_se), 
        .CLK(n1858), .Q(\mem3[51][24] ), .QN(n29288) );
  SDFFX1 \mem3_reg[50][31]  ( .D(n12867), .SI(\mem3[50][30] ), .SE(test_se), 
        .CLK(n1858), .Q(\mem3[50][31] ), .QN(n29289) );
  SDFFX1 \mem3_reg[50][30]  ( .D(n12866), .SI(\mem3[50][29] ), .SE(test_se), 
        .CLK(n1858), .Q(\mem3[50][30] ), .QN(n29290) );
  SDFFX1 \mem3_reg[50][29]  ( .D(n12865), .SI(\mem3[50][28] ), .SE(test_se), 
        .CLK(n1858), .Q(\mem3[50][29] ), .QN(n29291) );
  SDFFX1 \mem3_reg[50][28]  ( .D(n12864), .SI(\mem3[50][27] ), .SE(test_se), 
        .CLK(n1858), .Q(\mem3[50][28] ), .QN(n29292) );
  SDFFX1 \mem3_reg[50][27]  ( .D(n12863), .SI(\mem3[50][26] ), .SE(test_se), 
        .CLK(n1858), .Q(\mem3[50][27] ), .QN(n29293) );
  SDFFX1 \mem3_reg[50][26]  ( .D(n12862), .SI(\mem3[50][25] ), .SE(test_se), 
        .CLK(n1859), .Q(\mem3[50][26] ), .QN(n29294) );
  SDFFX1 \mem3_reg[50][25]  ( .D(n12861), .SI(\mem3[50][24] ), .SE(test_se), 
        .CLK(n1859), .Q(\mem3[50][25] ), .QN(n29295) );
  SDFFX1 \mem3_reg[50][24]  ( .D(n12860), .SI(\mem3[49][31] ), .SE(test_se), 
        .CLK(n1859), .Q(\mem3[50][24] ), .QN(n29296) );
  SDFFX1 \mem3_reg[49][31]  ( .D(n12859), .SI(\mem3[49][30] ), .SE(test_se), 
        .CLK(n1859), .Q(\mem3[49][31] ), .QN(n29297) );
  SDFFX1 \mem3_reg[49][30]  ( .D(n12858), .SI(\mem3[49][29] ), .SE(test_se), 
        .CLK(n1859), .Q(\mem3[49][30] ), .QN(n29298) );
  SDFFX1 \mem3_reg[49][29]  ( .D(n12857), .SI(\mem3[49][28] ), .SE(test_se), 
        .CLK(n1859), .Q(\mem3[49][29] ), .QN(n29299) );
  SDFFX1 \mem3_reg[49][28]  ( .D(n12856), .SI(\mem3[49][27] ), .SE(test_se), 
        .CLK(n1859), .Q(\mem3[49][28] ), .QN(n29300) );
  SDFFX1 \mem3_reg[49][27]  ( .D(n12855), .SI(\mem3[49][26] ), .SE(test_se), 
        .CLK(n1859), .Q(\mem3[49][27] ), .QN(n29301) );
  SDFFX1 \mem3_reg[49][26]  ( .D(n12854), .SI(\mem3[49][25] ), .SE(test_se), 
        .CLK(n1859), .Q(\mem3[49][26] ), .QN(n29302) );
  SDFFX1 \mem3_reg[49][25]  ( .D(n12853), .SI(\mem3[49][24] ), .SE(test_se), 
        .CLK(n1859), .Q(\mem3[49][25] ), .QN(n29303) );
  SDFFX1 \mem3_reg[49][24]  ( .D(n12852), .SI(\mem3[48][31] ), .SE(test_se), 
        .CLK(n1859), .Q(\mem3[49][24] ), .QN(n29304) );
  SDFFX1 \mem3_reg[48][31]  ( .D(n12851), .SI(\mem3[48][30] ), .SE(test_se), 
        .CLK(n1859), .Q(\mem3[48][31] ), .QN(n29305) );
  SDFFX1 \mem3_reg[48][30]  ( .D(n12850), .SI(\mem3[48][29] ), .SE(test_se), 
        .CLK(n1860), .Q(\mem3[48][30] ), .QN(n29306) );
  SDFFX1 \mem3_reg[48][29]  ( .D(n12849), .SI(\mem3[48][28] ), .SE(test_se), 
        .CLK(n1860), .Q(\mem3[48][29] ), .QN(n29307) );
  SDFFX1 \mem3_reg[48][28]  ( .D(n12848), .SI(\mem3[48][27] ), .SE(test_se), 
        .CLK(n1860), .Q(\mem3[48][28] ), .QN(n29308) );
  SDFFX1 \mem3_reg[48][27]  ( .D(n12847), .SI(\mem3[48][26] ), .SE(test_se), 
        .CLK(n1860), .Q(\mem3[48][27] ), .QN(n29309) );
  SDFFX1 \mem3_reg[48][26]  ( .D(n12846), .SI(\mem3[48][25] ), .SE(test_se), 
        .CLK(n1860), .Q(\mem3[48][26] ), .QN(n29310) );
  SDFFX1 \mem3_reg[48][25]  ( .D(n12845), .SI(\mem3[48][24] ), .SE(test_se), 
        .CLK(n1860), .Q(\mem3[48][25] ), .QN(n29311) );
  SDFFX1 \mem3_reg[48][24]  ( .D(n12844), .SI(\mem3[47][31] ), .SE(test_se), 
        .CLK(n1860), .Q(\mem3[48][24] ), .QN(n29312) );
  SDFFX1 \mem3_reg[47][31]  ( .D(n12843), .SI(\mem3[47][30] ), .SE(test_se), 
        .CLK(n1860), .Q(\mem3[47][31] ), .QN(n29313) );
  SDFFX1 \mem3_reg[47][30]  ( .D(n12842), .SI(\mem3[47][29] ), .SE(test_se), 
        .CLK(n1860), .Q(\mem3[47][30] ), .QN(n29314) );
  SDFFX1 \mem3_reg[47][29]  ( .D(n12841), .SI(\mem3[47][28] ), .SE(test_se), 
        .CLK(n1860), .Q(\mem3[47][29] ), .QN(n29315) );
  SDFFX1 \mem3_reg[47][28]  ( .D(n12840), .SI(\mem3[47][27] ), .SE(test_se), 
        .CLK(n1860), .Q(\mem3[47][28] ), .QN(n29316) );
  SDFFX1 \mem3_reg[47][27]  ( .D(n12839), .SI(\mem3[47][26] ), .SE(test_se), 
        .CLK(n1860), .Q(\mem3[47][27] ), .QN(n29317) );
  SDFFX1 \mem3_reg[47][26]  ( .D(n12838), .SI(\mem3[47][25] ), .SE(test_se), 
        .CLK(n1861), .Q(\mem3[47][26] ), .QN(n29318) );
  SDFFX1 \mem3_reg[47][25]  ( .D(n12837), .SI(\mem3[47][24] ), .SE(test_se), 
        .CLK(n1861), .Q(\mem3[47][25] ), .QN(n29319) );
  SDFFX1 \mem3_reg[47][24]  ( .D(n12836), .SI(\mem3[46][31] ), .SE(test_se), 
        .CLK(n1861), .Q(\mem3[47][24] ), .QN(n29320) );
  SDFFX1 \mem3_reg[46][31]  ( .D(n12835), .SI(\mem3[46][30] ), .SE(test_se), 
        .CLK(n1861), .Q(\mem3[46][31] ), .QN(n29321) );
  SDFFX1 \mem3_reg[46][30]  ( .D(n12834), .SI(\mem3[46][29] ), .SE(test_se), 
        .CLK(n1861), .Q(\mem3[46][30] ), .QN(n29322) );
  SDFFX1 \mem3_reg[46][29]  ( .D(n12833), .SI(\mem3[46][28] ), .SE(test_se), 
        .CLK(n1861), .Q(\mem3[46][29] ), .QN(n29323) );
  SDFFX1 \mem3_reg[46][28]  ( .D(n12832), .SI(\mem3[46][27] ), .SE(test_se), 
        .CLK(n1861), .Q(\mem3[46][28] ), .QN(n29324) );
  SDFFX1 \mem3_reg[46][27]  ( .D(n12831), .SI(\mem3[46][26] ), .SE(test_se), 
        .CLK(n1861), .Q(\mem3[46][27] ), .QN(n29325) );
  SDFFX1 \mem3_reg[46][26]  ( .D(n12830), .SI(\mem3[46][25] ), .SE(test_se), 
        .CLK(n1861), .Q(\mem3[46][26] ), .QN(n29326) );
  SDFFX1 \mem3_reg[46][25]  ( .D(n12829), .SI(\mem3[46][24] ), .SE(test_se), 
        .CLK(n1861), .Q(\mem3[46][25] ), .QN(n29327) );
  SDFFX1 \mem3_reg[46][24]  ( .D(n12828), .SI(\mem3[45][31] ), .SE(test_se), 
        .CLK(n1861), .Q(\mem3[46][24] ), .QN(n29328) );
  SDFFX1 \mem3_reg[45][31]  ( .D(n12827), .SI(\mem3[45][30] ), .SE(test_se), 
        .CLK(n1861), .Q(\mem3[45][31] ), .QN(n29329) );
  SDFFX1 \mem3_reg[45][30]  ( .D(n12826), .SI(\mem3[45][29] ), .SE(test_se), 
        .CLK(n1862), .Q(\mem3[45][30] ), .QN(n29330) );
  SDFFX1 \mem3_reg[45][29]  ( .D(n12825), .SI(\mem3[45][28] ), .SE(test_se), 
        .CLK(n1862), .Q(\mem3[45][29] ), .QN(n29331) );
  SDFFX1 \mem3_reg[45][28]  ( .D(n12824), .SI(\mem3[45][27] ), .SE(test_se), 
        .CLK(n1862), .Q(\mem3[45][28] ), .QN(n29332) );
  SDFFX1 \mem3_reg[45][27]  ( .D(n12823), .SI(\mem3[45][26] ), .SE(test_se), 
        .CLK(n1862), .Q(\mem3[45][27] ), .QN(n29333) );
  SDFFX1 \mem3_reg[45][26]  ( .D(n12822), .SI(\mem3[45][25] ), .SE(test_se), 
        .CLK(n1862), .Q(\mem3[45][26] ), .QN(n29334) );
  SDFFX1 \mem3_reg[45][25]  ( .D(n12821), .SI(\mem3[45][24] ), .SE(test_se), 
        .CLK(n1862), .Q(\mem3[45][25] ), .QN(n29335) );
  SDFFX1 \mem3_reg[45][24]  ( .D(n12820), .SI(\mem3[44][31] ), .SE(test_se), 
        .CLK(n1862), .Q(\mem3[45][24] ), .QN(n29336) );
  SDFFX1 \mem3_reg[44][31]  ( .D(n12819), .SI(\mem3[44][30] ), .SE(test_se), 
        .CLK(n1862), .Q(\mem3[44][31] ), .QN(n29337) );
  SDFFX1 \mem3_reg[44][30]  ( .D(n12818), .SI(\mem3[44][29] ), .SE(test_se), 
        .CLK(n1862), .Q(\mem3[44][30] ), .QN(n29338) );
  SDFFX1 \mem3_reg[44][29]  ( .D(n12817), .SI(\mem3[44][28] ), .SE(test_se), 
        .CLK(n1862), .Q(\mem3[44][29] ), .QN(n29339) );
  SDFFX1 \mem3_reg[44][28]  ( .D(n12816), .SI(\mem3[44][27] ), .SE(test_se), 
        .CLK(n1862), .Q(\mem3[44][28] ), .QN(n29340) );
  SDFFX1 \mem3_reg[44][27]  ( .D(n12815), .SI(\mem3[44][26] ), .SE(test_se), 
        .CLK(n1862), .Q(\mem3[44][27] ), .QN(n29341) );
  SDFFX1 \mem3_reg[44][26]  ( .D(n12814), .SI(\mem3[44][25] ), .SE(test_se), 
        .CLK(n1863), .Q(\mem3[44][26] ), .QN(n29342) );
  SDFFX1 \mem3_reg[44][25]  ( .D(n12813), .SI(\mem3[44][24] ), .SE(test_se), 
        .CLK(n1863), .Q(\mem3[44][25] ), .QN(n29343) );
  SDFFX1 \mem3_reg[44][24]  ( .D(n12812), .SI(\mem3[43][31] ), .SE(test_se), 
        .CLK(n1863), .Q(\mem3[44][24] ), .QN(n29344) );
  SDFFX1 \mem3_reg[43][31]  ( .D(n12811), .SI(\mem3[43][30] ), .SE(test_se), 
        .CLK(n1863), .Q(\mem3[43][31] ), .QN(n29345) );
  SDFFX1 \mem3_reg[43][30]  ( .D(n12810), .SI(\mem3[43][29] ), .SE(test_se), 
        .CLK(n1863), .Q(\mem3[43][30] ), .QN(n29346) );
  SDFFX1 \mem3_reg[43][29]  ( .D(n12809), .SI(\mem3[43][28] ), .SE(test_se), 
        .CLK(n1863), .Q(\mem3[43][29] ), .QN(n29347) );
  SDFFX1 \mem3_reg[43][28]  ( .D(n12808), .SI(\mem3[43][27] ), .SE(test_se), 
        .CLK(n1863), .Q(\mem3[43][28] ), .QN(n29348) );
  SDFFX1 \mem3_reg[43][27]  ( .D(n12807), .SI(\mem3[43][26] ), .SE(test_se), 
        .CLK(n1863), .Q(\mem3[43][27] ), .QN(n29349) );
  SDFFX1 \mem3_reg[43][26]  ( .D(n12806), .SI(\mem3[43][25] ), .SE(test_se), 
        .CLK(n1863), .Q(\mem3[43][26] ), .QN(n29350) );
  SDFFX1 \mem3_reg[43][25]  ( .D(n12805), .SI(\mem3[43][24] ), .SE(test_se), 
        .CLK(n1863), .Q(\mem3[43][25] ), .QN(n29351) );
  SDFFX1 \mem3_reg[43][24]  ( .D(n12804), .SI(\mem3[42][31] ), .SE(test_se), 
        .CLK(n1863), .Q(\mem3[43][24] ), .QN(n29352) );
  SDFFX1 \mem3_reg[42][31]  ( .D(n12803), .SI(\mem3[42][30] ), .SE(test_se), 
        .CLK(n1863), .Q(\mem3[42][31] ), .QN(n29353) );
  SDFFX1 \mem3_reg[42][30]  ( .D(n12802), .SI(\mem3[42][29] ), .SE(test_se), 
        .CLK(n1864), .Q(\mem3[42][30] ), .QN(n29354) );
  SDFFX1 \mem3_reg[42][29]  ( .D(n12801), .SI(\mem3[42][28] ), .SE(test_se), 
        .CLK(n1864), .Q(\mem3[42][29] ), .QN(n29355) );
  SDFFX1 \mem3_reg[42][28]  ( .D(n12800), .SI(\mem3[42][27] ), .SE(test_se), 
        .CLK(n1864), .Q(\mem3[42][28] ), .QN(n29356) );
  SDFFX1 \mem3_reg[42][27]  ( .D(n12799), .SI(\mem3[42][26] ), .SE(test_se), 
        .CLK(n1864), .Q(\mem3[42][27] ), .QN(n29357) );
  SDFFX1 \mem3_reg[42][26]  ( .D(n12798), .SI(\mem3[42][25] ), .SE(test_se), 
        .CLK(n1864), .Q(\mem3[42][26] ), .QN(n29358) );
  SDFFX1 \mem3_reg[42][25]  ( .D(n12797), .SI(\mem3[42][24] ), .SE(test_se), 
        .CLK(n1864), .Q(\mem3[42][25] ), .QN(n29359) );
  SDFFX1 \mem3_reg[42][24]  ( .D(n12796), .SI(\mem3[41][31] ), .SE(test_se), 
        .CLK(n1864), .Q(\mem3[42][24] ), .QN(n29360) );
  SDFFX1 \mem3_reg[41][31]  ( .D(n12795), .SI(\mem3[41][30] ), .SE(test_se), 
        .CLK(n1864), .Q(\mem3[41][31] ), .QN(n29361) );
  SDFFX1 \mem3_reg[41][30]  ( .D(n12794), .SI(\mem3[41][29] ), .SE(test_se), 
        .CLK(n1864), .Q(\mem3[41][30] ), .QN(n29362) );
  SDFFX1 \mem3_reg[41][29]  ( .D(n12793), .SI(\mem3[41][28] ), .SE(test_se), 
        .CLK(n1864), .Q(\mem3[41][29] ), .QN(n29363) );
  SDFFX1 \mem3_reg[41][28]  ( .D(n12792), .SI(\mem3[41][27] ), .SE(test_se), 
        .CLK(n1864), .Q(\mem3[41][28] ), .QN(n29364) );
  SDFFX1 \mem3_reg[41][27]  ( .D(n12791), .SI(\mem3[41][26] ), .SE(test_se), 
        .CLK(n1864), .Q(\mem3[41][27] ), .QN(n29365) );
  SDFFX1 \mem3_reg[41][26]  ( .D(n12790), .SI(\mem3[41][25] ), .SE(test_se), 
        .CLK(n1865), .Q(\mem3[41][26] ), .QN(n29366) );
  SDFFX1 \mem3_reg[41][25]  ( .D(n12789), .SI(\mem3[41][24] ), .SE(test_se), 
        .CLK(n1865), .Q(\mem3[41][25] ), .QN(n29367) );
  SDFFX1 \mem3_reg[41][24]  ( .D(n12788), .SI(\mem3[40][31] ), .SE(test_se), 
        .CLK(n1865), .Q(\mem3[41][24] ), .QN(n29368) );
  SDFFX1 \mem3_reg[40][31]  ( .D(n12787), .SI(\mem3[40][30] ), .SE(test_se), 
        .CLK(n1865), .Q(\mem3[40][31] ), .QN(n29369) );
  SDFFX1 \mem3_reg[40][30]  ( .D(n12786), .SI(\mem3[40][29] ), .SE(test_se), 
        .CLK(n1865), .Q(\mem3[40][30] ), .QN(n29370) );
  SDFFX1 \mem3_reg[40][29]  ( .D(n12785), .SI(\mem3[40][28] ), .SE(test_se), 
        .CLK(n1865), .Q(\mem3[40][29] ), .QN(n29371) );
  SDFFX1 \mem3_reg[40][28]  ( .D(n12784), .SI(\mem3[40][27] ), .SE(test_se), 
        .CLK(n1865), .Q(\mem3[40][28] ), .QN(n29372) );
  SDFFX1 \mem3_reg[40][27]  ( .D(n12783), .SI(\mem3[40][26] ), .SE(test_se), 
        .CLK(n1865), .Q(\mem3[40][27] ), .QN(n29373) );
  SDFFX1 \mem3_reg[40][26]  ( .D(n12782), .SI(\mem3[40][25] ), .SE(test_se), 
        .CLK(n1865), .Q(\mem3[40][26] ), .QN(n29374) );
  SDFFX1 \mem3_reg[40][25]  ( .D(n12781), .SI(\mem3[40][24] ), .SE(test_se), 
        .CLK(n1865), .Q(\mem3[40][25] ), .QN(n29375) );
  SDFFX1 \mem3_reg[40][24]  ( .D(n12780), .SI(\mem3[39][31] ), .SE(test_se), 
        .CLK(n1865), .Q(\mem3[40][24] ), .QN(n29376) );
  SDFFX1 \mem3_reg[39][31]  ( .D(n12779), .SI(\mem3[39][30] ), .SE(test_se), 
        .CLK(n1865), .Q(\mem3[39][31] ), .QN(n29377) );
  SDFFX1 \mem3_reg[39][30]  ( .D(n12778), .SI(\mem3[39][29] ), .SE(test_se), 
        .CLK(n1866), .Q(\mem3[39][30] ), .QN(n29378) );
  SDFFX1 \mem3_reg[39][29]  ( .D(n12777), .SI(\mem3[39][28] ), .SE(test_se), 
        .CLK(n1866), .Q(\mem3[39][29] ), .QN(n29379) );
  SDFFX1 \mem3_reg[39][28]  ( .D(n12776), .SI(\mem3[39][27] ), .SE(test_se), 
        .CLK(n1866), .Q(\mem3[39][28] ), .QN(n29380) );
  SDFFX1 \mem3_reg[39][27]  ( .D(n12775), .SI(\mem3[39][26] ), .SE(test_se), 
        .CLK(n1866), .Q(\mem3[39][27] ), .QN(n29381) );
  SDFFX1 \mem3_reg[39][26]  ( .D(n12774), .SI(\mem3[39][25] ), .SE(test_se), 
        .CLK(n1866), .Q(\mem3[39][26] ), .QN(n29382) );
  SDFFX1 \mem3_reg[39][25]  ( .D(n12773), .SI(\mem3[39][24] ), .SE(test_se), 
        .CLK(n1866), .Q(\mem3[39][25] ), .QN(n29383) );
  SDFFX1 \mem3_reg[39][24]  ( .D(n12772), .SI(\mem3[38][31] ), .SE(test_se), 
        .CLK(n1866), .Q(\mem3[39][24] ), .QN(n29384) );
  SDFFX1 \mem3_reg[38][31]  ( .D(n12771), .SI(\mem3[38][30] ), .SE(test_se), 
        .CLK(n1866), .Q(\mem3[38][31] ), .QN(n29385) );
  SDFFX1 \mem3_reg[38][30]  ( .D(n12770), .SI(\mem3[38][29] ), .SE(test_se), 
        .CLK(n1866), .Q(\mem3[38][30] ), .QN(n29386) );
  SDFFX1 \mem3_reg[38][29]  ( .D(n12769), .SI(\mem3[38][28] ), .SE(test_se), 
        .CLK(n1866), .Q(\mem3[38][29] ), .QN(n29387) );
  SDFFX1 \mem3_reg[38][28]  ( .D(n12768), .SI(\mem3[38][27] ), .SE(test_se), 
        .CLK(n1866), .Q(\mem3[38][28] ), .QN(n29388) );
  SDFFX1 \mem3_reg[38][27]  ( .D(n12767), .SI(\mem3[38][26] ), .SE(test_se), 
        .CLK(n1866), .Q(\mem3[38][27] ), .QN(n29389) );
  SDFFX1 \mem3_reg[38][26]  ( .D(n12766), .SI(\mem3[38][25] ), .SE(test_se), 
        .CLK(n1867), .Q(\mem3[38][26] ), .QN(n29390) );
  SDFFX1 \mem3_reg[38][25]  ( .D(n12765), .SI(\mem3[38][24] ), .SE(test_se), 
        .CLK(n1867), .Q(\mem3[38][25] ), .QN(n29391) );
  SDFFX1 \mem3_reg[38][24]  ( .D(n12764), .SI(\mem3[37][31] ), .SE(test_se), 
        .CLK(n1867), .Q(\mem3[38][24] ), .QN(n29392) );
  SDFFX1 \mem3_reg[37][31]  ( .D(n12763), .SI(\mem3[37][30] ), .SE(test_se), 
        .CLK(n1867), .Q(\mem3[37][31] ), .QN(n29393) );
  SDFFX1 \mem3_reg[37][30]  ( .D(n12762), .SI(\mem3[37][29] ), .SE(test_se), 
        .CLK(n1867), .Q(\mem3[37][30] ), .QN(n29394) );
  SDFFX1 \mem3_reg[37][29]  ( .D(n12761), .SI(\mem3[37][28] ), .SE(test_se), 
        .CLK(n1867), .Q(\mem3[37][29] ), .QN(n29395) );
  SDFFX1 \mem3_reg[37][28]  ( .D(n12760), .SI(\mem3[37][27] ), .SE(test_se), 
        .CLK(n1867), .Q(\mem3[37][28] ), .QN(n29396) );
  SDFFX1 \mem3_reg[37][27]  ( .D(n12759), .SI(\mem3[37][26] ), .SE(test_se), 
        .CLK(n1867), .Q(\mem3[37][27] ), .QN(n29397) );
  SDFFX1 \mem3_reg[37][26]  ( .D(n12758), .SI(\mem3[37][25] ), .SE(test_se), 
        .CLK(n1867), .Q(\mem3[37][26] ), .QN(n29398) );
  SDFFX1 \mem3_reg[37][25]  ( .D(n12757), .SI(\mem3[37][24] ), .SE(test_se), 
        .CLK(n1867), .Q(\mem3[37][25] ), .QN(n29399) );
  SDFFX1 \mem3_reg[37][24]  ( .D(n12756), .SI(\mem3[36][31] ), .SE(test_se), 
        .CLK(n1867), .Q(\mem3[37][24] ), .QN(n29400) );
  SDFFX1 \mem3_reg[36][31]  ( .D(n12755), .SI(\mem3[36][30] ), .SE(test_se), 
        .CLK(n1867), .Q(\mem3[36][31] ), .QN(n29401) );
  SDFFX1 \mem3_reg[36][30]  ( .D(n12754), .SI(\mem3[36][29] ), .SE(test_se), 
        .CLK(n1868), .Q(\mem3[36][30] ), .QN(n29402) );
  SDFFX1 \mem3_reg[36][29]  ( .D(n12753), .SI(\mem3[36][28] ), .SE(test_se), 
        .CLK(n1868), .Q(\mem3[36][29] ), .QN(n29403) );
  SDFFX1 \mem3_reg[36][28]  ( .D(n12752), .SI(\mem3[36][27] ), .SE(test_se), 
        .CLK(n1868), .Q(\mem3[36][28] ), .QN(n29404) );
  SDFFX1 \mem3_reg[36][27]  ( .D(n12751), .SI(\mem3[36][26] ), .SE(test_se), 
        .CLK(n1868), .Q(\mem3[36][27] ), .QN(n29405) );
  SDFFX1 \mem3_reg[36][26]  ( .D(n12750), .SI(\mem3[36][25] ), .SE(test_se), 
        .CLK(n1868), .Q(\mem3[36][26] ), .QN(n29406) );
  SDFFX1 \mem3_reg[36][25]  ( .D(n12749), .SI(\mem3[36][24] ), .SE(test_se), 
        .CLK(n1868), .Q(\mem3[36][25] ), .QN(n29407) );
  SDFFX1 \mem3_reg[36][24]  ( .D(n12748), .SI(\mem3[35][31] ), .SE(test_se), 
        .CLK(n1868), .Q(\mem3[36][24] ), .QN(n29408) );
  SDFFX1 \mem3_reg[35][31]  ( .D(n12747), .SI(\mem3[35][30] ), .SE(test_se), 
        .CLK(n1868), .Q(\mem3[35][31] ), .QN(n29409) );
  SDFFX1 \mem3_reg[35][30]  ( .D(n12746), .SI(\mem3[35][29] ), .SE(test_se), 
        .CLK(n1868), .Q(\mem3[35][30] ), .QN(n29410) );
  SDFFX1 \mem3_reg[35][29]  ( .D(n12745), .SI(\mem3[35][28] ), .SE(test_se), 
        .CLK(n1868), .Q(\mem3[35][29] ), .QN(n29411) );
  SDFFX1 \mem3_reg[35][28]  ( .D(n12744), .SI(\mem3[35][27] ), .SE(test_se), 
        .CLK(n1868), .Q(\mem3[35][28] ), .QN(n29412) );
  SDFFX1 \mem3_reg[35][27]  ( .D(n12743), .SI(\mem3[35][26] ), .SE(test_se), 
        .CLK(n1868), .Q(\mem3[35][27] ), .QN(n29413) );
  SDFFX1 \mem3_reg[35][26]  ( .D(n12742), .SI(\mem3[35][25] ), .SE(test_se), 
        .CLK(n1869), .Q(\mem3[35][26] ), .QN(n29414) );
  SDFFX1 \mem3_reg[35][25]  ( .D(n12741), .SI(\mem3[35][24] ), .SE(test_se), 
        .CLK(n1869), .Q(\mem3[35][25] ), .QN(n29415) );
  SDFFX1 \mem3_reg[35][24]  ( .D(n12740), .SI(\mem3[34][31] ), .SE(test_se), 
        .CLK(n1869), .Q(\mem3[35][24] ), .QN(n29416) );
  SDFFX1 \mem3_reg[34][31]  ( .D(n12739), .SI(\mem3[34][30] ), .SE(test_se), 
        .CLK(n1869), .Q(\mem3[34][31] ), .QN(n29417) );
  SDFFX1 \mem3_reg[34][30]  ( .D(n12738), .SI(\mem3[34][29] ), .SE(test_se), 
        .CLK(n1869), .Q(\mem3[34][30] ), .QN(n29418) );
  SDFFX1 \mem3_reg[34][29]  ( .D(n12737), .SI(\mem3[34][28] ), .SE(test_se), 
        .CLK(n1869), .Q(\mem3[34][29] ), .QN(n29419) );
  SDFFX1 \mem3_reg[34][28]  ( .D(n12736), .SI(\mem3[34][27] ), .SE(test_se), 
        .CLK(n1869), .Q(\mem3[34][28] ), .QN(n29420) );
  SDFFX1 \mem3_reg[34][27]  ( .D(n12735), .SI(\mem3[34][26] ), .SE(test_se), 
        .CLK(n1869), .Q(\mem3[34][27] ), .QN(n29421) );
  SDFFX1 \mem3_reg[34][26]  ( .D(n12734), .SI(\mem3[34][25] ), .SE(test_se), 
        .CLK(n1869), .Q(\mem3[34][26] ), .QN(n29422) );
  SDFFX1 \mem3_reg[34][25]  ( .D(n12733), .SI(\mem3[34][24] ), .SE(test_se), 
        .CLK(n1869), .Q(\mem3[34][25] ), .QN(n29423) );
  SDFFX1 \mem3_reg[34][24]  ( .D(n12732), .SI(\mem3[33][31] ), .SE(test_se), 
        .CLK(n1869), .Q(\mem3[34][24] ), .QN(n29424) );
  SDFFX1 \mem3_reg[33][31]  ( .D(n12731), .SI(\mem3[33][30] ), .SE(test_se), 
        .CLK(n1869), .Q(\mem3[33][31] ), .QN(n29425) );
  SDFFX1 \mem3_reg[33][30]  ( .D(n12730), .SI(\mem3[33][29] ), .SE(test_se), 
        .CLK(n1870), .Q(\mem3[33][30] ), .QN(n29426) );
  SDFFX1 \mem3_reg[33][29]  ( .D(n12729), .SI(\mem3[33][28] ), .SE(test_se), 
        .CLK(n1870), .Q(\mem3[33][29] ), .QN(n29427) );
  SDFFX1 \mem3_reg[33][28]  ( .D(n12728), .SI(\mem3[33][27] ), .SE(test_se), 
        .CLK(n1870), .Q(\mem3[33][28] ), .QN(n29428) );
  SDFFX1 \mem3_reg[33][27]  ( .D(n12727), .SI(\mem3[33][26] ), .SE(test_se), 
        .CLK(n1870), .Q(\mem3[33][27] ), .QN(n29429) );
  SDFFX1 \mem3_reg[33][26]  ( .D(n12726), .SI(\mem3[33][25] ), .SE(test_se), 
        .CLK(n1870), .Q(\mem3[33][26] ), .QN(n29430) );
  SDFFX1 \mem3_reg[33][25]  ( .D(n12725), .SI(\mem3[33][24] ), .SE(test_se), 
        .CLK(n1870), .Q(\mem3[33][25] ), .QN(n29431) );
  SDFFX1 \mem3_reg[33][24]  ( .D(n12724), .SI(\mem3[32][31] ), .SE(test_se), 
        .CLK(n1870), .Q(\mem3[33][24] ), .QN(n29432) );
  SDFFX1 \mem3_reg[32][31]  ( .D(n12723), .SI(\mem3[32][30] ), .SE(test_se), 
        .CLK(n1870), .Q(\mem3[32][31] ), .QN(n29433) );
  SDFFX1 \mem3_reg[32][30]  ( .D(n12722), .SI(\mem3[32][29] ), .SE(test_se), 
        .CLK(n1870), .Q(\mem3[32][30] ), .QN(n29434) );
  SDFFX1 \mem3_reg[32][29]  ( .D(n12721), .SI(\mem3[32][28] ), .SE(test_se), 
        .CLK(n1870), .Q(\mem3[32][29] ), .QN(n29435) );
  SDFFX1 \mem3_reg[32][28]  ( .D(n12720), .SI(\mem3[32][27] ), .SE(test_se), 
        .CLK(n1870), .Q(\mem3[32][28] ), .QN(n29436) );
  SDFFX1 \mem3_reg[32][27]  ( .D(n12719), .SI(\mem3[32][26] ), .SE(test_se), 
        .CLK(n1870), .Q(\mem3[32][27] ), .QN(n29437) );
  SDFFX1 \mem3_reg[32][26]  ( .D(n12718), .SI(\mem3[32][25] ), .SE(test_se), 
        .CLK(n1871), .Q(\mem3[32][26] ), .QN(n29438) );
  SDFFX1 \mem3_reg[32][25]  ( .D(n12717), .SI(\mem3[32][24] ), .SE(test_se), 
        .CLK(n1871), .Q(\mem3[32][25] ), .QN(n29439) );
  SDFFX1 \mem3_reg[32][24]  ( .D(n12716), .SI(\mem3[31][31] ), .SE(test_se), 
        .CLK(n1871), .Q(\mem3[32][24] ), .QN(n29440) );
  SDFFX1 \mem3_reg[31][31]  ( .D(n12715), .SI(\mem3[31][30] ), .SE(test_se), 
        .CLK(n1871), .Q(\mem3[31][31] ), .QN(n29441) );
  SDFFX1 \mem3_reg[31][30]  ( .D(n12714), .SI(\mem3[31][29] ), .SE(test_se), 
        .CLK(n1871), .Q(\mem3[31][30] ), .QN(n29442) );
  SDFFX1 \mem3_reg[31][29]  ( .D(n12713), .SI(\mem3[31][28] ), .SE(test_se), 
        .CLK(n1871), .Q(\mem3[31][29] ), .QN(n29443) );
  SDFFX1 \mem3_reg[31][28]  ( .D(n12712), .SI(\mem3[31][27] ), .SE(test_se), 
        .CLK(n1871), .Q(\mem3[31][28] ), .QN(n29444) );
  SDFFX1 \mem3_reg[31][27]  ( .D(n12711), .SI(\mem3[31][26] ), .SE(test_se), 
        .CLK(n1871), .Q(\mem3[31][27] ), .QN(n29445) );
  SDFFX1 \mem3_reg[31][26]  ( .D(n12710), .SI(\mem3[31][25] ), .SE(test_se), 
        .CLK(n1871), .Q(\mem3[31][26] ), .QN(n29446) );
  SDFFX1 \mem3_reg[31][25]  ( .D(n12709), .SI(\mem3[31][24] ), .SE(test_se), 
        .CLK(n1871), .Q(\mem3[31][25] ), .QN(n29447) );
  SDFFX1 \mem3_reg[31][24]  ( .D(n12708), .SI(\mem3[30][31] ), .SE(test_se), 
        .CLK(n1871), .Q(\mem3[31][24] ), .QN(n29448) );
  SDFFX1 \mem3_reg[30][31]  ( .D(n12707), .SI(\mem3[30][30] ), .SE(test_se), 
        .CLK(n1871), .Q(\mem3[30][31] ), .QN(n29449) );
  SDFFX1 \mem3_reg[30][30]  ( .D(n12706), .SI(\mem3[30][29] ), .SE(test_se), 
        .CLK(n1872), .Q(\mem3[30][30] ), .QN(n29450) );
  SDFFX1 \mem3_reg[30][29]  ( .D(n12705), .SI(\mem3[30][28] ), .SE(test_se), 
        .CLK(n1872), .Q(\mem3[30][29] ), .QN(n29451) );
  SDFFX1 \mem3_reg[30][28]  ( .D(n12704), .SI(\mem3[30][27] ), .SE(test_se), 
        .CLK(n1872), .Q(\mem3[30][28] ), .QN(n29452) );
  SDFFX1 \mem3_reg[30][27]  ( .D(n12703), .SI(\mem3[30][26] ), .SE(test_se), 
        .CLK(n1872), .Q(\mem3[30][27] ), .QN(n29453) );
  SDFFX1 \mem3_reg[30][26]  ( .D(n12702), .SI(\mem3[30][25] ), .SE(test_se), 
        .CLK(n1872), .Q(\mem3[30][26] ), .QN(n29454) );
  SDFFX1 \mem3_reg[30][25]  ( .D(n12701), .SI(\mem3[30][24] ), .SE(test_se), 
        .CLK(n1872), .Q(\mem3[30][25] ), .QN(n29455) );
  SDFFX1 \mem3_reg[30][24]  ( .D(n12700), .SI(\mem3[29][31] ), .SE(test_se), 
        .CLK(n1872), .Q(\mem3[30][24] ), .QN(n29456) );
  SDFFX1 \mem3_reg[29][31]  ( .D(n12699), .SI(\mem3[29][30] ), .SE(test_se), 
        .CLK(n1872), .Q(\mem3[29][31] ), .QN(n29457) );
  SDFFX1 \mem3_reg[29][30]  ( .D(n12698), .SI(\mem3[29][29] ), .SE(test_se), 
        .CLK(n1872), .Q(\mem3[29][30] ), .QN(n29458) );
  SDFFX1 \mem3_reg[29][29]  ( .D(n12697), .SI(\mem3[29][28] ), .SE(test_se), 
        .CLK(n1872), .Q(\mem3[29][29] ), .QN(n29459) );
  SDFFX1 \mem3_reg[29][28]  ( .D(n12696), .SI(\mem3[29][27] ), .SE(test_se), 
        .CLK(n1872), .Q(\mem3[29][28] ), .QN(n29460) );
  SDFFX1 \mem3_reg[29][27]  ( .D(n12695), .SI(\mem3[29][26] ), .SE(test_se), 
        .CLK(n1872), .Q(\mem3[29][27] ), .QN(n29461) );
  SDFFX1 \mem3_reg[29][26]  ( .D(n12694), .SI(\mem3[29][25] ), .SE(test_se), 
        .CLK(n1873), .Q(\mem3[29][26] ), .QN(n29462) );
  SDFFX1 \mem3_reg[29][25]  ( .D(n12693), .SI(\mem3[29][24] ), .SE(test_se), 
        .CLK(n1873), .Q(\mem3[29][25] ), .QN(n29463) );
  SDFFX1 \mem3_reg[29][24]  ( .D(n12692), .SI(\mem3[28][31] ), .SE(test_se), 
        .CLK(n1873), .Q(\mem3[29][24] ), .QN(n29464) );
  SDFFX1 \mem3_reg[28][31]  ( .D(n12691), .SI(\mem3[28][30] ), .SE(test_se), 
        .CLK(n1873), .Q(\mem3[28][31] ), .QN(n29465) );
  SDFFX1 \mem3_reg[28][30]  ( .D(n12690), .SI(\mem3[28][29] ), .SE(test_se), 
        .CLK(n1873), .Q(\mem3[28][30] ), .QN(n29466) );
  SDFFX1 \mem3_reg[28][29]  ( .D(n12689), .SI(\mem3[28][28] ), .SE(test_se), 
        .CLK(n1873), .Q(\mem3[28][29] ), .QN(n29467) );
  SDFFX1 \mem3_reg[28][28]  ( .D(n12688), .SI(\mem3[28][27] ), .SE(test_se), 
        .CLK(n1873), .Q(\mem3[28][28] ), .QN(n29468) );
  SDFFX1 \mem3_reg[28][27]  ( .D(n12687), .SI(\mem3[28][26] ), .SE(test_se), 
        .CLK(n1873), .Q(\mem3[28][27] ), .QN(n29469) );
  SDFFX1 \mem3_reg[28][26]  ( .D(n12686), .SI(\mem3[28][25] ), .SE(test_se), 
        .CLK(n1873), .Q(\mem3[28][26] ), .QN(n29470) );
  SDFFX1 \mem3_reg[28][25]  ( .D(n12685), .SI(\mem3[28][24] ), .SE(test_se), 
        .CLK(n1873), .Q(\mem3[28][25] ), .QN(n29471) );
  SDFFX1 \mem3_reg[28][24]  ( .D(n12684), .SI(\mem3[27][31] ), .SE(test_se), 
        .CLK(n1873), .Q(\mem3[28][24] ), .QN(n29472) );
  SDFFX1 \mem3_reg[27][31]  ( .D(n12683), .SI(\mem3[27][30] ), .SE(test_se), 
        .CLK(n1873), .Q(\mem3[27][31] ), .QN(n29473) );
  SDFFX1 \mem3_reg[27][30]  ( .D(n12682), .SI(\mem3[27][29] ), .SE(test_se), 
        .CLK(n1874), .Q(\mem3[27][30] ), .QN(n29474) );
  SDFFX1 \mem3_reg[27][29]  ( .D(n12681), .SI(\mem3[27][28] ), .SE(test_se), 
        .CLK(n1874), .Q(\mem3[27][29] ), .QN(n29475) );
  SDFFX1 \mem3_reg[27][28]  ( .D(n12680), .SI(\mem3[27][27] ), .SE(test_se), 
        .CLK(n1874), .Q(\mem3[27][28] ), .QN(n29476) );
  SDFFX1 \mem3_reg[27][27]  ( .D(n12679), .SI(\mem3[27][26] ), .SE(test_se), 
        .CLK(n1874), .Q(\mem3[27][27] ), .QN(n29477) );
  SDFFX1 \mem3_reg[27][26]  ( .D(n12678), .SI(\mem3[27][25] ), .SE(test_se), 
        .CLK(n1874), .Q(\mem3[27][26] ), .QN(n29478) );
  SDFFX1 \mem3_reg[27][25]  ( .D(n12677), .SI(\mem3[27][24] ), .SE(test_se), 
        .CLK(n1874), .Q(\mem3[27][25] ), .QN(n29479) );
  SDFFX1 \mem3_reg[27][24]  ( .D(n12676), .SI(\mem3[26][31] ), .SE(test_se), 
        .CLK(n1874), .Q(\mem3[27][24] ), .QN(n29480) );
  SDFFX1 \mem3_reg[26][31]  ( .D(n12675), .SI(\mem3[26][30] ), .SE(test_se), 
        .CLK(n1874), .Q(\mem3[26][31] ), .QN(n29481) );
  SDFFX1 \mem3_reg[26][30]  ( .D(n12674), .SI(\mem3[26][29] ), .SE(test_se), 
        .CLK(n1874), .Q(\mem3[26][30] ), .QN(n29482) );
  SDFFX1 \mem3_reg[26][29]  ( .D(n12673), .SI(\mem3[26][28] ), .SE(test_se), 
        .CLK(n1874), .Q(\mem3[26][29] ), .QN(n29483) );
  SDFFX1 \mem3_reg[26][28]  ( .D(n12672), .SI(\mem3[26][27] ), .SE(test_se), 
        .CLK(n1874), .Q(\mem3[26][28] ), .QN(n29484) );
  SDFFX1 \mem3_reg[26][27]  ( .D(n12671), .SI(\mem3[26][26] ), .SE(test_se), 
        .CLK(n1874), .Q(\mem3[26][27] ), .QN(n29485) );
  SDFFX1 \mem3_reg[26][26]  ( .D(n12670), .SI(\mem3[26][25] ), .SE(test_se), 
        .CLK(n1875), .Q(\mem3[26][26] ), .QN(n29486) );
  SDFFX1 \mem3_reg[26][25]  ( .D(n12669), .SI(\mem3[26][24] ), .SE(test_se), 
        .CLK(n1875), .Q(\mem3[26][25] ), .QN(n29487) );
  SDFFX1 \mem3_reg[26][24]  ( .D(n12668), .SI(\mem3[25][31] ), .SE(test_se), 
        .CLK(n1875), .Q(\mem3[26][24] ), .QN(n29488) );
  SDFFX1 \mem3_reg[25][31]  ( .D(n12667), .SI(\mem3[25][30] ), .SE(test_se), 
        .CLK(n1875), .Q(\mem3[25][31] ), .QN(n29489) );
  SDFFX1 \mem3_reg[25][30]  ( .D(n12666), .SI(\mem3[25][29] ), .SE(test_se), 
        .CLK(n1875), .Q(\mem3[25][30] ), .QN(n29490) );
  SDFFX1 \mem3_reg[25][29]  ( .D(n12665), .SI(\mem3[25][28] ), .SE(test_se), 
        .CLK(n1875), .Q(\mem3[25][29] ), .QN(n29491) );
  SDFFX1 \mem3_reg[25][28]  ( .D(n12664), .SI(\mem3[25][27] ), .SE(test_se), 
        .CLK(n1875), .Q(\mem3[25][28] ), .QN(n29492) );
  SDFFX1 \mem3_reg[25][27]  ( .D(n12663), .SI(\mem3[25][26] ), .SE(test_se), 
        .CLK(n1875), .Q(\mem3[25][27] ), .QN(n29493) );
  SDFFX1 \mem3_reg[25][26]  ( .D(n12662), .SI(\mem3[25][25] ), .SE(test_se), 
        .CLK(n1875), .Q(\mem3[25][26] ), .QN(n29494) );
  SDFFX1 \mem3_reg[25][25]  ( .D(n12661), .SI(\mem3[25][24] ), .SE(test_se), 
        .CLK(n1875), .Q(\mem3[25][25] ), .QN(n29495) );
  SDFFX1 \mem3_reg[25][24]  ( .D(n12660), .SI(\mem3[24][31] ), .SE(test_se), 
        .CLK(n1875), .Q(\mem3[25][24] ), .QN(n29496) );
  SDFFX1 \mem3_reg[24][31]  ( .D(n12659), .SI(\mem3[24][30] ), .SE(test_se), 
        .CLK(n1875), .Q(\mem3[24][31] ), .QN(n29497) );
  SDFFX1 \mem3_reg[24][30]  ( .D(n12658), .SI(\mem3[24][29] ), .SE(test_se), 
        .CLK(n1876), .Q(\mem3[24][30] ), .QN(n29498) );
  SDFFX1 \mem3_reg[24][29]  ( .D(n12657), .SI(\mem3[24][28] ), .SE(test_se), 
        .CLK(n1876), .Q(\mem3[24][29] ), .QN(n29499) );
  SDFFX1 \mem3_reg[24][28]  ( .D(n12656), .SI(\mem3[24][27] ), .SE(test_se), 
        .CLK(n1876), .Q(\mem3[24][28] ), .QN(n29500) );
  SDFFX1 \mem3_reg[24][27]  ( .D(n12655), .SI(\mem3[24][26] ), .SE(test_se), 
        .CLK(n1876), .Q(\mem3[24][27] ), .QN(n29501) );
  SDFFX1 \mem3_reg[24][26]  ( .D(n12654), .SI(\mem3[24][25] ), .SE(test_se), 
        .CLK(n1876), .Q(\mem3[24][26] ), .QN(n29502) );
  SDFFX1 \mem3_reg[24][25]  ( .D(n12653), .SI(\mem3[24][24] ), .SE(test_se), 
        .CLK(n1876), .Q(\mem3[24][25] ), .QN(n29503) );
  SDFFX1 \mem3_reg[24][24]  ( .D(n12652), .SI(\mem3[23][31] ), .SE(test_se), 
        .CLK(n1876), .Q(\mem3[24][24] ), .QN(n29504) );
  SDFFX1 \mem3_reg[23][31]  ( .D(n12651), .SI(\mem3[23][30] ), .SE(test_se), 
        .CLK(n1876), .Q(\mem3[23][31] ), .QN(n29505) );
  SDFFX1 \mem3_reg[23][30]  ( .D(n12650), .SI(\mem3[23][29] ), .SE(test_se), 
        .CLK(n1876), .Q(\mem3[23][30] ), .QN(n29506) );
  SDFFX1 \mem3_reg[23][29]  ( .D(n12649), .SI(\mem3[23][28] ), .SE(test_se), 
        .CLK(n1876), .Q(\mem3[23][29] ), .QN(n29507) );
  SDFFX1 \mem3_reg[23][28]  ( .D(n12648), .SI(\mem3[23][27] ), .SE(test_se), 
        .CLK(n1876), .Q(\mem3[23][28] ), .QN(n29508) );
  SDFFX1 \mem3_reg[23][27]  ( .D(n12647), .SI(\mem3[23][26] ), .SE(test_se), 
        .CLK(n1876), .Q(\mem3[23][27] ), .QN(n29509) );
  SDFFX1 \mem3_reg[23][26]  ( .D(n12646), .SI(\mem3[23][25] ), .SE(test_se), 
        .CLK(n1877), .Q(\mem3[23][26] ), .QN(n29510) );
  SDFFX1 \mem3_reg[23][25]  ( .D(n12645), .SI(\mem3[23][24] ), .SE(test_se), 
        .CLK(n1877), .Q(\mem3[23][25] ), .QN(n29511) );
  SDFFX1 \mem3_reg[23][24]  ( .D(n12644), .SI(\mem3[22][31] ), .SE(test_se), 
        .CLK(n1877), .Q(\mem3[23][24] ), .QN(n29512) );
  SDFFX1 \mem3_reg[22][31]  ( .D(n12643), .SI(\mem3[22][30] ), .SE(test_se), 
        .CLK(n1877), .Q(\mem3[22][31] ), .QN(n29513) );
  SDFFX1 \mem3_reg[22][30]  ( .D(n12642), .SI(\mem3[22][29] ), .SE(test_se), 
        .CLK(n1877), .Q(\mem3[22][30] ), .QN(n29514) );
  SDFFX1 \mem3_reg[22][29]  ( .D(n12641), .SI(\mem3[22][28] ), .SE(test_se), 
        .CLK(n1877), .Q(\mem3[22][29] ), .QN(n29515) );
  SDFFX1 \mem3_reg[22][28]  ( .D(n12640), .SI(\mem3[22][27] ), .SE(test_se), 
        .CLK(n1877), .Q(\mem3[22][28] ), .QN(n29516) );
  SDFFX1 \mem3_reg[22][27]  ( .D(n12639), .SI(\mem3[22][26] ), .SE(test_se), 
        .CLK(n1877), .Q(\mem3[22][27] ), .QN(n29517) );
  SDFFX1 \mem3_reg[22][26]  ( .D(n12638), .SI(\mem3[22][25] ), .SE(test_se), 
        .CLK(n1877), .Q(\mem3[22][26] ), .QN(n29518) );
  SDFFX1 \mem3_reg[22][25]  ( .D(n12637), .SI(\mem3[22][24] ), .SE(test_se), 
        .CLK(n1877), .Q(\mem3[22][25] ), .QN(n29519) );
  SDFFX1 \mem3_reg[22][24]  ( .D(n12636), .SI(\mem3[21][31] ), .SE(test_se), 
        .CLK(n1877), .Q(\mem3[22][24] ), .QN(n29520) );
  SDFFX1 \mem3_reg[21][31]  ( .D(n12635), .SI(\mem3[21][30] ), .SE(test_se), 
        .CLK(n1877), .Q(\mem3[21][31] ), .QN(n29521) );
  SDFFX1 \mem3_reg[21][30]  ( .D(n12634), .SI(\mem3[21][29] ), .SE(test_se), 
        .CLK(n1878), .Q(\mem3[21][30] ), .QN(n29522) );
  SDFFX1 \mem3_reg[21][29]  ( .D(n12633), .SI(\mem3[21][28] ), .SE(test_se), 
        .CLK(n1878), .Q(\mem3[21][29] ), .QN(n29523) );
  SDFFX1 \mem3_reg[21][28]  ( .D(n12632), .SI(\mem3[21][27] ), .SE(test_se), 
        .CLK(n1878), .Q(\mem3[21][28] ), .QN(n29524) );
  SDFFX1 \mem3_reg[21][27]  ( .D(n12631), .SI(\mem3[21][26] ), .SE(test_se), 
        .CLK(n1878), .Q(\mem3[21][27] ), .QN(n29525) );
  SDFFX1 \mem3_reg[21][26]  ( .D(n12630), .SI(\mem3[21][25] ), .SE(test_se), 
        .CLK(n1878), .Q(\mem3[21][26] ), .QN(n29526) );
  SDFFX1 \mem3_reg[21][25]  ( .D(n12629), .SI(\mem3[21][24] ), .SE(test_se), 
        .CLK(n1878), .Q(\mem3[21][25] ), .QN(n29527) );
  SDFFX1 \mem3_reg[21][24]  ( .D(n12628), .SI(\mem3[20][31] ), .SE(test_se), 
        .CLK(n1878), .Q(\mem3[21][24] ), .QN(n29528) );
  SDFFX1 \mem3_reg[20][31]  ( .D(n12627), .SI(\mem3[20][30] ), .SE(test_se), 
        .CLK(n1878), .Q(\mem3[20][31] ), .QN(n29529) );
  SDFFX1 \mem3_reg[20][30]  ( .D(n12626), .SI(\mem3[20][29] ), .SE(test_se), 
        .CLK(n1878), .Q(\mem3[20][30] ), .QN(n29530) );
  SDFFX1 \mem3_reg[20][29]  ( .D(n12625), .SI(\mem3[20][28] ), .SE(test_se), 
        .CLK(n1878), .Q(\mem3[20][29] ), .QN(n29531) );
  SDFFX1 \mem3_reg[20][28]  ( .D(n12624), .SI(\mem3[20][27] ), .SE(test_se), 
        .CLK(n1878), .Q(\mem3[20][28] ), .QN(n29532) );
  SDFFX1 \mem3_reg[20][27]  ( .D(n12623), .SI(\mem3[20][26] ), .SE(test_se), 
        .CLK(n1878), .Q(\mem3[20][27] ), .QN(n29533) );
  SDFFX1 \mem3_reg[20][26]  ( .D(n12622), .SI(\mem3[20][25] ), .SE(test_se), 
        .CLK(n1879), .Q(\mem3[20][26] ), .QN(n29534) );
  SDFFX1 \mem3_reg[20][25]  ( .D(n12621), .SI(\mem3[20][24] ), .SE(test_se), 
        .CLK(n1879), .Q(\mem3[20][25] ), .QN(n29535) );
  SDFFX1 \mem3_reg[20][24]  ( .D(n12620), .SI(\mem3[19][31] ), .SE(test_se), 
        .CLK(n1879), .Q(\mem3[20][24] ), .QN(n29536) );
  SDFFX1 \mem3_reg[19][31]  ( .D(n12619), .SI(\mem3[19][30] ), .SE(test_se), 
        .CLK(n1879), .Q(\mem3[19][31] ), .QN(n29537) );
  SDFFX1 \mem3_reg[19][30]  ( .D(n12618), .SI(\mem3[19][29] ), .SE(test_se), 
        .CLK(n1879), .Q(\mem3[19][30] ), .QN(n29538) );
  SDFFX1 \mem3_reg[19][29]  ( .D(n12617), .SI(\mem3[19][28] ), .SE(test_se), 
        .CLK(n1879), .Q(\mem3[19][29] ), .QN(n29539) );
  SDFFX1 \mem3_reg[19][28]  ( .D(n12616), .SI(\mem3[19][27] ), .SE(test_se), 
        .CLK(n1879), .Q(\mem3[19][28] ), .QN(n29540) );
  SDFFX1 \mem3_reg[19][27]  ( .D(n12615), .SI(\mem3[19][26] ), .SE(test_se), 
        .CLK(n1879), .Q(\mem3[19][27] ), .QN(n29541) );
  SDFFX1 \mem3_reg[19][26]  ( .D(n12614), .SI(\mem3[19][25] ), .SE(test_se), 
        .CLK(n1879), .Q(\mem3[19][26] ), .QN(n29542) );
  SDFFX1 \mem3_reg[19][25]  ( .D(n12613), .SI(\mem3[19][24] ), .SE(test_se), 
        .CLK(n1879), .Q(\mem3[19][25] ), .QN(n29543) );
  SDFFX1 \mem3_reg[19][24]  ( .D(n12612), .SI(\mem3[18][31] ), .SE(test_se), 
        .CLK(n1879), .Q(\mem3[19][24] ), .QN(n29544) );
  SDFFX1 \mem3_reg[18][31]  ( .D(n12611), .SI(\mem3[18][30] ), .SE(test_se), 
        .CLK(n1879), .Q(\mem3[18][31] ), .QN(n29545) );
  SDFFX1 \mem3_reg[18][30]  ( .D(n12610), .SI(\mem3[18][29] ), .SE(test_se), 
        .CLK(n1880), .Q(\mem3[18][30] ), .QN(n29546) );
  SDFFX1 \mem3_reg[18][29]  ( .D(n12609), .SI(\mem3[18][28] ), .SE(test_se), 
        .CLK(n1880), .Q(\mem3[18][29] ), .QN(n29547) );
  SDFFX1 \mem3_reg[18][28]  ( .D(n12608), .SI(\mem3[18][27] ), .SE(test_se), 
        .CLK(n1880), .Q(\mem3[18][28] ), .QN(n29548) );
  SDFFX1 \mem3_reg[18][27]  ( .D(n12607), .SI(\mem3[18][26] ), .SE(test_se), 
        .CLK(n1880), .Q(\mem3[18][27] ), .QN(n29549) );
  SDFFX1 \mem3_reg[18][26]  ( .D(n12606), .SI(\mem3[18][25] ), .SE(test_se), 
        .CLK(n1880), .Q(\mem3[18][26] ), .QN(n29550) );
  SDFFX1 \mem3_reg[18][25]  ( .D(n12605), .SI(\mem3[18][24] ), .SE(test_se), 
        .CLK(n1880), .Q(\mem3[18][25] ), .QN(n29551) );
  SDFFX1 \mem3_reg[18][24]  ( .D(n12604), .SI(\mem3[17][31] ), .SE(test_se), 
        .CLK(n1880), .Q(\mem3[18][24] ), .QN(n29552) );
  SDFFX1 \mem3_reg[17][31]  ( .D(n12603), .SI(\mem3[17][30] ), .SE(test_se), 
        .CLK(n1880), .Q(\mem3[17][31] ), .QN(n29553) );
  SDFFX1 \mem3_reg[17][30]  ( .D(n12602), .SI(\mem3[17][29] ), .SE(test_se), 
        .CLK(n1880), .Q(\mem3[17][30] ), .QN(n29554) );
  SDFFX1 \mem3_reg[17][29]  ( .D(n12601), .SI(\mem3[17][28] ), .SE(test_se), 
        .CLK(n1880), .Q(\mem3[17][29] ), .QN(n29555) );
  SDFFX1 \mem3_reg[17][28]  ( .D(n12600), .SI(\mem3[17][27] ), .SE(test_se), 
        .CLK(n1880), .Q(\mem3[17][28] ), .QN(n29556) );
  SDFFX1 \mem3_reg[17][27]  ( .D(n12599), .SI(\mem3[17][26] ), .SE(test_se), 
        .CLK(n1880), .Q(\mem3[17][27] ), .QN(n29557) );
  SDFFX1 \mem3_reg[17][26]  ( .D(n12598), .SI(\mem3[17][25] ), .SE(test_se), 
        .CLK(n1881), .Q(\mem3[17][26] ), .QN(n29558) );
  SDFFX1 \mem3_reg[17][25]  ( .D(n12597), .SI(\mem3[17][24] ), .SE(test_se), 
        .CLK(n1881), .Q(\mem3[17][25] ), .QN(n29559) );
  SDFFX1 \mem3_reg[17][24]  ( .D(n12596), .SI(\mem3[16][31] ), .SE(test_se), 
        .CLK(n1881), .Q(\mem3[17][24] ), .QN(n29560) );
  SDFFX1 \mem3_reg[16][31]  ( .D(n12595), .SI(\mem3[16][30] ), .SE(test_se), 
        .CLK(n1881), .Q(\mem3[16][31] ), .QN(n29561) );
  SDFFX1 \mem3_reg[16][30]  ( .D(n12594), .SI(\mem3[16][29] ), .SE(test_se), 
        .CLK(n1881), .Q(\mem3[16][30] ), .QN(n29562) );
  SDFFX1 \mem3_reg[16][29]  ( .D(n12593), .SI(\mem3[16][28] ), .SE(test_se), 
        .CLK(n1881), .Q(\mem3[16][29] ), .QN(n29563) );
  SDFFX1 \mem3_reg[16][28]  ( .D(n12592), .SI(\mem3[16][27] ), .SE(test_se), 
        .CLK(n1881), .Q(\mem3[16][28] ), .QN(n29564) );
  SDFFX1 \mem3_reg[16][27]  ( .D(n12591), .SI(\mem3[16][26] ), .SE(test_se), 
        .CLK(n1881), .Q(\mem3[16][27] ), .QN(n29565) );
  SDFFX1 \mem3_reg[16][26]  ( .D(n12590), .SI(\mem3[16][25] ), .SE(test_se), 
        .CLK(n1881), .Q(\mem3[16][26] ), .QN(n29566) );
  SDFFX1 \mem3_reg[16][25]  ( .D(n12589), .SI(\mem3[16][24] ), .SE(test_se), 
        .CLK(n1881), .Q(\mem3[16][25] ), .QN(n29567) );
  SDFFX1 \mem3_reg[16][24]  ( .D(n12588), .SI(\mem3[15][31] ), .SE(test_se), 
        .CLK(n1881), .Q(\mem3[16][24] ), .QN(n29568) );
  SDFFX1 \mem3_reg[15][31]  ( .D(n12587), .SI(\mem3[15][30] ), .SE(test_se), 
        .CLK(n1881), .Q(\mem3[15][31] ), .QN(n29569) );
  SDFFX1 \mem3_reg[15][30]  ( .D(n12586), .SI(\mem3[15][29] ), .SE(test_se), 
        .CLK(n1882), .Q(\mem3[15][30] ), .QN(n29570) );
  SDFFX1 \mem3_reg[15][29]  ( .D(n12585), .SI(\mem3[15][28] ), .SE(test_se), 
        .CLK(n1882), .Q(\mem3[15][29] ), .QN(n29571) );
  SDFFX1 \mem3_reg[15][28]  ( .D(n12584), .SI(\mem3[15][27] ), .SE(test_se), 
        .CLK(n1882), .Q(\mem3[15][28] ), .QN(n29572) );
  SDFFX1 \mem3_reg[15][27]  ( .D(n12583), .SI(\mem3[15][26] ), .SE(test_se), 
        .CLK(n1882), .Q(\mem3[15][27] ), .QN(n29573) );
  SDFFX1 \mem3_reg[15][26]  ( .D(n12582), .SI(\mem3[15][25] ), .SE(test_se), 
        .CLK(n1882), .Q(\mem3[15][26] ), .QN(n29574) );
  SDFFX1 \mem3_reg[15][25]  ( .D(n12581), .SI(\mem3[15][24] ), .SE(test_se), 
        .CLK(n1882), .Q(\mem3[15][25] ), .QN(n29575) );
  SDFFX1 \mem3_reg[15][24]  ( .D(n12580), .SI(\mem3[14][31] ), .SE(test_se), 
        .CLK(n1882), .Q(\mem3[15][24] ), .QN(n29576) );
  SDFFX1 \mem3_reg[14][31]  ( .D(n12579), .SI(\mem3[14][30] ), .SE(test_se), 
        .CLK(n1882), .Q(\mem3[14][31] ), .QN(n29577) );
  SDFFX1 \mem3_reg[14][30]  ( .D(n12578), .SI(\mem3[14][29] ), .SE(test_se), 
        .CLK(n1882), .Q(\mem3[14][30] ), .QN(n29578) );
  SDFFX1 \mem3_reg[14][29]  ( .D(n12577), .SI(\mem3[14][28] ), .SE(test_se), 
        .CLK(n1882), .Q(\mem3[14][29] ), .QN(n29579) );
  SDFFX1 \mem3_reg[14][28]  ( .D(n12576), .SI(\mem3[14][27] ), .SE(test_se), 
        .CLK(n1882), .Q(\mem3[14][28] ), .QN(n29580) );
  SDFFX1 \mem3_reg[14][27]  ( .D(n12575), .SI(\mem3[14][26] ), .SE(test_se), 
        .CLK(n1882), .Q(\mem3[14][27] ), .QN(n29581) );
  SDFFX1 \mem3_reg[14][26]  ( .D(n12574), .SI(\mem3[14][25] ), .SE(test_se), 
        .CLK(n1883), .Q(\mem3[14][26] ), .QN(n29582) );
  SDFFX1 \mem3_reg[14][25]  ( .D(n12573), .SI(\mem3[14][24] ), .SE(test_se), 
        .CLK(n1883), .Q(\mem3[14][25] ), .QN(n29583) );
  SDFFX1 \mem3_reg[14][24]  ( .D(n12572), .SI(\mem3[13][31] ), .SE(test_se), 
        .CLK(n1883), .Q(\mem3[14][24] ), .QN(n29584) );
  SDFFX1 \mem3_reg[13][31]  ( .D(n12571), .SI(\mem3[13][30] ), .SE(test_se), 
        .CLK(n1883), .Q(\mem3[13][31] ), .QN(n29585) );
  SDFFX1 \mem3_reg[13][30]  ( .D(n12570), .SI(\mem3[13][29] ), .SE(test_se), 
        .CLK(n1883), .Q(\mem3[13][30] ), .QN(n29586) );
  SDFFX1 \mem3_reg[13][29]  ( .D(n12569), .SI(\mem3[13][28] ), .SE(test_se), 
        .CLK(n1883), .Q(\mem3[13][29] ), .QN(n29587) );
  SDFFX1 \mem3_reg[13][28]  ( .D(n12568), .SI(\mem3[13][27] ), .SE(test_se), 
        .CLK(n1883), .Q(\mem3[13][28] ), .QN(n29588) );
  SDFFX1 \mem3_reg[13][27]  ( .D(n12567), .SI(\mem3[13][26] ), .SE(test_se), 
        .CLK(n1883), .Q(\mem3[13][27] ), .QN(n29589) );
  SDFFX1 \mem3_reg[13][26]  ( .D(n12566), .SI(\mem3[13][25] ), .SE(test_se), 
        .CLK(n1883), .Q(\mem3[13][26] ), .QN(n29590) );
  SDFFX1 \mem3_reg[13][25]  ( .D(n12565), .SI(\mem3[13][24] ), .SE(test_se), 
        .CLK(n1883), .Q(\mem3[13][25] ), .QN(n29591) );
  SDFFX1 \mem3_reg[13][24]  ( .D(n12564), .SI(\mem3[12][31] ), .SE(test_se), 
        .CLK(n1883), .Q(\mem3[13][24] ), .QN(n29592) );
  SDFFX1 \mem3_reg[12][31]  ( .D(n12563), .SI(\mem3[12][30] ), .SE(test_se), 
        .CLK(n1883), .Q(\mem3[12][31] ), .QN(n29593) );
  SDFFX1 \mem3_reg[12][30]  ( .D(n12562), .SI(\mem3[12][29] ), .SE(test_se), 
        .CLK(n1884), .Q(\mem3[12][30] ), .QN(n29594) );
  SDFFX1 \mem3_reg[12][29]  ( .D(n12561), .SI(\mem3[12][28] ), .SE(test_se), 
        .CLK(n1884), .Q(\mem3[12][29] ), .QN(n29595) );
  SDFFX1 \mem3_reg[12][28]  ( .D(n12560), .SI(\mem3[12][27] ), .SE(test_se), 
        .CLK(n1884), .Q(\mem3[12][28] ), .QN(n29596) );
  SDFFX1 \mem3_reg[12][27]  ( .D(n12559), .SI(\mem3[12][26] ), .SE(test_se), 
        .CLK(n1884), .Q(\mem3[12][27] ), .QN(n29597) );
  SDFFX1 \mem3_reg[12][26]  ( .D(n12558), .SI(\mem3[12][25] ), .SE(test_se), 
        .CLK(n1884), .Q(\mem3[12][26] ), .QN(n29598) );
  SDFFX1 \mem3_reg[12][25]  ( .D(n12557), .SI(\mem3[12][24] ), .SE(test_se), 
        .CLK(n1884), .Q(\mem3[12][25] ), .QN(n29599) );
  SDFFX1 \mem3_reg[12][24]  ( .D(n12556), .SI(\mem3[11][31] ), .SE(test_se), 
        .CLK(n1884), .Q(\mem3[12][24] ), .QN(n29600) );
  SDFFX1 \mem3_reg[11][31]  ( .D(n12555), .SI(\mem3[11][30] ), .SE(test_se), 
        .CLK(n2050), .Q(\mem3[11][31] ), .QN(n29601) );
  SDFFX1 \mem3_reg[11][30]  ( .D(n12554), .SI(\mem3[11][29] ), .SE(test_se), 
        .CLK(n2050), .Q(\mem3[11][30] ), .QN(n29602) );
  SDFFX1 \mem3_reg[11][29]  ( .D(n12553), .SI(\mem3[11][28] ), .SE(test_se), 
        .CLK(n2050), .Q(\mem3[11][29] ), .QN(n29603) );
  SDFFX1 \mem3_reg[11][28]  ( .D(n12552), .SI(\mem3[11][27] ), .SE(test_se), 
        .CLK(n2050), .Q(\mem3[11][28] ), .QN(n29604) );
  SDFFX1 \mem3_reg[11][27]  ( .D(n12551), .SI(\mem3[11][26] ), .SE(test_se), 
        .CLK(n2050), .Q(\mem3[11][27] ), .QN(n29605) );
  SDFFX1 \mem3_reg[11][26]  ( .D(n12550), .SI(\mem3[11][25] ), .SE(test_se), 
        .CLK(n2050), .Q(\mem3[11][26] ), .QN(n29606) );
  SDFFX1 \mem3_reg[11][25]  ( .D(n12549), .SI(\mem3[11][24] ), .SE(test_se), 
        .CLK(n2051), .Q(\mem3[11][25] ), .QN(n29607) );
  SDFFX1 \mem3_reg[11][24]  ( .D(n12548), .SI(\mem3[10][31] ), .SE(test_se), 
        .CLK(n2051), .Q(\mem3[11][24] ), .QN(n29608) );
  SDFFX1 \mem3_reg[10][31]  ( .D(n12547), .SI(\mem3[10][30] ), .SE(test_se), 
        .CLK(n2051), .Q(\mem3[10][31] ), .QN(n29609) );
  SDFFX1 \mem3_reg[10][30]  ( .D(n12546), .SI(\mem3[10][29] ), .SE(test_se), 
        .CLK(n2051), .Q(\mem3[10][30] ), .QN(n29610) );
  SDFFX1 \mem3_reg[10][29]  ( .D(n12545), .SI(\mem3[10][28] ), .SE(test_se), 
        .CLK(n2051), .Q(\mem3[10][29] ), .QN(n29611) );
  SDFFX1 \mem3_reg[10][28]  ( .D(n12544), .SI(\mem3[10][27] ), .SE(test_se), 
        .CLK(n2051), .Q(\mem3[10][28] ), .QN(n29612) );
  SDFFX1 \mem3_reg[10][27]  ( .D(n12543), .SI(\mem3[10][26] ), .SE(test_se), 
        .CLK(n2051), .Q(\mem3[10][27] ), .QN(n29613) );
  SDFFX1 \mem3_reg[10][26]  ( .D(n12542), .SI(\mem3[10][25] ), .SE(test_se), 
        .CLK(n2051), .Q(\mem3[10][26] ), .QN(n29614) );
  SDFFX1 \mem3_reg[10][25]  ( .D(n12541), .SI(\mem3[10][24] ), .SE(test_se), 
        .CLK(n2051), .Q(\mem3[10][25] ), .QN(n29615) );
  SDFFX1 \mem3_reg[10][24]  ( .D(n12540), .SI(\mem3[9][31] ), .SE(test_se), 
        .CLK(n2051), .Q(\mem3[10][24] ), .QN(n29616) );
  SDFFX1 \mem3_reg[9][31]  ( .D(n12539), .SI(\mem3[9][30] ), .SE(test_se), 
        .CLK(n2051), .Q(\mem3[9][31] ), .QN(n29617) );
  SDFFX1 \mem3_reg[9][30]  ( .D(n12538), .SI(\mem3[9][29] ), .SE(test_se), 
        .CLK(n2051), .Q(\mem3[9][30] ), .QN(n29618) );
  SDFFX1 \mem3_reg[9][29]  ( .D(n12537), .SI(\mem3[9][28] ), .SE(test_se), 
        .CLK(n2052), .Q(\mem3[9][29] ), .QN(n29619) );
  SDFFX1 \mem3_reg[9][28]  ( .D(n12536), .SI(\mem3[9][27] ), .SE(test_se), 
        .CLK(n2052), .Q(\mem3[9][28] ), .QN(n29620) );
  SDFFX1 \mem3_reg[9][27]  ( .D(n12535), .SI(\mem3[9][26] ), .SE(test_se), 
        .CLK(n2052), .Q(\mem3[9][27] ), .QN(n29621) );
  SDFFX1 \mem3_reg[9][26]  ( .D(n12534), .SI(\mem3[9][25] ), .SE(test_se), 
        .CLK(n2052), .Q(\mem3[9][26] ), .QN(n29622) );
  SDFFX1 \mem3_reg[9][25]  ( .D(n12533), .SI(\mem3[9][24] ), .SE(test_se), 
        .CLK(n2052), .Q(\mem3[9][25] ), .QN(n29623) );
  SDFFX1 \mem3_reg[9][24]  ( .D(n12532), .SI(\mem3[8][31] ), .SE(test_se), 
        .CLK(n2052), .Q(\mem3[9][24] ), .QN(n29624) );
  SDFFX1 \mem3_reg[8][31]  ( .D(n12531), .SI(\mem3[8][30] ), .SE(test_se), 
        .CLK(n2052), .Q(\mem3[8][31] ), .QN(n29625) );
  SDFFX1 \mem3_reg[8][30]  ( .D(n12530), .SI(\mem3[8][29] ), .SE(test_se), 
        .CLK(n2052), .Q(\mem3[8][30] ), .QN(n29626) );
  SDFFX1 \mem3_reg[8][29]  ( .D(n12529), .SI(\mem3[8][28] ), .SE(test_se), 
        .CLK(n2052), .Q(\mem3[8][29] ), .QN(n29627) );
  SDFFX1 \mem3_reg[8][28]  ( .D(n12528), .SI(\mem3[8][27] ), .SE(test_se), 
        .CLK(n2052), .Q(\mem3[8][28] ), .QN(n29628) );
  SDFFX1 \mem3_reg[8][27]  ( .D(n12527), .SI(\mem3[8][26] ), .SE(test_se), 
        .CLK(n2052), .Q(\mem3[8][27] ), .QN(n29629) );
  SDFFX1 \mem3_reg[8][26]  ( .D(n12526), .SI(\mem3[8][25] ), .SE(test_se), 
        .CLK(n2052), .Q(\mem3[8][26] ), .QN(n29630) );
  SDFFX1 \mem3_reg[8][25]  ( .D(n12525), .SI(\mem3[8][24] ), .SE(test_se), 
        .CLK(n2053), .Q(\mem3[8][25] ), .QN(n29631) );
  SDFFX1 \mem3_reg[8][24]  ( .D(n12524), .SI(\mem3[7][31] ), .SE(test_se), 
        .CLK(n2053), .Q(\mem3[8][24] ), .QN(n29632) );
  SDFFX1 \mem3_reg[7][31]  ( .D(n12523), .SI(\mem3[7][30] ), .SE(test_se), 
        .CLK(n2061), .Q(\mem3[7][31] ), .QN(n29633) );
  SDFFX1 \mem3_reg[7][30]  ( .D(n12522), .SI(\mem3[7][29] ), .SE(test_se), 
        .CLK(n2061), .Q(\mem3[7][30] ), .QN(n29634) );
  SDFFX1 \mem3_reg[7][29]  ( .D(n12521), .SI(\mem3[7][28] ), .SE(test_se), 
        .CLK(n2061), .Q(\mem3[7][29] ), .QN(n29635) );
  SDFFX1 \mem3_reg[7][28]  ( .D(n12520), .SI(\mem3[7][27] ), .SE(test_se), 
        .CLK(n2061), .Q(\mem3[7][28] ), .QN(n29636) );
  SDFFX1 \mem3_reg[7][27]  ( .D(n12519), .SI(\mem3[7][26] ), .SE(test_se), 
        .CLK(n2061), .Q(\mem3[7][27] ), .QN(n29637) );
  SDFFX1 \mem3_reg[7][26]  ( .D(n12518), .SI(\mem3[7][25] ), .SE(test_se), 
        .CLK(n2061), .Q(\mem3[7][26] ), .QN(n29638) );
  SDFFX1 \mem3_reg[7][25]  ( .D(n12517), .SI(\mem3[7][24] ), .SE(test_se), 
        .CLK(n2061), .Q(\mem3[7][25] ), .QN(n29639) );
  SDFFX1 \mem3_reg[7][24]  ( .D(n12516), .SI(\mem3[6][31] ), .SE(test_se), 
        .CLK(n2061), .Q(\mem3[7][24] ), .QN(n29640) );
  SDFFX1 \mem3_reg[6][31]  ( .D(n12515), .SI(\mem3[6][30] ), .SE(test_se), 
        .CLK(n2061), .Q(\mem3[6][31] ), .QN(n29641) );
  SDFFX1 \mem3_reg[6][30]  ( .D(n12514), .SI(\mem3[6][29] ), .SE(test_se), 
        .CLK(n2061), .Q(\mem3[6][30] ), .QN(n29642) );
  SDFFX1 \mem3_reg[6][29]  ( .D(n12513), .SI(\mem3[6][28] ), .SE(test_se), 
        .CLK(n2062), .Q(\mem3[6][29] ), .QN(n29643) );
  SDFFX1 \mem3_reg[6][28]  ( .D(n12512), .SI(\mem3[6][27] ), .SE(test_se), 
        .CLK(n2062), .Q(\mem3[6][28] ), .QN(n29644) );
  SDFFX1 \mem3_reg[6][27]  ( .D(n12511), .SI(\mem3[6][26] ), .SE(test_se), 
        .CLK(n2062), .Q(\mem3[6][27] ), .QN(n29645) );
  SDFFX1 \mem3_reg[6][26]  ( .D(n12510), .SI(\mem3[6][25] ), .SE(test_se), 
        .CLK(n2062), .Q(\mem3[6][26] ), .QN(n29646) );
  SDFFX1 \mem3_reg[6][25]  ( .D(n12509), .SI(\mem3[6][24] ), .SE(test_se), 
        .CLK(n2062), .Q(\mem3[6][25] ), .QN(n29647) );
  SDFFX1 \mem3_reg[6][24]  ( .D(n12508), .SI(\mem3[5][31] ), .SE(test_se), 
        .CLK(n2062), .Q(\mem3[6][24] ), .QN(n29648) );
  SDFFX1 \mem3_reg[5][31]  ( .D(n12507), .SI(\mem3[5][30] ), .SE(test_se), 
        .CLK(n2062), .Q(\mem3[5][31] ), .QN(n29649) );
  SDFFX1 \mem3_reg[5][30]  ( .D(n12506), .SI(\mem3[5][29] ), .SE(test_se), 
        .CLK(n2062), .Q(\mem3[5][30] ), .QN(n29650) );
  SDFFX1 \mem3_reg[5][29]  ( .D(n12505), .SI(\mem3[5][28] ), .SE(test_se), 
        .CLK(n2062), .Q(\mem3[5][29] ), .QN(n29651) );
  SDFFX1 \mem3_reg[5][28]  ( .D(n12504), .SI(\mem3[5][27] ), .SE(test_se), 
        .CLK(n2062), .Q(\mem3[5][28] ), .QN(n29652) );
  SDFFX1 \mem3_reg[5][27]  ( .D(n12503), .SI(\mem3[5][26] ), .SE(test_se), 
        .CLK(n2062), .Q(\mem3[5][27] ), .QN(n29653) );
  SDFFX1 \mem3_reg[5][26]  ( .D(n12502), .SI(\mem3[5][25] ), .SE(test_se), 
        .CLK(n2062), .Q(\mem3[5][26] ), .QN(n29654) );
  SDFFX1 \mem3_reg[5][25]  ( .D(n12501), .SI(\mem3[5][24] ), .SE(test_se), 
        .CLK(n2063), .Q(\mem3[5][25] ), .QN(n29655) );
  SDFFX1 \mem3_reg[5][24]  ( .D(n12500), .SI(\mem3[4][31] ), .SE(test_se), 
        .CLK(n2063), .Q(\mem3[5][24] ), .QN(n29656) );
  SDFFX1 \mem3_reg[4][31]  ( .D(n12499), .SI(\mem3[4][30] ), .SE(test_se), 
        .CLK(n2063), .Q(\mem3[4][31] ), .QN(n29657) );
  SDFFX1 \mem3_reg[4][30]  ( .D(n12498), .SI(\mem3[4][29] ), .SE(test_se), 
        .CLK(n2063), .Q(\mem3[4][30] ), .QN(n29658) );
  SDFFX1 \mem3_reg[4][29]  ( .D(n12497), .SI(\mem3[4][28] ), .SE(test_se), 
        .CLK(n2063), .Q(\mem3[4][29] ), .QN(n29659) );
  SDFFX1 \mem3_reg[4][28]  ( .D(n12496), .SI(\mem3[4][27] ), .SE(test_se), 
        .CLK(n2063), .Q(\mem3[4][28] ), .QN(n29660) );
  SDFFX1 \mem3_reg[4][27]  ( .D(n12495), .SI(\mem3[4][26] ), .SE(test_se), 
        .CLK(n2063), .Q(\mem3[4][27] ), .QN(n29661) );
  SDFFX1 \mem3_reg[4][26]  ( .D(n12494), .SI(\mem3[4][25] ), .SE(test_se), 
        .CLK(n2063), .Q(\mem3[4][26] ), .QN(n29662) );
  SDFFX1 \mem3_reg[4][25]  ( .D(n12493), .SI(\mem3[4][24] ), .SE(test_se), 
        .CLK(n2063), .Q(\mem3[4][25] ), .QN(n29663) );
  SDFFX1 \mem3_reg[4][24]  ( .D(n12492), .SI(\mem3[3][31] ), .SE(test_se), 
        .CLK(n2063), .Q(\mem3[4][24] ), .QN(n29664) );
  SDFFX1 \mem3_reg[3][31]  ( .D(n12491), .SI(\mem3[3][30] ), .SE(test_se), 
        .CLK(n2069), .Q(\mem3[3][31] ), .QN(n29665) );
  SDFFX1 \mem3_reg[3][30]  ( .D(n12490), .SI(\mem3[3][29] ), .SE(test_se), 
        .CLK(n2069), .Q(\mem3[3][30] ), .QN(n29666) );
  SDFFX1 \mem3_reg[3][29]  ( .D(n12489), .SI(\mem3[3][28] ), .SE(test_se), 
        .CLK(n2069), .Q(\mem3[3][29] ), .QN(n29667) );
  SDFFX1 \mem3_reg[3][28]  ( .D(n12488), .SI(\mem3[3][27] ), .SE(test_se), 
        .CLK(n2069), .Q(\mem3[3][28] ), .QN(n29668) );
  SDFFX1 \mem3_reg[3][27]  ( .D(n12487), .SI(\mem3[3][26] ), .SE(test_se), 
        .CLK(n2069), .Q(\mem3[3][27] ), .QN(n29669) );
  SDFFX1 \mem3_reg[3][26]  ( .D(n12486), .SI(\mem3[3][25] ), .SE(test_se), 
        .CLK(n2069), .Q(\mem3[3][26] ), .QN(n29670) );
  SDFFX1 \mem3_reg[3][25]  ( .D(n12485), .SI(\mem3[3][24] ), .SE(test_se), 
        .CLK(n2069), .Q(\mem3[3][25] ), .QN(n29671) );
  SDFFX1 \mem3_reg[3][24]  ( .D(n12484), .SI(\mem3[2][31] ), .SE(test_se), 
        .CLK(n2069), .Q(\mem3[3][24] ), .QN(n29672) );
  SDFFX1 \mem3_reg[2][31]  ( .D(n12483), .SI(\mem3[2][30] ), .SE(test_se), 
        .CLK(n2069), .Q(\mem3[2][31] ), .QN(n29673) );
  SDFFX1 \mem3_reg[2][30]  ( .D(n12482), .SI(\mem3[2][29] ), .SE(test_se), 
        .CLK(n2069), .Q(\mem3[2][30] ), .QN(n29674) );
  SDFFX1 \mem3_reg[2][29]  ( .D(n12481), .SI(\mem3[2][28] ), .SE(test_se), 
        .CLK(n2069), .Q(\mem3[2][29] ), .QN(n29675) );
  SDFFX1 \mem3_reg[2][28]  ( .D(n12480), .SI(\mem3[2][27] ), .SE(test_se), 
        .CLK(n2069), .Q(\mem3[2][28] ), .QN(n29676) );
  SDFFX1 \mem3_reg[2][27]  ( .D(n12479), .SI(\mem3[2][26] ), .SE(test_se), 
        .CLK(n2070), .Q(\mem3[2][27] ), .QN(n29677) );
  SDFFX1 \mem3_reg[2][26]  ( .D(n12478), .SI(\mem3[2][25] ), .SE(test_se), 
        .CLK(n2070), .Q(\mem3[2][26] ), .QN(n29678) );
  SDFFX1 \mem3_reg[2][25]  ( .D(n12477), .SI(\mem3[2][24] ), .SE(test_se), 
        .CLK(n2070), .Q(\mem3[2][25] ), .QN(n29679) );
  SDFFX1 \mem3_reg[2][24]  ( .D(n12476), .SI(\mem3[1][31] ), .SE(test_se), 
        .CLK(n2070), .Q(\mem3[2][24] ), .QN(n29680) );
  SDFFX1 \mem3_reg[1][31]  ( .D(n12475), .SI(\mem3[1][30] ), .SE(test_se), 
        .CLK(n2070), .Q(\mem3[1][31] ), .QN(n29681) );
  SDFFX1 \mem3_reg[1][30]  ( .D(n12474), .SI(\mem3[1][29] ), .SE(test_se), 
        .CLK(n2070), .Q(\mem3[1][30] ), .QN(n29682) );
  SDFFX1 \mem3_reg[1][29]  ( .D(n12473), .SI(\mem3[1][28] ), .SE(test_se), 
        .CLK(n2070), .Q(\mem3[1][29] ), .QN(n29683) );
  SDFFX1 \mem3_reg[1][28]  ( .D(n12472), .SI(\mem3[1][27] ), .SE(test_se), 
        .CLK(n2070), .Q(\mem3[1][28] ), .QN(n29684) );
  SDFFX1 \mem3_reg[1][27]  ( .D(n12471), .SI(\mem3[1][26] ), .SE(test_se), 
        .CLK(n2070), .Q(\mem3[1][27] ), .QN(n29685) );
  SDFFX1 \mem3_reg[1][26]  ( .D(n12470), .SI(\mem3[1][25] ), .SE(test_se), 
        .CLK(n2070), .Q(\mem3[1][26] ), .QN(n29686) );
  SDFFX1 \mem3_reg[1][25]  ( .D(n12469), .SI(\mem3[1][24] ), .SE(test_se), 
        .CLK(n2070), .Q(\mem3[1][25] ), .QN(n29687) );
  SDFFX1 \mem3_reg[1][24]  ( .D(n12468), .SI(\mem3[0][31] ), .SE(test_se), 
        .CLK(n2070), .Q(\mem3[1][24] ), .QN(n29688) );
  SDFFX1 \mem3_reg[0][31]  ( .D(n12467), .SI(\mem3[0][30] ), .SE(test_se), 
        .CLK(n2071), .Q(\mem3[0][31] ), .QN(n29689) );
  SDFFX1 \mem3_reg[0][30]  ( .D(n12466), .SI(\mem3[0][29] ), .SE(test_se), 
        .CLK(n2076), .Q(\mem3[0][30] ), .QN(n29690) );
  SDFFX1 \mem3_reg[0][29]  ( .D(n12465), .SI(\mem3[0][28] ), .SE(test_se), 
        .CLK(n2071), .Q(\mem3[0][29] ), .QN(n29691) );
  SDFFX1 \mem3_reg[0][28]  ( .D(n12464), .SI(\mem3[0][27] ), .SE(test_se), 
        .CLK(n2071), .Q(\mem3[0][28] ), .QN(n29692) );
  SDFFX1 \mem3_reg[0][27]  ( .D(n12463), .SI(\mem3[0][26] ), .SE(test_se), 
        .CLK(n2071), .Q(\mem3[0][27] ), .QN(n29693) );
  SDFFX1 \mem3_reg[0][26]  ( .D(n12462), .SI(\mem3[0][25] ), .SE(test_se), 
        .CLK(n2071), .Q(\mem3[0][26] ), .QN(n29694) );
  SDFFX1 \mem3_reg[0][25]  ( .D(n12461), .SI(\mem3[0][24] ), .SE(test_se), 
        .CLK(n2071), .Q(\mem3[0][25] ), .QN(n29695) );
  SDFFX1 \mem3_reg[0][24]  ( .D(n12460), .SI(\mem2[255][23] ), .SE(test_se), 
        .CLK(n2071), .Q(\mem3[0][24] ), .QN(n29696) );
  SDFFX1 \mem2_reg[255][23]  ( .D(n12459), .SI(\mem2[255][22] ), .SE(test_se), 
        .CLK(n2076), .Q(\mem2[255][23] ), .QN(n29697) );
  SDFFX1 \mem2_reg[255][22]  ( .D(n12458), .SI(\mem2[255][21] ), .SE(test_se), 
        .CLK(n1884), .Q(\mem2[255][22] ), .QN(n29698) );
  SDFFX1 \mem2_reg[255][21]  ( .D(n12457), .SI(\mem2[255][20] ), .SE(test_se), 
        .CLK(n1884), .Q(\mem2[255][21] ), .QN(n29699) );
  SDFFX1 \mem2_reg[255][20]  ( .D(n12456), .SI(\mem2[255][19] ), .SE(test_se), 
        .CLK(n1884), .Q(\mem2[255][20] ), .QN(n29700) );
  SDFFX1 \mem2_reg[255][19]  ( .D(n12455), .SI(\mem2[255][18] ), .SE(test_se), 
        .CLK(n1884), .Q(\mem2[255][19] ), .QN(n29701) );
  SDFFX1 \mem2_reg[255][18]  ( .D(n12454), .SI(\mem2[255][17] ), .SE(test_se), 
        .CLK(n1884), .Q(\mem2[255][18] ), .QN(n29702) );
  SDFFX1 \mem2_reg[255][17]  ( .D(n12453), .SI(\mem2[255][16] ), .SE(test_se), 
        .CLK(n1885), .Q(\mem2[255][17] ), .QN(n29703) );
  SDFFX1 \mem2_reg[255][16]  ( .D(n12452), .SI(\mem2[254][23] ), .SE(test_se), 
        .CLK(n1885), .Q(\mem2[255][16] ), .QN(n29704) );
  SDFFX1 \mem2_reg[254][23]  ( .D(n12451), .SI(\mem2[254][22] ), .SE(test_se), 
        .CLK(n1885), .Q(\mem2[254][23] ), .QN(n29705) );
  SDFFX1 \mem2_reg[254][22]  ( .D(n12450), .SI(\mem2[254][21] ), .SE(test_se), 
        .CLK(n1885), .Q(\mem2[254][22] ), .QN(n29706) );
  SDFFX1 \mem2_reg[254][21]  ( .D(n12449), .SI(\mem2[254][20] ), .SE(test_se), 
        .CLK(n1885), .Q(\mem2[254][21] ), .QN(n29707) );
  SDFFX1 \mem2_reg[254][20]  ( .D(n12448), .SI(\mem2[254][19] ), .SE(test_se), 
        .CLK(n1885), .Q(\mem2[254][20] ), .QN(n29708) );
  SDFFX1 \mem2_reg[254][19]  ( .D(n12447), .SI(\mem2[254][18] ), .SE(test_se), 
        .CLK(n1885), .Q(\mem2[254][19] ), .QN(n29709) );
  SDFFX1 \mem2_reg[254][18]  ( .D(n12446), .SI(\mem2[254][17] ), .SE(test_se), 
        .CLK(n1885), .Q(\mem2[254][18] ), .QN(n29710) );
  SDFFX1 \mem2_reg[254][17]  ( .D(n12445), .SI(\mem2[254][16] ), .SE(test_se), 
        .CLK(n1885), .Q(\mem2[254][17] ), .QN(n29711) );
  SDFFX1 \mem2_reg[254][16]  ( .D(n12444), .SI(\mem2[253][23] ), .SE(test_se), 
        .CLK(n1885), .Q(\mem2[254][16] ), .QN(n29712) );
  SDFFX1 \mem2_reg[253][23]  ( .D(n12443), .SI(\mem2[253][22] ), .SE(test_se), 
        .CLK(n1885), .Q(\mem2[253][23] ), .QN(n29713) );
  SDFFX1 \mem2_reg[253][22]  ( .D(n12442), .SI(\mem2[253][21] ), .SE(test_se), 
        .CLK(n1885), .Q(\mem2[253][22] ), .QN(n29714) );
  SDFFX1 \mem2_reg[253][21]  ( .D(n12441), .SI(\mem2[253][20] ), .SE(test_se), 
        .CLK(n1886), .Q(\mem2[253][21] ), .QN(n29715) );
  SDFFX1 \mem2_reg[253][20]  ( .D(n12440), .SI(\mem2[253][19] ), .SE(test_se), 
        .CLK(n1886), .Q(\mem2[253][20] ), .QN(n29716) );
  SDFFX1 \mem2_reg[253][19]  ( .D(n12439), .SI(\mem2[253][18] ), .SE(test_se), 
        .CLK(n1886), .Q(\mem2[253][19] ), .QN(n29717) );
  SDFFX1 \mem2_reg[253][18]  ( .D(n12438), .SI(\mem2[253][17] ), .SE(test_se), 
        .CLK(n1886), .Q(\mem2[253][18] ), .QN(n29718) );
  SDFFX1 \mem2_reg[253][17]  ( .D(n12437), .SI(\mem2[253][16] ), .SE(test_se), 
        .CLK(n1886), .Q(\mem2[253][17] ), .QN(n29719) );
  SDFFX1 \mem2_reg[253][16]  ( .D(n12436), .SI(\mem2[252][23] ), .SE(test_se), 
        .CLK(n1886), .Q(\mem2[253][16] ), .QN(n29720) );
  SDFFX1 \mem2_reg[252][23]  ( .D(n12435), .SI(\mem2[252][22] ), .SE(test_se), 
        .CLK(n1886), .Q(\mem2[252][23] ), .QN(n29721) );
  SDFFX1 \mem2_reg[252][22]  ( .D(n12434), .SI(\mem2[252][21] ), .SE(test_se), 
        .CLK(n1886), .Q(\mem2[252][22] ), .QN(n29722) );
  SDFFX1 \mem2_reg[252][21]  ( .D(n12433), .SI(\mem2[252][20] ), .SE(test_se), 
        .CLK(n1886), .Q(\mem2[252][21] ), .QN(n29723) );
  SDFFX1 \mem2_reg[252][20]  ( .D(n12432), .SI(\mem2[252][19] ), .SE(test_se), 
        .CLK(n1886), .Q(\mem2[252][20] ), .QN(n29724) );
  SDFFX1 \mem2_reg[252][19]  ( .D(n12431), .SI(\mem2[252][18] ), .SE(test_se), 
        .CLK(n1886), .Q(\mem2[252][19] ), .QN(n29725) );
  SDFFX1 \mem2_reg[252][18]  ( .D(n12430), .SI(\mem2[252][17] ), .SE(test_se), 
        .CLK(n1886), .Q(\mem2[252][18] ), .QN(n29726) );
  SDFFX1 \mem2_reg[252][17]  ( .D(n12429), .SI(\mem2[252][16] ), .SE(test_se), 
        .CLK(n1887), .Q(\mem2[252][17] ), .QN(n29727) );
  SDFFX1 \mem2_reg[252][16]  ( .D(n12428), .SI(\mem2[251][23] ), .SE(test_se), 
        .CLK(n1887), .Q(\mem2[252][16] ), .QN(n29728) );
  SDFFX1 \mem2_reg[251][23]  ( .D(n12427), .SI(\mem2[251][22] ), .SE(test_se), 
        .CLK(n1887), .Q(\mem2[251][23] ), .QN(n29729) );
  SDFFX1 \mem2_reg[251][22]  ( .D(n12426), .SI(\mem2[251][21] ), .SE(test_se), 
        .CLK(n1887), .Q(\mem2[251][22] ), .QN(n29730) );
  SDFFX1 \mem2_reg[251][21]  ( .D(n12425), .SI(\mem2[251][20] ), .SE(test_se), 
        .CLK(n1887), .Q(\mem2[251][21] ), .QN(n29731) );
  SDFFX1 \mem2_reg[251][20]  ( .D(n12424), .SI(\mem2[251][19] ), .SE(test_se), 
        .CLK(n1887), .Q(\mem2[251][20] ), .QN(n29732) );
  SDFFX1 \mem2_reg[251][19]  ( .D(n12423), .SI(\mem2[251][18] ), .SE(test_se), 
        .CLK(n1887), .Q(\mem2[251][19] ), .QN(n29733) );
  SDFFX1 \mem2_reg[251][18]  ( .D(n12422), .SI(\mem2[251][17] ), .SE(test_se), 
        .CLK(n1887), .Q(\mem2[251][18] ), .QN(n29734) );
  SDFFX1 \mem2_reg[251][17]  ( .D(n12421), .SI(\mem2[251][16] ), .SE(test_se), 
        .CLK(n1887), .Q(\mem2[251][17] ), .QN(n29735) );
  SDFFX1 \mem2_reg[251][16]  ( .D(n12420), .SI(\mem2[250][23] ), .SE(test_se), 
        .CLK(n1887), .Q(\mem2[251][16] ), .QN(n29736) );
  SDFFX1 \mem2_reg[250][23]  ( .D(n12419), .SI(\mem2[250][22] ), .SE(test_se), 
        .CLK(n1887), .Q(\mem2[250][23] ), .QN(n29737) );
  SDFFX1 \mem2_reg[250][22]  ( .D(n12418), .SI(\mem2[250][21] ), .SE(test_se), 
        .CLK(n1887), .Q(\mem2[250][22] ), .QN(n29738) );
  SDFFX1 \mem2_reg[250][21]  ( .D(n12417), .SI(\mem2[250][20] ), .SE(test_se), 
        .CLK(n1888), .Q(\mem2[250][21] ), .QN(n29739) );
  SDFFX1 \mem2_reg[250][20]  ( .D(n12416), .SI(\mem2[250][19] ), .SE(test_se), 
        .CLK(n1888), .Q(\mem2[250][20] ), .QN(n29740) );
  SDFFX1 \mem2_reg[250][19]  ( .D(n12415), .SI(\mem2[250][18] ), .SE(test_se), 
        .CLK(n1888), .Q(\mem2[250][19] ), .QN(n29741) );
  SDFFX1 \mem2_reg[250][18]  ( .D(n12414), .SI(\mem2[250][17] ), .SE(test_se), 
        .CLK(n1888), .Q(\mem2[250][18] ), .QN(n29742) );
  SDFFX1 \mem2_reg[250][17]  ( .D(n12413), .SI(\mem2[250][16] ), .SE(test_se), 
        .CLK(n1888), .Q(\mem2[250][17] ), .QN(n29743) );
  SDFFX1 \mem2_reg[250][16]  ( .D(n12412), .SI(\mem2[249][23] ), .SE(test_se), 
        .CLK(n1888), .Q(\mem2[250][16] ), .QN(n29744) );
  SDFFX1 \mem2_reg[249][23]  ( .D(n12411), .SI(\mem2[249][22] ), .SE(test_se), 
        .CLK(n1888), .Q(\mem2[249][23] ), .QN(n29745) );
  SDFFX1 \mem2_reg[249][22]  ( .D(n12410), .SI(\mem2[249][21] ), .SE(test_se), 
        .CLK(n1888), .Q(\mem2[249][22] ), .QN(n29746) );
  SDFFX1 \mem2_reg[249][21]  ( .D(n12409), .SI(\mem2[249][20] ), .SE(test_se), 
        .CLK(n1888), .Q(\mem2[249][21] ), .QN(n29747) );
  SDFFX1 \mem2_reg[249][20]  ( .D(n12408), .SI(\mem2[249][19] ), .SE(test_se), 
        .CLK(n1888), .Q(\mem2[249][20] ), .QN(n29748) );
  SDFFX1 \mem2_reg[249][19]  ( .D(n12407), .SI(\mem2[249][18] ), .SE(test_se), 
        .CLK(n1888), .Q(\mem2[249][19] ), .QN(n29749) );
  SDFFX1 \mem2_reg[249][18]  ( .D(n12406), .SI(\mem2[249][17] ), .SE(test_se), 
        .CLK(n1888), .Q(\mem2[249][18] ), .QN(n29750) );
  SDFFX1 \mem2_reg[249][17]  ( .D(n12405), .SI(\mem2[249][16] ), .SE(test_se), 
        .CLK(n1889), .Q(\mem2[249][17] ), .QN(n29751) );
  SDFFX1 \mem2_reg[249][16]  ( .D(n12404), .SI(\mem2[248][23] ), .SE(test_se), 
        .CLK(n1889), .Q(\mem2[249][16] ), .QN(n29752) );
  SDFFX1 \mem2_reg[248][23]  ( .D(n12403), .SI(\mem2[248][22] ), .SE(test_se), 
        .CLK(n1889), .Q(\mem2[248][23] ), .QN(n29753) );
  SDFFX1 \mem2_reg[248][22]  ( .D(n12402), .SI(\mem2[248][21] ), .SE(test_se), 
        .CLK(n1889), .Q(\mem2[248][22] ), .QN(n29754) );
  SDFFX1 \mem2_reg[248][21]  ( .D(n12401), .SI(\mem2[248][20] ), .SE(test_se), 
        .CLK(n1889), .Q(\mem2[248][21] ), .QN(n29755) );
  SDFFX1 \mem2_reg[248][20]  ( .D(n12400), .SI(\mem2[248][19] ), .SE(test_se), 
        .CLK(n1889), .Q(\mem2[248][20] ), .QN(n29756) );
  SDFFX1 \mem2_reg[248][19]  ( .D(n12399), .SI(\mem2[248][18] ), .SE(test_se), 
        .CLK(n1889), .Q(\mem2[248][19] ), .QN(n29757) );
  SDFFX1 \mem2_reg[248][18]  ( .D(n12398), .SI(\mem2[248][17] ), .SE(test_se), 
        .CLK(n1889), .Q(\mem2[248][18] ), .QN(n29758) );
  SDFFX1 \mem2_reg[248][17]  ( .D(n12397), .SI(\mem2[248][16] ), .SE(test_se), 
        .CLK(n1889), .Q(\mem2[248][17] ), .QN(n29759) );
  SDFFX1 \mem2_reg[248][16]  ( .D(n12396), .SI(\mem2[247][23] ), .SE(test_se), 
        .CLK(n1889), .Q(\mem2[248][16] ), .QN(n29760) );
  SDFFX1 \mem2_reg[247][23]  ( .D(n12395), .SI(\mem2[247][22] ), .SE(test_se), 
        .CLK(n1889), .Q(\mem2[247][23] ), .QN(n29761) );
  SDFFX1 \mem2_reg[247][22]  ( .D(n12394), .SI(\mem2[247][21] ), .SE(test_se), 
        .CLK(n1889), .Q(\mem2[247][22] ), .QN(n29762) );
  SDFFX1 \mem2_reg[247][21]  ( .D(n12393), .SI(\mem2[247][20] ), .SE(test_se), 
        .CLK(n1890), .Q(\mem2[247][21] ), .QN(n29763) );
  SDFFX1 \mem2_reg[247][20]  ( .D(n12392), .SI(\mem2[247][19] ), .SE(test_se), 
        .CLK(n1890), .Q(\mem2[247][20] ), .QN(n29764) );
  SDFFX1 \mem2_reg[247][19]  ( .D(n12391), .SI(\mem2[247][18] ), .SE(test_se), 
        .CLK(n1890), .Q(\mem2[247][19] ), .QN(n29765) );
  SDFFX1 \mem2_reg[247][18]  ( .D(n12390), .SI(\mem2[247][17] ), .SE(test_se), 
        .CLK(n1890), .Q(\mem2[247][18] ), .QN(n29766) );
  SDFFX1 \mem2_reg[247][17]  ( .D(n12389), .SI(\mem2[247][16] ), .SE(test_se), 
        .CLK(n1890), .Q(\mem2[247][17] ), .QN(n29767) );
  SDFFX1 \mem2_reg[247][16]  ( .D(n12388), .SI(\mem2[246][23] ), .SE(test_se), 
        .CLK(n1890), .Q(\mem2[247][16] ), .QN(n29768) );
  SDFFX1 \mem2_reg[246][23]  ( .D(n12387), .SI(\mem2[246][22] ), .SE(test_se), 
        .CLK(n1890), .Q(\mem2[246][23] ), .QN(n29769) );
  SDFFX1 \mem2_reg[246][22]  ( .D(n12386), .SI(\mem2[246][21] ), .SE(test_se), 
        .CLK(n1890), .Q(\mem2[246][22] ), .QN(n29770) );
  SDFFX1 \mem2_reg[246][21]  ( .D(n12385), .SI(\mem2[246][20] ), .SE(test_se), 
        .CLK(n1890), .Q(\mem2[246][21] ), .QN(n29771) );
  SDFFX1 \mem2_reg[246][20]  ( .D(n12384), .SI(\mem2[246][19] ), .SE(test_se), 
        .CLK(n1890), .Q(\mem2[246][20] ), .QN(n29772) );
  SDFFX1 \mem2_reg[246][19]  ( .D(n12383), .SI(\mem2[246][18] ), .SE(test_se), 
        .CLK(n1890), .Q(\mem2[246][19] ), .QN(n29773) );
  SDFFX1 \mem2_reg[246][18]  ( .D(n12382), .SI(\mem2[246][17] ), .SE(test_se), 
        .CLK(n1890), .Q(\mem2[246][18] ), .QN(n29774) );
  SDFFX1 \mem2_reg[246][17]  ( .D(n12381), .SI(\mem2[246][16] ), .SE(test_se), 
        .CLK(n1891), .Q(\mem2[246][17] ), .QN(n29775) );
  SDFFX1 \mem2_reg[246][16]  ( .D(n12380), .SI(\mem2[245][23] ), .SE(test_se), 
        .CLK(n1891), .Q(\mem2[246][16] ), .QN(n29776) );
  SDFFX1 \mem2_reg[245][23]  ( .D(n12379), .SI(\mem2[245][22] ), .SE(test_se), 
        .CLK(n1891), .Q(\mem2[245][23] ), .QN(n29777) );
  SDFFX1 \mem2_reg[245][22]  ( .D(n12378), .SI(\mem2[245][21] ), .SE(test_se), 
        .CLK(n1891), .Q(\mem2[245][22] ), .QN(n29778) );
  SDFFX1 \mem2_reg[245][21]  ( .D(n12377), .SI(\mem2[245][20] ), .SE(test_se), 
        .CLK(n1891), .Q(\mem2[245][21] ), .QN(n29779) );
  SDFFX1 \mem2_reg[245][20]  ( .D(n12376), .SI(\mem2[245][19] ), .SE(test_se), 
        .CLK(n1891), .Q(\mem2[245][20] ), .QN(n29780) );
  SDFFX1 \mem2_reg[245][19]  ( .D(n12375), .SI(\mem2[245][18] ), .SE(test_se), 
        .CLK(n1891), .Q(\mem2[245][19] ), .QN(n29781) );
  SDFFX1 \mem2_reg[245][18]  ( .D(n12374), .SI(\mem2[245][17] ), .SE(test_se), 
        .CLK(n1891), .Q(\mem2[245][18] ), .QN(n29782) );
  SDFFX1 \mem2_reg[245][17]  ( .D(n12373), .SI(\mem2[245][16] ), .SE(test_se), 
        .CLK(n1891), .Q(\mem2[245][17] ), .QN(n29783) );
  SDFFX1 \mem2_reg[245][16]  ( .D(n12372), .SI(\mem2[244][23] ), .SE(test_se), 
        .CLK(n1891), .Q(\mem2[245][16] ), .QN(n29784) );
  SDFFX1 \mem2_reg[244][23]  ( .D(n12371), .SI(\mem2[244][22] ), .SE(test_se), 
        .CLK(n1891), .Q(\mem2[244][23] ), .QN(n29785) );
  SDFFX1 \mem2_reg[244][22]  ( .D(n12370), .SI(\mem2[244][21] ), .SE(test_se), 
        .CLK(n1891), .Q(\mem2[244][22] ), .QN(n29786) );
  SDFFX1 \mem2_reg[244][21]  ( .D(n12369), .SI(\mem2[244][20] ), .SE(test_se), 
        .CLK(n1892), .Q(\mem2[244][21] ), .QN(n29787) );
  SDFFX1 \mem2_reg[244][20]  ( .D(n12368), .SI(\mem2[244][19] ), .SE(test_se), 
        .CLK(n1892), .Q(\mem2[244][20] ), .QN(n29788) );
  SDFFX1 \mem2_reg[244][19]  ( .D(n12367), .SI(\mem2[244][18] ), .SE(test_se), 
        .CLK(n1892), .Q(\mem2[244][19] ), .QN(n29789) );
  SDFFX1 \mem2_reg[244][18]  ( .D(n12366), .SI(\mem2[244][17] ), .SE(test_se), 
        .CLK(n1892), .Q(\mem2[244][18] ), .QN(n29790) );
  SDFFX1 \mem2_reg[244][17]  ( .D(n12365), .SI(\mem2[244][16] ), .SE(test_se), 
        .CLK(n1892), .Q(\mem2[244][17] ), .QN(n29791) );
  SDFFX1 \mem2_reg[244][16]  ( .D(n12364), .SI(\mem2[243][23] ), .SE(test_se), 
        .CLK(n1892), .Q(\mem2[244][16] ), .QN(n29792) );
  SDFFX1 \mem2_reg[243][23]  ( .D(n12363), .SI(\mem2[243][22] ), .SE(test_se), 
        .CLK(n1892), .Q(\mem2[243][23] ), .QN(n29793) );
  SDFFX1 \mem2_reg[243][22]  ( .D(n12362), .SI(\mem2[243][21] ), .SE(test_se), 
        .CLK(n1892), .Q(\mem2[243][22] ), .QN(n29794) );
  SDFFX1 \mem2_reg[243][21]  ( .D(n12361), .SI(\mem2[243][20] ), .SE(test_se), 
        .CLK(n1892), .Q(\mem2[243][21] ), .QN(n29795) );
  SDFFX1 \mem2_reg[243][20]  ( .D(n12360), .SI(\mem2[243][19] ), .SE(test_se), 
        .CLK(n1892), .Q(\mem2[243][20] ), .QN(n29796) );
  SDFFX1 \mem2_reg[243][19]  ( .D(n12359), .SI(\mem2[243][18] ), .SE(test_se), 
        .CLK(n1892), .Q(\mem2[243][19] ), .QN(n29797) );
  SDFFX1 \mem2_reg[243][18]  ( .D(n12358), .SI(\mem2[243][17] ), .SE(test_se), 
        .CLK(n1892), .Q(\mem2[243][18] ), .QN(n29798) );
  SDFFX1 \mem2_reg[243][17]  ( .D(n12357), .SI(\mem2[243][16] ), .SE(test_se), 
        .CLK(n1893), .Q(\mem2[243][17] ), .QN(n29799) );
  SDFFX1 \mem2_reg[243][16]  ( .D(n12356), .SI(\mem2[242][23] ), .SE(test_se), 
        .CLK(n1893), .Q(\mem2[243][16] ), .QN(n29800) );
  SDFFX1 \mem2_reg[242][23]  ( .D(n12355), .SI(\mem2[242][22] ), .SE(test_se), 
        .CLK(n1893), .Q(\mem2[242][23] ), .QN(n29801) );
  SDFFX1 \mem2_reg[242][22]  ( .D(n12354), .SI(\mem2[242][21] ), .SE(test_se), 
        .CLK(n1893), .Q(\mem2[242][22] ), .QN(n29802) );
  SDFFX1 \mem2_reg[242][21]  ( .D(n12353), .SI(\mem2[242][20] ), .SE(test_se), 
        .CLK(n1893), .Q(\mem2[242][21] ), .QN(n29803) );
  SDFFX1 \mem2_reg[242][20]  ( .D(n12352), .SI(\mem2[242][19] ), .SE(test_se), 
        .CLK(n1893), .Q(\mem2[242][20] ), .QN(n29804) );
  SDFFX1 \mem2_reg[242][19]  ( .D(n12351), .SI(\mem2[242][18] ), .SE(test_se), 
        .CLK(n1893), .Q(\mem2[242][19] ), .QN(n29805) );
  SDFFX1 \mem2_reg[242][18]  ( .D(n12350), .SI(\mem2[242][17] ), .SE(test_se), 
        .CLK(n1893), .Q(\mem2[242][18] ), .QN(n29806) );
  SDFFX1 \mem2_reg[242][17]  ( .D(n12349), .SI(\mem2[242][16] ), .SE(test_se), 
        .CLK(n1893), .Q(\mem2[242][17] ), .QN(n29807) );
  SDFFX1 \mem2_reg[242][16]  ( .D(n12348), .SI(\mem2[241][23] ), .SE(test_se), 
        .CLK(n1893), .Q(\mem2[242][16] ), .QN(n29808) );
  SDFFX1 \mem2_reg[241][23]  ( .D(n12347), .SI(\mem2[241][22] ), .SE(test_se), 
        .CLK(n1893), .Q(\mem2[241][23] ), .QN(n29809) );
  SDFFX1 \mem2_reg[241][22]  ( .D(n12346), .SI(\mem2[241][21] ), .SE(test_se), 
        .CLK(n1893), .Q(\mem2[241][22] ), .QN(n29810) );
  SDFFX1 \mem2_reg[241][21]  ( .D(n12345), .SI(\mem2[241][20] ), .SE(test_se), 
        .CLK(n1894), .Q(\mem2[241][21] ), .QN(n29811) );
  SDFFX1 \mem2_reg[241][20]  ( .D(n12344), .SI(\mem2[241][19] ), .SE(test_se), 
        .CLK(n1894), .Q(\mem2[241][20] ), .QN(n29812) );
  SDFFX1 \mem2_reg[241][19]  ( .D(n12343), .SI(\mem2[241][18] ), .SE(test_se), 
        .CLK(n1894), .Q(\mem2[241][19] ), .QN(n29813) );
  SDFFX1 \mem2_reg[241][18]  ( .D(n12342), .SI(\mem2[241][17] ), .SE(test_se), 
        .CLK(n1894), .Q(\mem2[241][18] ), .QN(n29814) );
  SDFFX1 \mem2_reg[241][17]  ( .D(n12341), .SI(\mem2[241][16] ), .SE(test_se), 
        .CLK(n1894), .Q(\mem2[241][17] ), .QN(n29815) );
  SDFFX1 \mem2_reg[241][16]  ( .D(n12340), .SI(\mem2[240][23] ), .SE(test_se), 
        .CLK(n1894), .Q(\mem2[241][16] ), .QN(n29816) );
  SDFFX1 \mem2_reg[240][23]  ( .D(n12339), .SI(\mem2[240][22] ), .SE(test_se), 
        .CLK(n1894), .Q(\mem2[240][23] ), .QN(n29817) );
  SDFFX1 \mem2_reg[240][22]  ( .D(n12338), .SI(\mem2[240][21] ), .SE(test_se), 
        .CLK(n1894), .Q(\mem2[240][22] ), .QN(n29818) );
  SDFFX1 \mem2_reg[240][21]  ( .D(n12337), .SI(\mem2[240][20] ), .SE(test_se), 
        .CLK(n1894), .Q(\mem2[240][21] ), .QN(n29819) );
  SDFFX1 \mem2_reg[240][20]  ( .D(n12336), .SI(\mem2[240][19] ), .SE(test_se), 
        .CLK(n1894), .Q(\mem2[240][20] ), .QN(n29820) );
  SDFFX1 \mem2_reg[240][19]  ( .D(n12335), .SI(\mem2[240][18] ), .SE(test_se), 
        .CLK(n1894), .Q(\mem2[240][19] ), .QN(n29821) );
  SDFFX1 \mem2_reg[240][18]  ( .D(n12334), .SI(\mem2[240][17] ), .SE(test_se), 
        .CLK(n1894), .Q(\mem2[240][18] ), .QN(n29822) );
  SDFFX1 \mem2_reg[240][17]  ( .D(n12333), .SI(\mem2[240][16] ), .SE(test_se), 
        .CLK(n1895), .Q(\mem2[240][17] ), .QN(n29823) );
  SDFFX1 \mem2_reg[240][16]  ( .D(n12332), .SI(\mem2[239][23] ), .SE(test_se), 
        .CLK(n1895), .Q(\mem2[240][16] ), .QN(n29824) );
  SDFFX1 \mem2_reg[239][23]  ( .D(n12331), .SI(\mem2[239][22] ), .SE(test_se), 
        .CLK(n1895), .Q(\mem2[239][23] ), .QN(n29825) );
  SDFFX1 \mem2_reg[239][22]  ( .D(n12330), .SI(\mem2[239][21] ), .SE(test_se), 
        .CLK(n1895), .Q(\mem2[239][22] ), .QN(n29826) );
  SDFFX1 \mem2_reg[239][21]  ( .D(n12329), .SI(\mem2[239][20] ), .SE(test_se), 
        .CLK(n1895), .Q(\mem2[239][21] ), .QN(n29827) );
  SDFFX1 \mem2_reg[239][20]  ( .D(n12328), .SI(\mem2[239][19] ), .SE(test_se), 
        .CLK(n1895), .Q(\mem2[239][20] ), .QN(n29828) );
  SDFFX1 \mem2_reg[239][19]  ( .D(n12327), .SI(\mem2[239][18] ), .SE(test_se), 
        .CLK(n1895), .Q(\mem2[239][19] ), .QN(n29829) );
  SDFFX1 \mem2_reg[239][18]  ( .D(n12326), .SI(\mem2[239][17] ), .SE(test_se), 
        .CLK(n1895), .Q(\mem2[239][18] ), .QN(n29830) );
  SDFFX1 \mem2_reg[239][17]  ( .D(n12325), .SI(\mem2[239][16] ), .SE(test_se), 
        .CLK(n1895), .Q(\mem2[239][17] ), .QN(n29831) );
  SDFFX1 \mem2_reg[239][16]  ( .D(n12324), .SI(\mem2[238][23] ), .SE(test_se), 
        .CLK(n1895), .Q(\mem2[239][16] ), .QN(n29832) );
  SDFFX1 \mem2_reg[238][23]  ( .D(n12323), .SI(\mem2[238][22] ), .SE(test_se), 
        .CLK(n1895), .Q(\mem2[238][23] ), .QN(n29833) );
  SDFFX1 \mem2_reg[238][22]  ( .D(n12322), .SI(\mem2[238][21] ), .SE(test_se), 
        .CLK(n1895), .Q(\mem2[238][22] ), .QN(n29834) );
  SDFFX1 \mem2_reg[238][21]  ( .D(n12321), .SI(\mem2[238][20] ), .SE(test_se), 
        .CLK(n1896), .Q(\mem2[238][21] ), .QN(n29835) );
  SDFFX1 \mem2_reg[238][20]  ( .D(n12320), .SI(\mem2[238][19] ), .SE(test_se), 
        .CLK(n1896), .Q(\mem2[238][20] ), .QN(n29836) );
  SDFFX1 \mem2_reg[238][19]  ( .D(n12319), .SI(\mem2[238][18] ), .SE(test_se), 
        .CLK(n1896), .Q(\mem2[238][19] ), .QN(n29837) );
  SDFFX1 \mem2_reg[238][18]  ( .D(n12318), .SI(\mem2[238][17] ), .SE(test_se), 
        .CLK(n1896), .Q(\mem2[238][18] ), .QN(n29838) );
  SDFFX1 \mem2_reg[238][17]  ( .D(n12317), .SI(\mem2[238][16] ), .SE(test_se), 
        .CLK(n1896), .Q(\mem2[238][17] ), .QN(n29839) );
  SDFFX1 \mem2_reg[238][16]  ( .D(n12316), .SI(\mem2[237][23] ), .SE(test_se), 
        .CLK(n1896), .Q(\mem2[238][16] ), .QN(n29840) );
  SDFFX1 \mem2_reg[237][23]  ( .D(n12315), .SI(\mem2[237][22] ), .SE(test_se), 
        .CLK(n1896), .Q(\mem2[237][23] ), .QN(n29841) );
  SDFFX1 \mem2_reg[237][22]  ( .D(n12314), .SI(\mem2[237][21] ), .SE(test_se), 
        .CLK(n1896), .Q(\mem2[237][22] ), .QN(n29842) );
  SDFFX1 \mem2_reg[237][21]  ( .D(n12313), .SI(\mem2[237][20] ), .SE(test_se), 
        .CLK(n1896), .Q(\mem2[237][21] ), .QN(n29843) );
  SDFFX1 \mem2_reg[237][20]  ( .D(n12312), .SI(\mem2[237][19] ), .SE(test_se), 
        .CLK(n1896), .Q(\mem2[237][20] ), .QN(n29844) );
  SDFFX1 \mem2_reg[237][19]  ( .D(n12311), .SI(\mem2[237][18] ), .SE(test_se), 
        .CLK(n1896), .Q(\mem2[237][19] ), .QN(n29845) );
  SDFFX1 \mem2_reg[237][18]  ( .D(n12310), .SI(\mem2[237][17] ), .SE(test_se), 
        .CLK(n1896), .Q(\mem2[237][18] ), .QN(n29846) );
  SDFFX1 \mem2_reg[237][17]  ( .D(n12309), .SI(\mem2[237][16] ), .SE(test_se), 
        .CLK(n1897), .Q(\mem2[237][17] ), .QN(n29847) );
  SDFFX1 \mem2_reg[237][16]  ( .D(n12308), .SI(\mem2[236][23] ), .SE(test_se), 
        .CLK(n1897), .Q(\mem2[237][16] ), .QN(n29848) );
  SDFFX1 \mem2_reg[236][23]  ( .D(n12307), .SI(\mem2[236][22] ), .SE(test_se), 
        .CLK(n1897), .Q(\mem2[236][23] ), .QN(n29849) );
  SDFFX1 \mem2_reg[236][22]  ( .D(n12306), .SI(\mem2[236][21] ), .SE(test_se), 
        .CLK(n1897), .Q(\mem2[236][22] ), .QN(n29850) );
  SDFFX1 \mem2_reg[236][21]  ( .D(n12305), .SI(\mem2[236][20] ), .SE(test_se), 
        .CLK(n1897), .Q(\mem2[236][21] ), .QN(n29851) );
  SDFFX1 \mem2_reg[236][20]  ( .D(n12304), .SI(\mem2[236][19] ), .SE(test_se), 
        .CLK(n1897), .Q(\mem2[236][20] ), .QN(n29852) );
  SDFFX1 \mem2_reg[236][19]  ( .D(n12303), .SI(\mem2[236][18] ), .SE(test_se), 
        .CLK(n1897), .Q(\mem2[236][19] ), .QN(n29853) );
  SDFFX1 \mem2_reg[236][18]  ( .D(n12302), .SI(\mem2[236][17] ), .SE(test_se), 
        .CLK(n1897), .Q(\mem2[236][18] ), .QN(n29854) );
  SDFFX1 \mem2_reg[236][17]  ( .D(n12301), .SI(\mem2[236][16] ), .SE(test_se), 
        .CLK(n1897), .Q(\mem2[236][17] ), .QN(n29855) );
  SDFFX1 \mem2_reg[236][16]  ( .D(n12300), .SI(\mem2[235][23] ), .SE(test_se), 
        .CLK(n1897), .Q(\mem2[236][16] ), .QN(n29856) );
  SDFFX1 \mem2_reg[235][23]  ( .D(n12299), .SI(\mem2[235][22] ), .SE(test_se), 
        .CLK(n1897), .Q(\mem2[235][23] ), .QN(n29857) );
  SDFFX1 \mem2_reg[235][22]  ( .D(n12298), .SI(\mem2[235][21] ), .SE(test_se), 
        .CLK(n1897), .Q(\mem2[235][22] ), .QN(n29858) );
  SDFFX1 \mem2_reg[235][21]  ( .D(n12297), .SI(\mem2[235][20] ), .SE(test_se), 
        .CLK(n1898), .Q(\mem2[235][21] ), .QN(n29859) );
  SDFFX1 \mem2_reg[235][20]  ( .D(n12296), .SI(\mem2[235][19] ), .SE(test_se), 
        .CLK(n1898), .Q(\mem2[235][20] ), .QN(n29860) );
  SDFFX1 \mem2_reg[235][19]  ( .D(n12295), .SI(\mem2[235][18] ), .SE(test_se), 
        .CLK(n1898), .Q(\mem2[235][19] ), .QN(n29861) );
  SDFFX1 \mem2_reg[235][18]  ( .D(n12294), .SI(\mem2[235][17] ), .SE(test_se), 
        .CLK(n1898), .Q(\mem2[235][18] ), .QN(n29862) );
  SDFFX1 \mem2_reg[235][17]  ( .D(n12293), .SI(\mem2[235][16] ), .SE(test_se), 
        .CLK(n1898), .Q(\mem2[235][17] ), .QN(n29863) );
  SDFFX1 \mem2_reg[235][16]  ( .D(n12292), .SI(\mem2[234][23] ), .SE(test_se), 
        .CLK(n1898), .Q(\mem2[235][16] ), .QN(n29864) );
  SDFFX1 \mem2_reg[234][23]  ( .D(n12291), .SI(\mem2[234][22] ), .SE(test_se), 
        .CLK(n1898), .Q(\mem2[234][23] ), .QN(n29865) );
  SDFFX1 \mem2_reg[234][22]  ( .D(n12290), .SI(\mem2[234][21] ), .SE(test_se), 
        .CLK(n1898), .Q(\mem2[234][22] ), .QN(n29866) );
  SDFFX1 \mem2_reg[234][21]  ( .D(n12289), .SI(\mem2[234][20] ), .SE(test_se), 
        .CLK(n1898), .Q(\mem2[234][21] ), .QN(n29867) );
  SDFFX1 \mem2_reg[234][20]  ( .D(n12288), .SI(\mem2[234][19] ), .SE(test_se), 
        .CLK(n1898), .Q(\mem2[234][20] ), .QN(n29868) );
  SDFFX1 \mem2_reg[234][19]  ( .D(n12287), .SI(\mem2[234][18] ), .SE(test_se), 
        .CLK(n1898), .Q(\mem2[234][19] ), .QN(n29869) );
  SDFFX1 \mem2_reg[234][18]  ( .D(n12286), .SI(\mem2[234][17] ), .SE(test_se), 
        .CLK(n1898), .Q(\mem2[234][18] ), .QN(n29870) );
  SDFFX1 \mem2_reg[234][17]  ( .D(n12285), .SI(\mem2[234][16] ), .SE(test_se), 
        .CLK(n1899), .Q(\mem2[234][17] ), .QN(n29871) );
  SDFFX1 \mem2_reg[234][16]  ( .D(n12284), .SI(\mem2[233][23] ), .SE(test_se), 
        .CLK(n1899), .Q(\mem2[234][16] ), .QN(n29872) );
  SDFFX1 \mem2_reg[233][23]  ( .D(n12283), .SI(\mem2[233][22] ), .SE(test_se), 
        .CLK(n1899), .Q(\mem2[233][23] ), .QN(n29873) );
  SDFFX1 \mem2_reg[233][22]  ( .D(n12282), .SI(\mem2[233][21] ), .SE(test_se), 
        .CLK(n1899), .Q(\mem2[233][22] ), .QN(n29874) );
  SDFFX1 \mem2_reg[233][21]  ( .D(n12281), .SI(\mem2[233][20] ), .SE(test_se), 
        .CLK(n1899), .Q(\mem2[233][21] ), .QN(n29875) );
  SDFFX1 \mem2_reg[233][20]  ( .D(n12280), .SI(\mem2[233][19] ), .SE(test_se), 
        .CLK(n1899), .Q(\mem2[233][20] ), .QN(n29876) );
  SDFFX1 \mem2_reg[233][19]  ( .D(n12279), .SI(\mem2[233][18] ), .SE(test_se), 
        .CLK(n1899), .Q(\mem2[233][19] ), .QN(n29877) );
  SDFFX1 \mem2_reg[233][18]  ( .D(n12278), .SI(\mem2[233][17] ), .SE(test_se), 
        .CLK(n1899), .Q(\mem2[233][18] ), .QN(n29878) );
  SDFFX1 \mem2_reg[233][17]  ( .D(n12277), .SI(\mem2[233][16] ), .SE(test_se), 
        .CLK(n1899), .Q(\mem2[233][17] ), .QN(n29879) );
  SDFFX1 \mem2_reg[233][16]  ( .D(n12276), .SI(\mem2[232][23] ), .SE(test_se), 
        .CLK(n1899), .Q(\mem2[233][16] ), .QN(n29880) );
  SDFFX1 \mem2_reg[232][23]  ( .D(n12275), .SI(\mem2[232][22] ), .SE(test_se), 
        .CLK(n1899), .Q(\mem2[232][23] ), .QN(n29881) );
  SDFFX1 \mem2_reg[232][22]  ( .D(n12274), .SI(\mem2[232][21] ), .SE(test_se), 
        .CLK(n1899), .Q(\mem2[232][22] ), .QN(n29882) );
  SDFFX1 \mem2_reg[232][21]  ( .D(n12273), .SI(\mem2[232][20] ), .SE(test_se), 
        .CLK(n1900), .Q(\mem2[232][21] ), .QN(n29883) );
  SDFFX1 \mem2_reg[232][20]  ( .D(n12272), .SI(\mem2[232][19] ), .SE(test_se), 
        .CLK(n1900), .Q(\mem2[232][20] ), .QN(n29884) );
  SDFFX1 \mem2_reg[232][19]  ( .D(n12271), .SI(\mem2[232][18] ), .SE(test_se), 
        .CLK(n1900), .Q(\mem2[232][19] ), .QN(n29885) );
  SDFFX1 \mem2_reg[232][18]  ( .D(n12270), .SI(\mem2[232][17] ), .SE(test_se), 
        .CLK(n1900), .Q(\mem2[232][18] ), .QN(n29886) );
  SDFFX1 \mem2_reg[232][17]  ( .D(n12269), .SI(\mem2[232][16] ), .SE(test_se), 
        .CLK(n1900), .Q(\mem2[232][17] ), .QN(n29887) );
  SDFFX1 \mem2_reg[232][16]  ( .D(n12268), .SI(\mem2[231][23] ), .SE(test_se), 
        .CLK(n1900), .Q(\mem2[232][16] ), .QN(n29888) );
  SDFFX1 \mem2_reg[231][23]  ( .D(n12267), .SI(\mem2[231][22] ), .SE(test_se), 
        .CLK(n1900), .Q(\mem2[231][23] ), .QN(n29889) );
  SDFFX1 \mem2_reg[231][22]  ( .D(n12266), .SI(\mem2[231][21] ), .SE(test_se), 
        .CLK(n1900), .Q(\mem2[231][22] ), .QN(n29890) );
  SDFFX1 \mem2_reg[231][21]  ( .D(n12265), .SI(\mem2[231][20] ), .SE(test_se), 
        .CLK(n1900), .Q(\mem2[231][21] ), .QN(n29891) );
  SDFFX1 \mem2_reg[231][20]  ( .D(n12264), .SI(\mem2[231][19] ), .SE(test_se), 
        .CLK(n1900), .Q(\mem2[231][20] ), .QN(n29892) );
  SDFFX1 \mem2_reg[231][19]  ( .D(n12263), .SI(\mem2[231][18] ), .SE(test_se), 
        .CLK(n1900), .Q(\mem2[231][19] ), .QN(n29893) );
  SDFFX1 \mem2_reg[231][18]  ( .D(n12262), .SI(\mem2[231][17] ), .SE(test_se), 
        .CLK(n1900), .Q(\mem2[231][18] ), .QN(n29894) );
  SDFFX1 \mem2_reg[231][17]  ( .D(n12261), .SI(\mem2[231][16] ), .SE(test_se), 
        .CLK(n1901), .Q(\mem2[231][17] ), .QN(n29895) );
  SDFFX1 \mem2_reg[231][16]  ( .D(n12260), .SI(\mem2[230][23] ), .SE(test_se), 
        .CLK(n1901), .Q(\mem2[231][16] ), .QN(n29896) );
  SDFFX1 \mem2_reg[230][23]  ( .D(n12259), .SI(\mem2[230][22] ), .SE(test_se), 
        .CLK(n1901), .Q(\mem2[230][23] ), .QN(n29897) );
  SDFFX1 \mem2_reg[230][22]  ( .D(n12258), .SI(\mem2[230][21] ), .SE(test_se), 
        .CLK(n1901), .Q(\mem2[230][22] ), .QN(n29898) );
  SDFFX1 \mem2_reg[230][21]  ( .D(n12257), .SI(\mem2[230][20] ), .SE(test_se), 
        .CLK(n1901), .Q(\mem2[230][21] ), .QN(n29899) );
  SDFFX1 \mem2_reg[230][20]  ( .D(n12256), .SI(\mem2[230][19] ), .SE(test_se), 
        .CLK(n1901), .Q(\mem2[230][20] ), .QN(n29900) );
  SDFFX1 \mem2_reg[230][19]  ( .D(n12255), .SI(\mem2[230][18] ), .SE(test_se), 
        .CLK(n1901), .Q(\mem2[230][19] ), .QN(n29901) );
  SDFFX1 \mem2_reg[230][18]  ( .D(n12254), .SI(\mem2[230][17] ), .SE(test_se), 
        .CLK(n1901), .Q(\mem2[230][18] ), .QN(n29902) );
  SDFFX1 \mem2_reg[230][17]  ( .D(n12253), .SI(\mem2[230][16] ), .SE(test_se), 
        .CLK(n1901), .Q(\mem2[230][17] ), .QN(n29903) );
  SDFFX1 \mem2_reg[230][16]  ( .D(n12252), .SI(\mem2[229][23] ), .SE(test_se), 
        .CLK(n1901), .Q(\mem2[230][16] ), .QN(n29904) );
  SDFFX1 \mem2_reg[229][23]  ( .D(n12251), .SI(\mem2[229][22] ), .SE(test_se), 
        .CLK(n1901), .Q(\mem2[229][23] ), .QN(n29905) );
  SDFFX1 \mem2_reg[229][22]  ( .D(n12250), .SI(\mem2[229][21] ), .SE(test_se), 
        .CLK(n1901), .Q(\mem2[229][22] ), .QN(n29906) );
  SDFFX1 \mem2_reg[229][21]  ( .D(n12249), .SI(\mem2[229][20] ), .SE(test_se), 
        .CLK(n1902), .Q(\mem2[229][21] ), .QN(n29907) );
  SDFFX1 \mem2_reg[229][20]  ( .D(n12248), .SI(\mem2[229][19] ), .SE(test_se), 
        .CLK(n1902), .Q(\mem2[229][20] ), .QN(n29908) );
  SDFFX1 \mem2_reg[229][19]  ( .D(n12247), .SI(\mem2[229][18] ), .SE(test_se), 
        .CLK(n1902), .Q(\mem2[229][19] ), .QN(n29909) );
  SDFFX1 \mem2_reg[229][18]  ( .D(n12246), .SI(\mem2[229][17] ), .SE(test_se), 
        .CLK(n1902), .Q(\mem2[229][18] ), .QN(n29910) );
  SDFFX1 \mem2_reg[229][17]  ( .D(n12245), .SI(\mem2[229][16] ), .SE(test_se), 
        .CLK(n1902), .Q(\mem2[229][17] ), .QN(n29911) );
  SDFFX1 \mem2_reg[229][16]  ( .D(n12244), .SI(\mem2[228][23] ), .SE(test_se), 
        .CLK(n1902), .Q(\mem2[229][16] ), .QN(n29912) );
  SDFFX1 \mem2_reg[228][23]  ( .D(n12243), .SI(\mem2[228][22] ), .SE(test_se), 
        .CLK(n1902), .Q(\mem2[228][23] ), .QN(n29913) );
  SDFFX1 \mem2_reg[228][22]  ( .D(n12242), .SI(\mem2[228][21] ), .SE(test_se), 
        .CLK(n1902), .Q(\mem2[228][22] ), .QN(n29914) );
  SDFFX1 \mem2_reg[228][21]  ( .D(n12241), .SI(\mem2[228][20] ), .SE(test_se), 
        .CLK(n1902), .Q(\mem2[228][21] ), .QN(n29915) );
  SDFFX1 \mem2_reg[228][20]  ( .D(n12240), .SI(\mem2[228][19] ), .SE(test_se), 
        .CLK(n1902), .Q(\mem2[228][20] ), .QN(n29916) );
  SDFFX1 \mem2_reg[228][19]  ( .D(n12239), .SI(\mem2[228][18] ), .SE(test_se), 
        .CLK(n1902), .Q(\mem2[228][19] ), .QN(n29917) );
  SDFFX1 \mem2_reg[228][18]  ( .D(n12238), .SI(\mem2[228][17] ), .SE(test_se), 
        .CLK(n1902), .Q(\mem2[228][18] ), .QN(n29918) );
  SDFFX1 \mem2_reg[228][17]  ( .D(n12237), .SI(\mem2[228][16] ), .SE(test_se), 
        .CLK(n1903), .Q(\mem2[228][17] ), .QN(n29919) );
  SDFFX1 \mem2_reg[228][16]  ( .D(n12236), .SI(\mem2[227][23] ), .SE(test_se), 
        .CLK(n1903), .Q(\mem2[228][16] ), .QN(n29920) );
  SDFFX1 \mem2_reg[227][23]  ( .D(n12235), .SI(\mem2[227][22] ), .SE(test_se), 
        .CLK(n1903), .Q(\mem2[227][23] ), .QN(n29921) );
  SDFFX1 \mem2_reg[227][22]  ( .D(n12234), .SI(\mem2[227][21] ), .SE(test_se), 
        .CLK(n1903), .Q(\mem2[227][22] ), .QN(n29922) );
  SDFFX1 \mem2_reg[227][21]  ( .D(n12233), .SI(\mem2[227][20] ), .SE(test_se), 
        .CLK(n1903), .Q(\mem2[227][21] ), .QN(n29923) );
  SDFFX1 \mem2_reg[227][20]  ( .D(n12232), .SI(\mem2[227][19] ), .SE(test_se), 
        .CLK(n1903), .Q(\mem2[227][20] ), .QN(n29924) );
  SDFFX1 \mem2_reg[227][19]  ( .D(n12231), .SI(\mem2[227][18] ), .SE(test_se), 
        .CLK(n1903), .Q(\mem2[227][19] ), .QN(n29925) );
  SDFFX1 \mem2_reg[227][18]  ( .D(n12230), .SI(\mem2[227][17] ), .SE(test_se), 
        .CLK(n1903), .Q(\mem2[227][18] ), .QN(n29926) );
  SDFFX1 \mem2_reg[227][17]  ( .D(n12229), .SI(\mem2[227][16] ), .SE(test_se), 
        .CLK(n1903), .Q(\mem2[227][17] ), .QN(n29927) );
  SDFFX1 \mem2_reg[227][16]  ( .D(n12228), .SI(\mem2[226][23] ), .SE(test_se), 
        .CLK(n1903), .Q(\mem2[227][16] ), .QN(n29928) );
  SDFFX1 \mem2_reg[226][23]  ( .D(n12227), .SI(\mem2[226][22] ), .SE(test_se), 
        .CLK(n1903), .Q(\mem2[226][23] ), .QN(n29929) );
  SDFFX1 \mem2_reg[226][22]  ( .D(n12226), .SI(\mem2[226][21] ), .SE(test_se), 
        .CLK(n1903), .Q(\mem2[226][22] ), .QN(n29930) );
  SDFFX1 \mem2_reg[226][21]  ( .D(n12225), .SI(\mem2[226][20] ), .SE(test_se), 
        .CLK(n1904), .Q(\mem2[226][21] ), .QN(n29931) );
  SDFFX1 \mem2_reg[226][20]  ( .D(n12224), .SI(\mem2[226][19] ), .SE(test_se), 
        .CLK(n1904), .Q(\mem2[226][20] ), .QN(n29932) );
  SDFFX1 \mem2_reg[226][19]  ( .D(n12223), .SI(\mem2[226][18] ), .SE(test_se), 
        .CLK(n1904), .Q(\mem2[226][19] ), .QN(n29933) );
  SDFFX1 \mem2_reg[226][18]  ( .D(n12222), .SI(\mem2[226][17] ), .SE(test_se), 
        .CLK(n1904), .Q(\mem2[226][18] ), .QN(n29934) );
  SDFFX1 \mem2_reg[226][17]  ( .D(n12221), .SI(\mem2[226][16] ), .SE(test_se), 
        .CLK(n1904), .Q(\mem2[226][17] ), .QN(n29935) );
  SDFFX1 \mem2_reg[226][16]  ( .D(n12220), .SI(\mem2[225][23] ), .SE(test_se), 
        .CLK(n1904), .Q(\mem2[226][16] ), .QN(n29936) );
  SDFFX1 \mem2_reg[225][23]  ( .D(n12219), .SI(\mem2[225][22] ), .SE(test_se), 
        .CLK(n1904), .Q(\mem2[225][23] ), .QN(n29937) );
  SDFFX1 \mem2_reg[225][22]  ( .D(n12218), .SI(\mem2[225][21] ), .SE(test_se), 
        .CLK(n1904), .Q(\mem2[225][22] ), .QN(n29938) );
  SDFFX1 \mem2_reg[225][21]  ( .D(n12217), .SI(\mem2[225][20] ), .SE(test_se), 
        .CLK(n1904), .Q(\mem2[225][21] ), .QN(n29939) );
  SDFFX1 \mem2_reg[225][20]  ( .D(n12216), .SI(\mem2[225][19] ), .SE(test_se), 
        .CLK(n1904), .Q(\mem2[225][20] ), .QN(n29940) );
  SDFFX1 \mem2_reg[225][19]  ( .D(n12215), .SI(\mem2[225][18] ), .SE(test_se), 
        .CLK(n1904), .Q(\mem2[225][19] ), .QN(n29941) );
  SDFFX1 \mem2_reg[225][18]  ( .D(n12214), .SI(\mem2[225][17] ), .SE(test_se), 
        .CLK(n1904), .Q(\mem2[225][18] ), .QN(n29942) );
  SDFFX1 \mem2_reg[225][17]  ( .D(n12213), .SI(\mem2[225][16] ), .SE(test_se), 
        .CLK(n1905), .Q(\mem2[225][17] ), .QN(n29943) );
  SDFFX1 \mem2_reg[225][16]  ( .D(n12212), .SI(\mem2[224][23] ), .SE(test_se), 
        .CLK(n1905), .Q(\mem2[225][16] ), .QN(n29944) );
  SDFFX1 \mem2_reg[224][23]  ( .D(n12211), .SI(\mem2[224][22] ), .SE(test_se), 
        .CLK(n1905), .Q(\mem2[224][23] ), .QN(n29945) );
  SDFFX1 \mem2_reg[224][22]  ( .D(n12210), .SI(\mem2[224][21] ), .SE(test_se), 
        .CLK(n1905), .Q(\mem2[224][22] ), .QN(n29946) );
  SDFFX1 \mem2_reg[224][21]  ( .D(n12209), .SI(\mem2[224][20] ), .SE(test_se), 
        .CLK(n1905), .Q(\mem2[224][21] ), .QN(n29947) );
  SDFFX1 \mem2_reg[224][20]  ( .D(n12208), .SI(\mem2[224][19] ), .SE(test_se), 
        .CLK(n1905), .Q(\mem2[224][20] ), .QN(n29948) );
  SDFFX1 \mem2_reg[224][19]  ( .D(n12207), .SI(\mem2[224][18] ), .SE(test_se), 
        .CLK(n1905), .Q(\mem2[224][19] ), .QN(n29949) );
  SDFFX1 \mem2_reg[224][18]  ( .D(n12206), .SI(\mem2[224][17] ), .SE(test_se), 
        .CLK(n1905), .Q(\mem2[224][18] ), .QN(n29950) );
  SDFFX1 \mem2_reg[224][17]  ( .D(n12205), .SI(\mem2[224][16] ), .SE(test_se), 
        .CLK(n1905), .Q(\mem2[224][17] ), .QN(n29951) );
  SDFFX1 \mem2_reg[224][16]  ( .D(n12204), .SI(\mem2[223][23] ), .SE(test_se), 
        .CLK(n1905), .Q(\mem2[224][16] ), .QN(n29952) );
  SDFFX1 \mem2_reg[223][23]  ( .D(n12203), .SI(\mem2[223][22] ), .SE(test_se), 
        .CLK(n1905), .Q(\mem2[223][23] ), .QN(n29953) );
  SDFFX1 \mem2_reg[223][22]  ( .D(n12202), .SI(\mem2[223][21] ), .SE(test_se), 
        .CLK(n1905), .Q(\mem2[223][22] ), .QN(n29954) );
  SDFFX1 \mem2_reg[223][21]  ( .D(n12201), .SI(\mem2[223][20] ), .SE(test_se), 
        .CLK(n1906), .Q(\mem2[223][21] ), .QN(n29955) );
  SDFFX1 \mem2_reg[223][20]  ( .D(n12200), .SI(\mem2[223][19] ), .SE(test_se), 
        .CLK(n1906), .Q(\mem2[223][20] ), .QN(n29956) );
  SDFFX1 \mem2_reg[223][19]  ( .D(n12199), .SI(\mem2[223][18] ), .SE(test_se), 
        .CLK(n1906), .Q(\mem2[223][19] ), .QN(n29957) );
  SDFFX1 \mem2_reg[223][18]  ( .D(n12198), .SI(\mem2[223][17] ), .SE(test_se), 
        .CLK(n1906), .Q(\mem2[223][18] ), .QN(n29958) );
  SDFFX1 \mem2_reg[223][17]  ( .D(n12197), .SI(\mem2[223][16] ), .SE(test_se), 
        .CLK(n1906), .Q(\mem2[223][17] ), .QN(n29959) );
  SDFFX1 \mem2_reg[223][16]  ( .D(n12196), .SI(\mem2[222][23] ), .SE(test_se), 
        .CLK(n1906), .Q(\mem2[223][16] ), .QN(n29960) );
  SDFFX1 \mem2_reg[222][23]  ( .D(n12195), .SI(\mem2[222][22] ), .SE(test_se), 
        .CLK(n1906), .Q(\mem2[222][23] ), .QN(n29961) );
  SDFFX1 \mem2_reg[222][22]  ( .D(n12194), .SI(\mem2[222][21] ), .SE(test_se), 
        .CLK(n1906), .Q(\mem2[222][22] ), .QN(n29962) );
  SDFFX1 \mem2_reg[222][21]  ( .D(n12193), .SI(\mem2[222][20] ), .SE(test_se), 
        .CLK(n1906), .Q(\mem2[222][21] ), .QN(n29963) );
  SDFFX1 \mem2_reg[222][20]  ( .D(n12192), .SI(\mem2[222][19] ), .SE(test_se), 
        .CLK(n1906), .Q(\mem2[222][20] ), .QN(n29964) );
  SDFFX1 \mem2_reg[222][19]  ( .D(n12191), .SI(\mem2[222][18] ), .SE(test_se), 
        .CLK(n1906), .Q(\mem2[222][19] ), .QN(n29965) );
  SDFFX1 \mem2_reg[222][18]  ( .D(n12190), .SI(\mem2[222][17] ), .SE(test_se), 
        .CLK(n1906), .Q(\mem2[222][18] ), .QN(n29966) );
  SDFFX1 \mem2_reg[222][17]  ( .D(n12189), .SI(\mem2[222][16] ), .SE(test_se), 
        .CLK(n1907), .Q(\mem2[222][17] ), .QN(n29967) );
  SDFFX1 \mem2_reg[222][16]  ( .D(n12188), .SI(\mem2[221][23] ), .SE(test_se), 
        .CLK(n1907), .Q(\mem2[222][16] ), .QN(n29968) );
  SDFFX1 \mem2_reg[221][23]  ( .D(n12187), .SI(\mem2[221][22] ), .SE(test_se), 
        .CLK(n1907), .Q(\mem2[221][23] ), .QN(n29969) );
  SDFFX1 \mem2_reg[221][22]  ( .D(n12186), .SI(\mem2[221][21] ), .SE(test_se), 
        .CLK(n1907), .Q(\mem2[221][22] ), .QN(n29970) );
  SDFFX1 \mem2_reg[221][21]  ( .D(n12185), .SI(\mem2[221][20] ), .SE(test_se), 
        .CLK(n1907), .Q(\mem2[221][21] ), .QN(n29971) );
  SDFFX1 \mem2_reg[221][20]  ( .D(n12184), .SI(\mem2[221][19] ), .SE(test_se), 
        .CLK(n1907), .Q(\mem2[221][20] ), .QN(n29972) );
  SDFFX1 \mem2_reg[221][19]  ( .D(n12183), .SI(\mem2[221][18] ), .SE(test_se), 
        .CLK(n1907), .Q(\mem2[221][19] ), .QN(n29973) );
  SDFFX1 \mem2_reg[221][18]  ( .D(n12182), .SI(\mem2[221][17] ), .SE(test_se), 
        .CLK(n1907), .Q(\mem2[221][18] ), .QN(n29974) );
  SDFFX1 \mem2_reg[221][17]  ( .D(n12181), .SI(\mem2[221][16] ), .SE(test_se), 
        .CLK(n1907), .Q(\mem2[221][17] ), .QN(n29975) );
  SDFFX1 \mem2_reg[221][16]  ( .D(n12180), .SI(\mem2[220][23] ), .SE(test_se), 
        .CLK(n1907), .Q(\mem2[221][16] ), .QN(n29976) );
  SDFFX1 \mem2_reg[220][23]  ( .D(n12179), .SI(\mem2[220][22] ), .SE(test_se), 
        .CLK(n1907), .Q(\mem2[220][23] ), .QN(n29977) );
  SDFFX1 \mem2_reg[220][22]  ( .D(n12178), .SI(\mem2[220][21] ), .SE(test_se), 
        .CLK(n1907), .Q(\mem2[220][22] ), .QN(n29978) );
  SDFFX1 \mem2_reg[220][21]  ( .D(n12177), .SI(\mem2[220][20] ), .SE(test_se), 
        .CLK(n1908), .Q(\mem2[220][21] ), .QN(n29979) );
  SDFFX1 \mem2_reg[220][20]  ( .D(n12176), .SI(\mem2[220][19] ), .SE(test_se), 
        .CLK(n1908), .Q(\mem2[220][20] ), .QN(n29980) );
  SDFFX1 \mem2_reg[220][19]  ( .D(n12175), .SI(\mem2[220][18] ), .SE(test_se), 
        .CLK(n1908), .Q(\mem2[220][19] ), .QN(n29981) );
  SDFFX1 \mem2_reg[220][18]  ( .D(n12174), .SI(\mem2[220][17] ), .SE(test_se), 
        .CLK(n1908), .Q(\mem2[220][18] ), .QN(n29982) );
  SDFFX1 \mem2_reg[220][17]  ( .D(n12173), .SI(\mem2[220][16] ), .SE(test_se), 
        .CLK(n1908), .Q(\mem2[220][17] ), .QN(n29983) );
  SDFFX1 \mem2_reg[220][16]  ( .D(n12172), .SI(\mem2[219][23] ), .SE(test_se), 
        .CLK(n1908), .Q(\mem2[220][16] ), .QN(n29984) );
  SDFFX1 \mem2_reg[219][23]  ( .D(n12171), .SI(\mem2[219][22] ), .SE(test_se), 
        .CLK(n1908), .Q(\mem2[219][23] ), .QN(n29985) );
  SDFFX1 \mem2_reg[219][22]  ( .D(n12170), .SI(\mem2[219][21] ), .SE(test_se), 
        .CLK(n1908), .Q(\mem2[219][22] ), .QN(n29986) );
  SDFFX1 \mem2_reg[219][21]  ( .D(n12169), .SI(\mem2[219][20] ), .SE(test_se), 
        .CLK(n1908), .Q(\mem2[219][21] ), .QN(n29987) );
  SDFFX1 \mem2_reg[219][20]  ( .D(n12168), .SI(\mem2[219][19] ), .SE(test_se), 
        .CLK(n1908), .Q(\mem2[219][20] ), .QN(n29988) );
  SDFFX1 \mem2_reg[219][19]  ( .D(n12167), .SI(\mem2[219][18] ), .SE(test_se), 
        .CLK(n1908), .Q(\mem2[219][19] ), .QN(n29989) );
  SDFFX1 \mem2_reg[219][18]  ( .D(n12166), .SI(\mem2[219][17] ), .SE(test_se), 
        .CLK(n1908), .Q(\mem2[219][18] ), .QN(n29990) );
  SDFFX1 \mem2_reg[219][17]  ( .D(n12165), .SI(\mem2[219][16] ), .SE(test_se), 
        .CLK(n1909), .Q(\mem2[219][17] ), .QN(n29991) );
  SDFFX1 \mem2_reg[219][16]  ( .D(n12164), .SI(\mem2[218][23] ), .SE(test_se), 
        .CLK(n1909), .Q(\mem2[219][16] ), .QN(n29992) );
  SDFFX1 \mem2_reg[218][23]  ( .D(n12163), .SI(\mem2[218][22] ), .SE(test_se), 
        .CLK(n1909), .Q(\mem2[218][23] ), .QN(n29993) );
  SDFFX1 \mem2_reg[218][22]  ( .D(n12162), .SI(\mem2[218][21] ), .SE(test_se), 
        .CLK(n1909), .Q(\mem2[218][22] ), .QN(n29994) );
  SDFFX1 \mem2_reg[218][21]  ( .D(n12161), .SI(\mem2[218][20] ), .SE(test_se), 
        .CLK(n1909), .Q(\mem2[218][21] ), .QN(n29995) );
  SDFFX1 \mem2_reg[218][20]  ( .D(n12160), .SI(\mem2[218][19] ), .SE(test_se), 
        .CLK(n1909), .Q(\mem2[218][20] ), .QN(n29996) );
  SDFFX1 \mem2_reg[218][19]  ( .D(n12159), .SI(\mem2[218][18] ), .SE(test_se), 
        .CLK(n1909), .Q(\mem2[218][19] ), .QN(n29997) );
  SDFFX1 \mem2_reg[218][18]  ( .D(n12158), .SI(\mem2[218][17] ), .SE(test_se), 
        .CLK(n1909), .Q(\mem2[218][18] ), .QN(n29998) );
  SDFFX1 \mem2_reg[218][17]  ( .D(n12157), .SI(\mem2[218][16] ), .SE(test_se), 
        .CLK(n1909), .Q(\mem2[218][17] ), .QN(n29999) );
  SDFFX1 \mem2_reg[218][16]  ( .D(n12156), .SI(\mem2[217][23] ), .SE(test_se), 
        .CLK(n1909), .Q(\mem2[218][16] ), .QN(n30000) );
  SDFFX1 \mem2_reg[217][23]  ( .D(n12155), .SI(\mem2[217][22] ), .SE(test_se), 
        .CLK(n1909), .Q(\mem2[217][23] ), .QN(n30001) );
  SDFFX1 \mem2_reg[217][22]  ( .D(n12154), .SI(\mem2[217][21] ), .SE(test_se), 
        .CLK(n1909), .Q(\mem2[217][22] ), .QN(n30002) );
  SDFFX1 \mem2_reg[217][21]  ( .D(n12153), .SI(\mem2[217][20] ), .SE(test_se), 
        .CLK(n1910), .Q(\mem2[217][21] ), .QN(n30003) );
  SDFFX1 \mem2_reg[217][20]  ( .D(n12152), .SI(\mem2[217][19] ), .SE(test_se), 
        .CLK(n1910), .Q(\mem2[217][20] ), .QN(n30004) );
  SDFFX1 \mem2_reg[217][19]  ( .D(n12151), .SI(\mem2[217][18] ), .SE(test_se), 
        .CLK(n1910), .Q(\mem2[217][19] ), .QN(n30005) );
  SDFFX1 \mem2_reg[217][18]  ( .D(n12150), .SI(\mem2[217][17] ), .SE(test_se), 
        .CLK(n1910), .Q(\mem2[217][18] ), .QN(n30006) );
  SDFFX1 \mem2_reg[217][17]  ( .D(n12149), .SI(\mem2[217][16] ), .SE(test_se), 
        .CLK(n1910), .Q(\mem2[217][17] ), .QN(n30007) );
  SDFFX1 \mem2_reg[217][16]  ( .D(n12148), .SI(\mem2[216][23] ), .SE(test_se), 
        .CLK(n1910), .Q(\mem2[217][16] ), .QN(n30008) );
  SDFFX1 \mem2_reg[216][23]  ( .D(n12147), .SI(\mem2[216][22] ), .SE(test_se), 
        .CLK(n1910), .Q(\mem2[216][23] ), .QN(n30009) );
  SDFFX1 \mem2_reg[216][22]  ( .D(n12146), .SI(\mem2[216][21] ), .SE(test_se), 
        .CLK(n1910), .Q(\mem2[216][22] ), .QN(n30010) );
  SDFFX1 \mem2_reg[216][21]  ( .D(n12145), .SI(\mem2[216][20] ), .SE(test_se), 
        .CLK(n1910), .Q(\mem2[216][21] ), .QN(n30011) );
  SDFFX1 \mem2_reg[216][20]  ( .D(n12144), .SI(\mem2[216][19] ), .SE(test_se), 
        .CLK(n1910), .Q(\mem2[216][20] ), .QN(n30012) );
  SDFFX1 \mem2_reg[216][19]  ( .D(n12143), .SI(\mem2[216][18] ), .SE(test_se), 
        .CLK(n1910), .Q(\mem2[216][19] ), .QN(n30013) );
  SDFFX1 \mem2_reg[216][18]  ( .D(n12142), .SI(\mem2[216][17] ), .SE(test_se), 
        .CLK(n1910), .Q(\mem2[216][18] ), .QN(n30014) );
  SDFFX1 \mem2_reg[216][17]  ( .D(n12141), .SI(\mem2[216][16] ), .SE(test_se), 
        .CLK(n1911), .Q(\mem2[216][17] ), .QN(n30015) );
  SDFFX1 \mem2_reg[216][16]  ( .D(n12140), .SI(\mem2[215][23] ), .SE(test_se), 
        .CLK(n1911), .Q(\mem2[216][16] ), .QN(n30016) );
  SDFFX1 \mem2_reg[215][23]  ( .D(n12139), .SI(\mem2[215][22] ), .SE(test_se), 
        .CLK(n1911), .Q(\mem2[215][23] ), .QN(n30017) );
  SDFFX1 \mem2_reg[215][22]  ( .D(n12138), .SI(\mem2[215][21] ), .SE(test_se), 
        .CLK(n1911), .Q(\mem2[215][22] ), .QN(n30018) );
  SDFFX1 \mem2_reg[215][21]  ( .D(n12137), .SI(\mem2[215][20] ), .SE(test_se), 
        .CLK(n1911), .Q(\mem2[215][21] ), .QN(n30019) );
  SDFFX1 \mem2_reg[215][20]  ( .D(n12136), .SI(\mem2[215][19] ), .SE(test_se), 
        .CLK(n1911), .Q(\mem2[215][20] ), .QN(n30020) );
  SDFFX1 \mem2_reg[215][19]  ( .D(n12135), .SI(\mem2[215][18] ), .SE(test_se), 
        .CLK(n1911), .Q(\mem2[215][19] ), .QN(n30021) );
  SDFFX1 \mem2_reg[215][18]  ( .D(n12134), .SI(\mem2[215][17] ), .SE(test_se), 
        .CLK(n1911), .Q(\mem2[215][18] ), .QN(n30022) );
  SDFFX1 \mem2_reg[215][17]  ( .D(n12133), .SI(\mem2[215][16] ), .SE(test_se), 
        .CLK(n1911), .Q(\mem2[215][17] ), .QN(n30023) );
  SDFFX1 \mem2_reg[215][16]  ( .D(n12132), .SI(\mem2[214][23] ), .SE(test_se), 
        .CLK(n1911), .Q(\mem2[215][16] ), .QN(n30024) );
  SDFFX1 \mem2_reg[214][23]  ( .D(n12131), .SI(\mem2[214][22] ), .SE(test_se), 
        .CLK(n1911), .Q(\mem2[214][23] ), .QN(n30025) );
  SDFFX1 \mem2_reg[214][22]  ( .D(n12130), .SI(\mem2[214][21] ), .SE(test_se), 
        .CLK(n1911), .Q(\mem2[214][22] ), .QN(n30026) );
  SDFFX1 \mem2_reg[214][21]  ( .D(n12129), .SI(\mem2[214][20] ), .SE(test_se), 
        .CLK(n1912), .Q(\mem2[214][21] ), .QN(n30027) );
  SDFFX1 \mem2_reg[214][20]  ( .D(n12128), .SI(\mem2[214][19] ), .SE(test_se), 
        .CLK(n1912), .Q(\mem2[214][20] ), .QN(n30028) );
  SDFFX1 \mem2_reg[214][19]  ( .D(n12127), .SI(\mem2[214][18] ), .SE(test_se), 
        .CLK(n1912), .Q(\mem2[214][19] ), .QN(n30029) );
  SDFFX1 \mem2_reg[214][18]  ( .D(n12126), .SI(\mem2[214][17] ), .SE(test_se), 
        .CLK(n1912), .Q(\mem2[214][18] ), .QN(n30030) );
  SDFFX1 \mem2_reg[214][17]  ( .D(n12125), .SI(\mem2[214][16] ), .SE(test_se), 
        .CLK(n1912), .Q(\mem2[214][17] ), .QN(n30031) );
  SDFFX1 \mem2_reg[214][16]  ( .D(n12124), .SI(\mem2[213][23] ), .SE(test_se), 
        .CLK(n1912), .Q(\mem2[214][16] ), .QN(n30032) );
  SDFFX1 \mem2_reg[213][23]  ( .D(n12123), .SI(\mem2[213][22] ), .SE(test_se), 
        .CLK(n1912), .Q(\mem2[213][23] ), .QN(n30033) );
  SDFFX1 \mem2_reg[213][22]  ( .D(n12122), .SI(\mem2[213][21] ), .SE(test_se), 
        .CLK(n1912), .Q(\mem2[213][22] ), .QN(n30034) );
  SDFFX1 \mem2_reg[213][21]  ( .D(n12121), .SI(\mem2[213][20] ), .SE(test_se), 
        .CLK(n1912), .Q(\mem2[213][21] ), .QN(n30035) );
  SDFFX1 \mem2_reg[213][20]  ( .D(n12120), .SI(\mem2[213][19] ), .SE(test_se), 
        .CLK(n1912), .Q(\mem2[213][20] ), .QN(n30036) );
  SDFFX1 \mem2_reg[213][19]  ( .D(n12119), .SI(\mem2[213][18] ), .SE(test_se), 
        .CLK(n1912), .Q(\mem2[213][19] ), .QN(n30037) );
  SDFFX1 \mem2_reg[213][18]  ( .D(n12118), .SI(\mem2[213][17] ), .SE(test_se), 
        .CLK(n1912), .Q(\mem2[213][18] ), .QN(n30038) );
  SDFFX1 \mem2_reg[213][17]  ( .D(n12117), .SI(\mem2[213][16] ), .SE(test_se), 
        .CLK(n1913), .Q(\mem2[213][17] ), .QN(n30039) );
  SDFFX1 \mem2_reg[213][16]  ( .D(n12116), .SI(\mem2[212][23] ), .SE(test_se), 
        .CLK(n1913), .Q(\mem2[213][16] ), .QN(n30040) );
  SDFFX1 \mem2_reg[212][23]  ( .D(n12115), .SI(\mem2[212][22] ), .SE(test_se), 
        .CLK(n1913), .Q(\mem2[212][23] ), .QN(n30041) );
  SDFFX1 \mem2_reg[212][22]  ( .D(n12114), .SI(\mem2[212][21] ), .SE(test_se), 
        .CLK(n1913), .Q(\mem2[212][22] ), .QN(n30042) );
  SDFFX1 \mem2_reg[212][21]  ( .D(n12113), .SI(\mem2[212][20] ), .SE(test_se), 
        .CLK(n1913), .Q(\mem2[212][21] ), .QN(n30043) );
  SDFFX1 \mem2_reg[212][20]  ( .D(n12112), .SI(\mem2[212][19] ), .SE(test_se), 
        .CLK(n1913), .Q(\mem2[212][20] ), .QN(n30044) );
  SDFFX1 \mem2_reg[212][19]  ( .D(n12111), .SI(\mem2[212][18] ), .SE(test_se), 
        .CLK(n1913), .Q(\mem2[212][19] ), .QN(n30045) );
  SDFFX1 \mem2_reg[212][18]  ( .D(n12110), .SI(\mem2[212][17] ), .SE(test_se), 
        .CLK(n1913), .Q(\mem2[212][18] ), .QN(n30046) );
  SDFFX1 \mem2_reg[212][17]  ( .D(n12109), .SI(\mem2[212][16] ), .SE(test_se), 
        .CLK(n1913), .Q(\mem2[212][17] ), .QN(n30047) );
  SDFFX1 \mem2_reg[212][16]  ( .D(n12108), .SI(\mem2[211][23] ), .SE(test_se), 
        .CLK(n1913), .Q(\mem2[212][16] ), .QN(n30048) );
  SDFFX1 \mem2_reg[211][23]  ( .D(n12107), .SI(\mem2[211][22] ), .SE(test_se), 
        .CLK(n1913), .Q(\mem2[211][23] ), .QN(n30049) );
  SDFFX1 \mem2_reg[211][22]  ( .D(n12106), .SI(\mem2[211][21] ), .SE(test_se), 
        .CLK(n1913), .Q(\mem2[211][22] ), .QN(n30050) );
  SDFFX1 \mem2_reg[211][21]  ( .D(n12105), .SI(\mem2[211][20] ), .SE(test_se), 
        .CLK(n1914), .Q(\mem2[211][21] ), .QN(n30051) );
  SDFFX1 \mem2_reg[211][20]  ( .D(n12104), .SI(\mem2[211][19] ), .SE(test_se), 
        .CLK(n1914), .Q(\mem2[211][20] ), .QN(n30052) );
  SDFFX1 \mem2_reg[211][19]  ( .D(n12103), .SI(\mem2[211][18] ), .SE(test_se), 
        .CLK(n1914), .Q(\mem2[211][19] ), .QN(n30053) );
  SDFFX1 \mem2_reg[211][18]  ( .D(n12102), .SI(\mem2[211][17] ), .SE(test_se), 
        .CLK(n1914), .Q(\mem2[211][18] ), .QN(n30054) );
  SDFFX1 \mem2_reg[211][17]  ( .D(n12101), .SI(\mem2[211][16] ), .SE(test_se), 
        .CLK(n1914), .Q(\mem2[211][17] ), .QN(n30055) );
  SDFFX1 \mem2_reg[211][16]  ( .D(n12100), .SI(\mem2[210][23] ), .SE(test_se), 
        .CLK(n1914), .Q(\mem2[211][16] ), .QN(n30056) );
  SDFFX1 \mem2_reg[210][23]  ( .D(n12099), .SI(\mem2[210][22] ), .SE(test_se), 
        .CLK(n1914), .Q(\mem2[210][23] ), .QN(n30057) );
  SDFFX1 \mem2_reg[210][22]  ( .D(n12098), .SI(\mem2[210][21] ), .SE(test_se), 
        .CLK(n1914), .Q(\mem2[210][22] ), .QN(n30058) );
  SDFFX1 \mem2_reg[210][21]  ( .D(n12097), .SI(\mem2[210][20] ), .SE(test_se), 
        .CLK(n1914), .Q(\mem2[210][21] ), .QN(n30059) );
  SDFFX1 \mem2_reg[210][20]  ( .D(n12096), .SI(\mem2[210][19] ), .SE(test_se), 
        .CLK(n1914), .Q(\mem2[210][20] ), .QN(n30060) );
  SDFFX1 \mem2_reg[210][19]  ( .D(n12095), .SI(\mem2[210][18] ), .SE(test_se), 
        .CLK(n1914), .Q(\mem2[210][19] ), .QN(n30061) );
  SDFFX1 \mem2_reg[210][18]  ( .D(n12094), .SI(\mem2[210][17] ), .SE(test_se), 
        .CLK(n1914), .Q(\mem2[210][18] ), .QN(n30062) );
  SDFFX1 \mem2_reg[210][17]  ( .D(n12093), .SI(\mem2[210][16] ), .SE(test_se), 
        .CLK(n1915), .Q(\mem2[210][17] ), .QN(n30063) );
  SDFFX1 \mem2_reg[210][16]  ( .D(n12092), .SI(\mem2[209][23] ), .SE(test_se), 
        .CLK(n1915), .Q(\mem2[210][16] ), .QN(n30064) );
  SDFFX1 \mem2_reg[209][23]  ( .D(n12091), .SI(\mem2[209][22] ), .SE(test_se), 
        .CLK(n1915), .Q(\mem2[209][23] ), .QN(n30065) );
  SDFFX1 \mem2_reg[209][22]  ( .D(n12090), .SI(\mem2[209][21] ), .SE(test_se), 
        .CLK(n1915), .Q(\mem2[209][22] ), .QN(n30066) );
  SDFFX1 \mem2_reg[209][21]  ( .D(n12089), .SI(\mem2[209][20] ), .SE(test_se), 
        .CLK(n1915), .Q(\mem2[209][21] ), .QN(n30067) );
  SDFFX1 \mem2_reg[209][20]  ( .D(n12088), .SI(\mem2[209][19] ), .SE(test_se), 
        .CLK(n1915), .Q(\mem2[209][20] ), .QN(n30068) );
  SDFFX1 \mem2_reg[209][19]  ( .D(n12087), .SI(\mem2[209][18] ), .SE(test_se), 
        .CLK(n1915), .Q(\mem2[209][19] ), .QN(n30069) );
  SDFFX1 \mem2_reg[209][18]  ( .D(n12086), .SI(\mem2[209][17] ), .SE(test_se), 
        .CLK(n1915), .Q(\mem2[209][18] ), .QN(n30070) );
  SDFFX1 \mem2_reg[209][17]  ( .D(n12085), .SI(\mem2[209][16] ), .SE(test_se), 
        .CLK(n1915), .Q(\mem2[209][17] ), .QN(n30071) );
  SDFFX1 \mem2_reg[209][16]  ( .D(n12084), .SI(\mem2[208][23] ), .SE(test_se), 
        .CLK(n1915), .Q(\mem2[209][16] ), .QN(n30072) );
  SDFFX1 \mem2_reg[208][23]  ( .D(n12083), .SI(\mem2[208][22] ), .SE(test_se), 
        .CLK(n1915), .Q(\mem2[208][23] ), .QN(n30073) );
  SDFFX1 \mem2_reg[208][22]  ( .D(n12082), .SI(\mem2[208][21] ), .SE(test_se), 
        .CLK(n1915), .Q(\mem2[208][22] ), .QN(n30074) );
  SDFFX1 \mem2_reg[208][21]  ( .D(n12081), .SI(\mem2[208][20] ), .SE(test_se), 
        .CLK(n1916), .Q(\mem2[208][21] ), .QN(n30075) );
  SDFFX1 \mem2_reg[208][20]  ( .D(n12080), .SI(\mem2[208][19] ), .SE(test_se), 
        .CLK(n1916), .Q(\mem2[208][20] ), .QN(n30076) );
  SDFFX1 \mem2_reg[208][19]  ( .D(n12079), .SI(\mem2[208][18] ), .SE(test_se), 
        .CLK(n1916), .Q(\mem2[208][19] ), .QN(n30077) );
  SDFFX1 \mem2_reg[208][18]  ( .D(n12078), .SI(\mem2[208][17] ), .SE(test_se), 
        .CLK(n1916), .Q(\mem2[208][18] ), .QN(n30078) );
  SDFFX1 \mem2_reg[208][17]  ( .D(n12077), .SI(\mem2[208][16] ), .SE(test_se), 
        .CLK(n1916), .Q(\mem2[208][17] ), .QN(n30079) );
  SDFFX1 \mem2_reg[208][16]  ( .D(n12076), .SI(\mem2[207][23] ), .SE(test_se), 
        .CLK(n1916), .Q(\mem2[208][16] ), .QN(n30080) );
  SDFFX1 \mem2_reg[207][23]  ( .D(n12075), .SI(\mem2[207][22] ), .SE(test_se), 
        .CLK(n1916), .Q(\mem2[207][23] ), .QN(n30081) );
  SDFFX1 \mem2_reg[207][22]  ( .D(n12074), .SI(\mem2[207][21] ), .SE(test_se), 
        .CLK(n1916), .Q(\mem2[207][22] ), .QN(n30082) );
  SDFFX1 \mem2_reg[207][21]  ( .D(n12073), .SI(\mem2[207][20] ), .SE(test_se), 
        .CLK(n1916), .Q(\mem2[207][21] ), .QN(n30083) );
  SDFFX1 \mem2_reg[207][20]  ( .D(n12072), .SI(\mem2[207][19] ), .SE(test_se), 
        .CLK(n1916), .Q(\mem2[207][20] ), .QN(n30084) );
  SDFFX1 \mem2_reg[207][19]  ( .D(n12071), .SI(\mem2[207][18] ), .SE(test_se), 
        .CLK(n1916), .Q(\mem2[207][19] ), .QN(n30085) );
  SDFFX1 \mem2_reg[207][18]  ( .D(n12070), .SI(\mem2[207][17] ), .SE(test_se), 
        .CLK(n1916), .Q(\mem2[207][18] ), .QN(n30086) );
  SDFFX1 \mem2_reg[207][17]  ( .D(n12069), .SI(\mem2[207][16] ), .SE(test_se), 
        .CLK(n1917), .Q(\mem2[207][17] ), .QN(n30087) );
  SDFFX1 \mem2_reg[207][16]  ( .D(n12068), .SI(\mem2[206][23] ), .SE(test_se), 
        .CLK(n1917), .Q(\mem2[207][16] ), .QN(n30088) );
  SDFFX1 \mem2_reg[206][23]  ( .D(n12067), .SI(\mem2[206][22] ), .SE(test_se), 
        .CLK(n1917), .Q(\mem2[206][23] ), .QN(n30089) );
  SDFFX1 \mem2_reg[206][22]  ( .D(n12066), .SI(\mem2[206][21] ), .SE(test_se), 
        .CLK(n1917), .Q(\mem2[206][22] ), .QN(n30090) );
  SDFFX1 \mem2_reg[206][21]  ( .D(n12065), .SI(\mem2[206][20] ), .SE(test_se), 
        .CLK(n1917), .Q(\mem2[206][21] ), .QN(n30091) );
  SDFFX1 \mem2_reg[206][20]  ( .D(n12064), .SI(\mem2[206][19] ), .SE(test_se), 
        .CLK(n1917), .Q(\mem2[206][20] ), .QN(n30092) );
  SDFFX1 \mem2_reg[206][19]  ( .D(n12063), .SI(\mem2[206][18] ), .SE(test_se), 
        .CLK(n1917), .Q(\mem2[206][19] ), .QN(n30093) );
  SDFFX1 \mem2_reg[206][18]  ( .D(n12062), .SI(\mem2[206][17] ), .SE(test_se), 
        .CLK(n1917), .Q(\mem2[206][18] ), .QN(n30094) );
  SDFFX1 \mem2_reg[206][17]  ( .D(n12061), .SI(\mem2[206][16] ), .SE(test_se), 
        .CLK(n1917), .Q(\mem2[206][17] ), .QN(n30095) );
  SDFFX1 \mem2_reg[206][16]  ( .D(n12060), .SI(\mem2[205][23] ), .SE(test_se), 
        .CLK(n1917), .Q(\mem2[206][16] ), .QN(n30096) );
  SDFFX1 \mem2_reg[205][23]  ( .D(n12059), .SI(\mem2[205][22] ), .SE(test_se), 
        .CLK(n1917), .Q(\mem2[205][23] ), .QN(n30097) );
  SDFFX1 \mem2_reg[205][22]  ( .D(n12058), .SI(\mem2[205][21] ), .SE(test_se), 
        .CLK(n1917), .Q(\mem2[205][22] ), .QN(n30098) );
  SDFFX1 \mem2_reg[205][21]  ( .D(n12057), .SI(\mem2[205][20] ), .SE(test_se), 
        .CLK(n1918), .Q(\mem2[205][21] ), .QN(n30099) );
  SDFFX1 \mem2_reg[205][20]  ( .D(n12056), .SI(\mem2[205][19] ), .SE(test_se), 
        .CLK(n1918), .Q(\mem2[205][20] ), .QN(n30100) );
  SDFFX1 \mem2_reg[205][19]  ( .D(n12055), .SI(\mem2[205][18] ), .SE(test_se), 
        .CLK(n1918), .Q(\mem2[205][19] ), .QN(n30101) );
  SDFFX1 \mem2_reg[205][18]  ( .D(n12054), .SI(\mem2[205][17] ), .SE(test_se), 
        .CLK(n1918), .Q(\mem2[205][18] ), .QN(n30102) );
  SDFFX1 \mem2_reg[205][17]  ( .D(n12053), .SI(\mem2[205][16] ), .SE(test_se), 
        .CLK(n1918), .Q(\mem2[205][17] ), .QN(n30103) );
  SDFFX1 \mem2_reg[205][16]  ( .D(n12052), .SI(\mem2[204][23] ), .SE(test_se), 
        .CLK(n1918), .Q(\mem2[205][16] ), .QN(n30104) );
  SDFFX1 \mem2_reg[204][23]  ( .D(n12051), .SI(\mem2[204][22] ), .SE(test_se), 
        .CLK(n1918), .Q(\mem2[204][23] ), .QN(n30105) );
  SDFFX1 \mem2_reg[204][22]  ( .D(n12050), .SI(\mem2[204][21] ), .SE(test_se), 
        .CLK(n1918), .Q(\mem2[204][22] ), .QN(n30106) );
  SDFFX1 \mem2_reg[204][21]  ( .D(n12049), .SI(\mem2[204][20] ), .SE(test_se), 
        .CLK(n1918), .Q(\mem2[204][21] ), .QN(n30107) );
  SDFFX1 \mem2_reg[204][20]  ( .D(n12048), .SI(\mem2[204][19] ), .SE(test_se), 
        .CLK(n1918), .Q(\mem2[204][20] ), .QN(n30108) );
  SDFFX1 \mem2_reg[204][19]  ( .D(n12047), .SI(\mem2[204][18] ), .SE(test_se), 
        .CLK(n1918), .Q(\mem2[204][19] ), .QN(n30109) );
  SDFFX1 \mem2_reg[204][18]  ( .D(n12046), .SI(\mem2[204][17] ), .SE(test_se), 
        .CLK(n1918), .Q(\mem2[204][18] ), .QN(n30110) );
  SDFFX1 \mem2_reg[204][17]  ( .D(n12045), .SI(\mem2[204][16] ), .SE(test_se), 
        .CLK(n1919), .Q(\mem2[204][17] ), .QN(n30111) );
  SDFFX1 \mem2_reg[204][16]  ( .D(n12044), .SI(\mem2[203][23] ), .SE(test_se), 
        .CLK(n1919), .Q(\mem2[204][16] ), .QN(n30112) );
  SDFFX1 \mem2_reg[203][23]  ( .D(n12043), .SI(\mem2[203][22] ), .SE(test_se), 
        .CLK(n1919), .Q(\mem2[203][23] ), .QN(n30113) );
  SDFFX1 \mem2_reg[203][22]  ( .D(n12042), .SI(\mem2[203][21] ), .SE(test_se), 
        .CLK(n1919), .Q(\mem2[203][22] ), .QN(n30114) );
  SDFFX1 \mem2_reg[203][21]  ( .D(n12041), .SI(\mem2[203][20] ), .SE(test_se), 
        .CLK(n1919), .Q(\mem2[203][21] ), .QN(n30115) );
  SDFFX1 \mem2_reg[203][20]  ( .D(n12040), .SI(\mem2[203][19] ), .SE(test_se), 
        .CLK(n1919), .Q(\mem2[203][20] ), .QN(n30116) );
  SDFFX1 \mem2_reg[203][19]  ( .D(n12039), .SI(\mem2[203][18] ), .SE(test_se), 
        .CLK(n1919), .Q(\mem2[203][19] ), .QN(n30117) );
  SDFFX1 \mem2_reg[203][18]  ( .D(n12038), .SI(\mem2[203][17] ), .SE(test_se), 
        .CLK(n1919), .Q(\mem2[203][18] ), .QN(n30118) );
  SDFFX1 \mem2_reg[203][17]  ( .D(n12037), .SI(\mem2[203][16] ), .SE(test_se), 
        .CLK(n1919), .Q(\mem2[203][17] ), .QN(n30119) );
  SDFFX1 \mem2_reg[203][16]  ( .D(n12036), .SI(\mem2[202][23] ), .SE(test_se), 
        .CLK(n1919), .Q(\mem2[203][16] ), .QN(n30120) );
  SDFFX1 \mem2_reg[202][23]  ( .D(n12035), .SI(\mem2[202][22] ), .SE(test_se), 
        .CLK(n1919), .Q(\mem2[202][23] ), .QN(n30121) );
  SDFFX1 \mem2_reg[202][22]  ( .D(n12034), .SI(\mem2[202][21] ), .SE(test_se), 
        .CLK(n1919), .Q(\mem2[202][22] ), .QN(n30122) );
  SDFFX1 \mem2_reg[202][21]  ( .D(n12033), .SI(\mem2[202][20] ), .SE(test_se), 
        .CLK(n1920), .Q(\mem2[202][21] ), .QN(n30123) );
  SDFFX1 \mem2_reg[202][20]  ( .D(n12032), .SI(\mem2[202][19] ), .SE(test_se), 
        .CLK(n1920), .Q(\mem2[202][20] ), .QN(n30124) );
  SDFFX1 \mem2_reg[202][19]  ( .D(n12031), .SI(\mem2[202][18] ), .SE(test_se), 
        .CLK(n1920), .Q(\mem2[202][19] ), .QN(n30125) );
  SDFFX1 \mem2_reg[202][18]  ( .D(n12030), .SI(\mem2[202][17] ), .SE(test_se), 
        .CLK(n1920), .Q(\mem2[202][18] ), .QN(n30126) );
  SDFFX1 \mem2_reg[202][17]  ( .D(n12029), .SI(\mem2[202][16] ), .SE(test_se), 
        .CLK(n1920), .Q(\mem2[202][17] ), .QN(n30127) );
  SDFFX1 \mem2_reg[202][16]  ( .D(n12028), .SI(\mem2[201][23] ), .SE(test_se), 
        .CLK(n1920), .Q(\mem2[202][16] ), .QN(n30128) );
  SDFFX1 \mem2_reg[201][23]  ( .D(n12027), .SI(\mem2[201][22] ), .SE(test_se), 
        .CLK(n1920), .Q(\mem2[201][23] ), .QN(n30129) );
  SDFFX1 \mem2_reg[201][22]  ( .D(n12026), .SI(\mem2[201][21] ), .SE(test_se), 
        .CLK(n1920), .Q(\mem2[201][22] ), .QN(n30130) );
  SDFFX1 \mem2_reg[201][21]  ( .D(n12025), .SI(\mem2[201][20] ), .SE(test_se), 
        .CLK(n1920), .Q(\mem2[201][21] ), .QN(n30131) );
  SDFFX1 \mem2_reg[201][20]  ( .D(n12024), .SI(\mem2[201][19] ), .SE(test_se), 
        .CLK(n1920), .Q(\mem2[201][20] ), .QN(n30132) );
  SDFFX1 \mem2_reg[201][19]  ( .D(n12023), .SI(\mem2[201][18] ), .SE(test_se), 
        .CLK(n1920), .Q(\mem2[201][19] ), .QN(n30133) );
  SDFFX1 \mem2_reg[201][18]  ( .D(n12022), .SI(\mem2[201][17] ), .SE(test_se), 
        .CLK(n1920), .Q(\mem2[201][18] ), .QN(n30134) );
  SDFFX1 \mem2_reg[201][17]  ( .D(n12021), .SI(\mem2[201][16] ), .SE(test_se), 
        .CLK(n1921), .Q(\mem2[201][17] ), .QN(n30135) );
  SDFFX1 \mem2_reg[201][16]  ( .D(n12020), .SI(\mem2[200][23] ), .SE(test_se), 
        .CLK(n1921), .Q(\mem2[201][16] ), .QN(n30136) );
  SDFFX1 \mem2_reg[200][23]  ( .D(n12019), .SI(\mem2[200][22] ), .SE(test_se), 
        .CLK(n1921), .Q(\mem2[200][23] ), .QN(n30137) );
  SDFFX1 \mem2_reg[200][22]  ( .D(n12018), .SI(\mem2[200][21] ), .SE(test_se), 
        .CLK(n1921), .Q(\mem2[200][22] ), .QN(n30138) );
  SDFFX1 \mem2_reg[200][21]  ( .D(n12017), .SI(\mem2[200][20] ), .SE(test_se), 
        .CLK(n1921), .Q(\mem2[200][21] ), .QN(n30139) );
  SDFFX1 \mem2_reg[200][20]  ( .D(n12016), .SI(\mem2[200][19] ), .SE(test_se), 
        .CLK(n1921), .Q(\mem2[200][20] ), .QN(n30140) );
  SDFFX1 \mem2_reg[200][19]  ( .D(n12015), .SI(\mem2[200][18] ), .SE(test_se), 
        .CLK(n1921), .Q(\mem2[200][19] ), .QN(n30141) );
  SDFFX1 \mem2_reg[200][18]  ( .D(n12014), .SI(\mem2[200][17] ), .SE(test_se), 
        .CLK(n1921), .Q(\mem2[200][18] ), .QN(n30142) );
  SDFFX1 \mem2_reg[200][17]  ( .D(n12013), .SI(\mem2[200][16] ), .SE(test_se), 
        .CLK(n1921), .Q(\mem2[200][17] ), .QN(n30143) );
  SDFFX1 \mem2_reg[200][16]  ( .D(n12012), .SI(\mem2[199][23] ), .SE(test_se), 
        .CLK(n1921), .Q(\mem2[200][16] ), .QN(n30144) );
  SDFFX1 \mem2_reg[199][23]  ( .D(n12011), .SI(\mem2[199][22] ), .SE(test_se), 
        .CLK(n1921), .Q(\mem2[199][23] ), .QN(n30145) );
  SDFFX1 \mem2_reg[199][22]  ( .D(n12010), .SI(\mem2[199][21] ), .SE(test_se), 
        .CLK(n1921), .Q(\mem2[199][22] ), .QN(n30146) );
  SDFFX1 \mem2_reg[199][21]  ( .D(n12009), .SI(\mem2[199][20] ), .SE(test_se), 
        .CLK(n1922), .Q(\mem2[199][21] ), .QN(n30147) );
  SDFFX1 \mem2_reg[199][20]  ( .D(n12008), .SI(\mem2[199][19] ), .SE(test_se), 
        .CLK(n1922), .Q(\mem2[199][20] ), .QN(n30148) );
  SDFFX1 \mem2_reg[199][19]  ( .D(n12007), .SI(\mem2[199][18] ), .SE(test_se), 
        .CLK(n1922), .Q(\mem2[199][19] ), .QN(n30149) );
  SDFFX1 \mem2_reg[199][18]  ( .D(n12006), .SI(\mem2[199][17] ), .SE(test_se), 
        .CLK(n1922), .Q(\mem2[199][18] ), .QN(n30150) );
  SDFFX1 \mem2_reg[199][17]  ( .D(n12005), .SI(\mem2[199][16] ), .SE(test_se), 
        .CLK(n1922), .Q(\mem2[199][17] ), .QN(n30151) );
  SDFFX1 \mem2_reg[199][16]  ( .D(n12004), .SI(\mem2[198][23] ), .SE(test_se), 
        .CLK(n1922), .Q(\mem2[199][16] ), .QN(n30152) );
  SDFFX1 \mem2_reg[198][23]  ( .D(n12003), .SI(\mem2[198][22] ), .SE(test_se), 
        .CLK(n1922), .Q(\mem2[198][23] ), .QN(n30153) );
  SDFFX1 \mem2_reg[198][22]  ( .D(n12002), .SI(\mem2[198][21] ), .SE(test_se), 
        .CLK(n1922), .Q(\mem2[198][22] ), .QN(n30154) );
  SDFFX1 \mem2_reg[198][21]  ( .D(n12001), .SI(\mem2[198][20] ), .SE(test_se), 
        .CLK(n1922), .Q(\mem2[198][21] ), .QN(n30155) );
  SDFFX1 \mem2_reg[198][20]  ( .D(n12000), .SI(\mem2[198][19] ), .SE(test_se), 
        .CLK(n1922), .Q(\mem2[198][20] ), .QN(n30156) );
  SDFFX1 \mem2_reg[198][19]  ( .D(n11999), .SI(\mem2[198][18] ), .SE(test_se), 
        .CLK(n1922), .Q(\mem2[198][19] ), .QN(n30157) );
  SDFFX1 \mem2_reg[198][18]  ( .D(n11998), .SI(\mem2[198][17] ), .SE(test_se), 
        .CLK(n1922), .Q(\mem2[198][18] ), .QN(n30158) );
  SDFFX1 \mem2_reg[198][17]  ( .D(n11997), .SI(\mem2[198][16] ), .SE(test_se), 
        .CLK(n1923), .Q(\mem2[198][17] ), .QN(n30159) );
  SDFFX1 \mem2_reg[198][16]  ( .D(n11996), .SI(\mem2[197][23] ), .SE(test_se), 
        .CLK(n1923), .Q(\mem2[198][16] ), .QN(n30160) );
  SDFFX1 \mem2_reg[197][23]  ( .D(n11995), .SI(\mem2[197][22] ), .SE(test_se), 
        .CLK(n1923), .Q(\mem2[197][23] ), .QN(n30161) );
  SDFFX1 \mem2_reg[197][22]  ( .D(n11994), .SI(\mem2[197][21] ), .SE(test_se), 
        .CLK(n1923), .Q(\mem2[197][22] ), .QN(n30162) );
  SDFFX1 \mem2_reg[197][21]  ( .D(n11993), .SI(\mem2[197][20] ), .SE(test_se), 
        .CLK(n1923), .Q(\mem2[197][21] ), .QN(n30163) );
  SDFFX1 \mem2_reg[197][20]  ( .D(n11992), .SI(\mem2[197][19] ), .SE(test_se), 
        .CLK(n1923), .Q(\mem2[197][20] ), .QN(n30164) );
  SDFFX1 \mem2_reg[197][19]  ( .D(n11991), .SI(\mem2[197][18] ), .SE(test_se), 
        .CLK(n1923), .Q(\mem2[197][19] ), .QN(n30165) );
  SDFFX1 \mem2_reg[197][18]  ( .D(n11990), .SI(\mem2[197][17] ), .SE(test_se), 
        .CLK(n1923), .Q(\mem2[197][18] ), .QN(n30166) );
  SDFFX1 \mem2_reg[197][17]  ( .D(n11989), .SI(\mem2[197][16] ), .SE(test_se), 
        .CLK(n1923), .Q(\mem2[197][17] ), .QN(n30167) );
  SDFFX1 \mem2_reg[197][16]  ( .D(n11988), .SI(\mem2[196][23] ), .SE(test_se), 
        .CLK(n1923), .Q(\mem2[197][16] ), .QN(n30168) );
  SDFFX1 \mem2_reg[196][23]  ( .D(n11987), .SI(\mem2[196][22] ), .SE(test_se), 
        .CLK(n1923), .Q(\mem2[196][23] ), .QN(n30169) );
  SDFFX1 \mem2_reg[196][22]  ( .D(n11986), .SI(\mem2[196][21] ), .SE(test_se), 
        .CLK(n1923), .Q(\mem2[196][22] ), .QN(n30170) );
  SDFFX1 \mem2_reg[196][21]  ( .D(n11985), .SI(\mem2[196][20] ), .SE(test_se), 
        .CLK(n1924), .Q(\mem2[196][21] ), .QN(n30171) );
  SDFFX1 \mem2_reg[196][20]  ( .D(n11984), .SI(\mem2[196][19] ), .SE(test_se), 
        .CLK(n1924), .Q(\mem2[196][20] ), .QN(n30172) );
  SDFFX1 \mem2_reg[196][19]  ( .D(n11983), .SI(\mem2[196][18] ), .SE(test_se), 
        .CLK(n1924), .Q(\mem2[196][19] ), .QN(n30173) );
  SDFFX1 \mem2_reg[196][18]  ( .D(n11982), .SI(\mem2[196][17] ), .SE(test_se), 
        .CLK(n1924), .Q(\mem2[196][18] ), .QN(n30174) );
  SDFFX1 \mem2_reg[196][17]  ( .D(n11981), .SI(\mem2[196][16] ), .SE(test_se), 
        .CLK(n1924), .Q(\mem2[196][17] ), .QN(n30175) );
  SDFFX1 \mem2_reg[196][16]  ( .D(n11980), .SI(\mem2[195][23] ), .SE(test_se), 
        .CLK(n1924), .Q(\mem2[196][16] ), .QN(n30176) );
  SDFFX1 \mem2_reg[195][23]  ( .D(n11979), .SI(\mem2[195][22] ), .SE(test_se), 
        .CLK(n1924), .Q(\mem2[195][23] ), .QN(n30177) );
  SDFFX1 \mem2_reg[195][22]  ( .D(n11978), .SI(\mem2[195][21] ), .SE(test_se), 
        .CLK(n1924), .Q(\mem2[195][22] ), .QN(n30178) );
  SDFFX1 \mem2_reg[195][21]  ( .D(n11977), .SI(\mem2[195][20] ), .SE(test_se), 
        .CLK(n1924), .Q(\mem2[195][21] ), .QN(n30179) );
  SDFFX1 \mem2_reg[195][20]  ( .D(n11976), .SI(\mem2[195][19] ), .SE(test_se), 
        .CLK(n1924), .Q(\mem2[195][20] ), .QN(n30180) );
  SDFFX1 \mem2_reg[195][19]  ( .D(n11975), .SI(\mem2[195][18] ), .SE(test_se), 
        .CLK(n1924), .Q(\mem2[195][19] ), .QN(n30181) );
  SDFFX1 \mem2_reg[195][18]  ( .D(n11974), .SI(\mem2[195][17] ), .SE(test_se), 
        .CLK(n1924), .Q(\mem2[195][18] ), .QN(n30182) );
  SDFFX1 \mem2_reg[195][17]  ( .D(n11973), .SI(\mem2[195][16] ), .SE(test_se), 
        .CLK(n1925), .Q(\mem2[195][17] ), .QN(n30183) );
  SDFFX1 \mem2_reg[195][16]  ( .D(n11972), .SI(\mem2[194][23] ), .SE(test_se), 
        .CLK(n1925), .Q(\mem2[195][16] ), .QN(n30184) );
  SDFFX1 \mem2_reg[194][23]  ( .D(n11971), .SI(\mem2[194][22] ), .SE(test_se), 
        .CLK(n1925), .Q(\mem2[194][23] ), .QN(n30185) );
  SDFFX1 \mem2_reg[194][22]  ( .D(n11970), .SI(\mem2[194][21] ), .SE(test_se), 
        .CLK(n1925), .Q(\mem2[194][22] ), .QN(n30186) );
  SDFFX1 \mem2_reg[194][21]  ( .D(n11969), .SI(\mem2[194][20] ), .SE(test_se), 
        .CLK(n1925), .Q(\mem2[194][21] ), .QN(n30187) );
  SDFFX1 \mem2_reg[194][20]  ( .D(n11968), .SI(\mem2[194][19] ), .SE(test_se), 
        .CLK(n1925), .Q(\mem2[194][20] ), .QN(n30188) );
  SDFFX1 \mem2_reg[194][19]  ( .D(n11967), .SI(\mem2[194][18] ), .SE(test_se), 
        .CLK(n1925), .Q(\mem2[194][19] ), .QN(n30189) );
  SDFFX1 \mem2_reg[194][18]  ( .D(n11966), .SI(\mem2[194][17] ), .SE(test_se), 
        .CLK(n1925), .Q(\mem2[194][18] ), .QN(n30190) );
  SDFFX1 \mem2_reg[194][17]  ( .D(n11965), .SI(\mem2[194][16] ), .SE(test_se), 
        .CLK(n1925), .Q(\mem2[194][17] ), .QN(n30191) );
  SDFFX1 \mem2_reg[194][16]  ( .D(n11964), .SI(\mem2[193][23] ), .SE(test_se), 
        .CLK(n1925), .Q(\mem2[194][16] ), .QN(n30192) );
  SDFFX1 \mem2_reg[193][23]  ( .D(n11963), .SI(\mem2[193][22] ), .SE(test_se), 
        .CLK(n1925), .Q(\mem2[193][23] ), .QN(n30193) );
  SDFFX1 \mem2_reg[193][22]  ( .D(n11962), .SI(\mem2[193][21] ), .SE(test_se), 
        .CLK(n1925), .Q(\mem2[193][22] ), .QN(n30194) );
  SDFFX1 \mem2_reg[193][21]  ( .D(n11961), .SI(\mem2[193][20] ), .SE(test_se), 
        .CLK(n1926), .Q(\mem2[193][21] ), .QN(n30195) );
  SDFFX1 \mem2_reg[193][20]  ( .D(n11960), .SI(\mem2[193][19] ), .SE(test_se), 
        .CLK(n1926), .Q(\mem2[193][20] ), .QN(n30196) );
  SDFFX1 \mem2_reg[193][19]  ( .D(n11959), .SI(\mem2[193][18] ), .SE(test_se), 
        .CLK(n1926), .Q(\mem2[193][19] ), .QN(n30197) );
  SDFFX1 \mem2_reg[193][18]  ( .D(n11958), .SI(\mem2[193][17] ), .SE(test_se), 
        .CLK(n1926), .Q(\mem2[193][18] ), .QN(n30198) );
  SDFFX1 \mem2_reg[193][17]  ( .D(n11957), .SI(\mem2[193][16] ), .SE(test_se), 
        .CLK(n1926), .Q(\mem2[193][17] ), .QN(n30199) );
  SDFFX1 \mem2_reg[193][16]  ( .D(n11956), .SI(\mem2[192][23] ), .SE(test_se), 
        .CLK(n1926), .Q(\mem2[193][16] ), .QN(n30200) );
  SDFFX1 \mem2_reg[192][23]  ( .D(n11955), .SI(\mem2[192][22] ), .SE(test_se), 
        .CLK(n1926), .Q(\mem2[192][23] ), .QN(n30201) );
  SDFFX1 \mem2_reg[192][22]  ( .D(n11954), .SI(\mem2[192][21] ), .SE(test_se), 
        .CLK(n1926), .Q(\mem2[192][22] ), .QN(n30202) );
  SDFFX1 \mem2_reg[192][21]  ( .D(n11953), .SI(\mem2[192][20] ), .SE(test_se), 
        .CLK(n1926), .Q(\mem2[192][21] ), .QN(n30203) );
  SDFFX1 \mem2_reg[192][20]  ( .D(n11952), .SI(\mem2[192][19] ), .SE(test_se), 
        .CLK(n1926), .Q(\mem2[192][20] ), .QN(n30204) );
  SDFFX1 \mem2_reg[192][19]  ( .D(n11951), .SI(\mem2[192][18] ), .SE(test_se), 
        .CLK(n1926), .Q(\mem2[192][19] ), .QN(n30205) );
  SDFFX1 \mem2_reg[192][18]  ( .D(n11950), .SI(\mem2[192][17] ), .SE(test_se), 
        .CLK(n1926), .Q(\mem2[192][18] ), .QN(n30206) );
  SDFFX1 \mem2_reg[192][17]  ( .D(n11949), .SI(\mem2[192][16] ), .SE(test_se), 
        .CLK(n1927), .Q(\mem2[192][17] ), .QN(n30207) );
  SDFFX1 \mem2_reg[192][16]  ( .D(n11948), .SI(\mem2[191][23] ), .SE(test_se), 
        .CLK(n1927), .Q(\mem2[192][16] ), .QN(n30208) );
  SDFFX1 \mem2_reg[191][23]  ( .D(n11947), .SI(\mem2[191][22] ), .SE(test_se), 
        .CLK(n1927), .Q(\mem2[191][23] ), .QN(n30209) );
  SDFFX1 \mem2_reg[191][22]  ( .D(n11946), .SI(\mem2[191][21] ), .SE(test_se), 
        .CLK(n1927), .Q(\mem2[191][22] ), .QN(n30210) );
  SDFFX1 \mem2_reg[191][21]  ( .D(n11945), .SI(\mem2[191][20] ), .SE(test_se), 
        .CLK(n1927), .Q(\mem2[191][21] ), .QN(n30211) );
  SDFFX1 \mem2_reg[191][20]  ( .D(n11944), .SI(\mem2[191][19] ), .SE(test_se), 
        .CLK(n1927), .Q(\mem2[191][20] ), .QN(n30212) );
  SDFFX1 \mem2_reg[191][19]  ( .D(n11943), .SI(\mem2[191][18] ), .SE(test_se), 
        .CLK(n1927), .Q(\mem2[191][19] ), .QN(n30213) );
  SDFFX1 \mem2_reg[191][18]  ( .D(n11942), .SI(\mem2[191][17] ), .SE(test_se), 
        .CLK(n1927), .Q(\mem2[191][18] ), .QN(n30214) );
  SDFFX1 \mem2_reg[191][17]  ( .D(n11941), .SI(\mem2[191][16] ), .SE(test_se), 
        .CLK(n1927), .Q(\mem2[191][17] ), .QN(n30215) );
  SDFFX1 \mem2_reg[191][16]  ( .D(n11940), .SI(\mem2[190][23] ), .SE(test_se), 
        .CLK(n1927), .Q(\mem2[191][16] ), .QN(n30216) );
  SDFFX1 \mem2_reg[190][23]  ( .D(n11939), .SI(\mem2[190][22] ), .SE(test_se), 
        .CLK(n1927), .Q(\mem2[190][23] ), .QN(n30217) );
  SDFFX1 \mem2_reg[190][22]  ( .D(n11938), .SI(\mem2[190][21] ), .SE(test_se), 
        .CLK(n1927), .Q(\mem2[190][22] ), .QN(n30218) );
  SDFFX1 \mem2_reg[190][21]  ( .D(n11937), .SI(\mem2[190][20] ), .SE(test_se), 
        .CLK(n1928), .Q(\mem2[190][21] ), .QN(n30219) );
  SDFFX1 \mem2_reg[190][20]  ( .D(n11936), .SI(\mem2[190][19] ), .SE(test_se), 
        .CLK(n1928), .Q(\mem2[190][20] ), .QN(n30220) );
  SDFFX1 \mem2_reg[190][19]  ( .D(n11935), .SI(\mem2[190][18] ), .SE(test_se), 
        .CLK(n1928), .Q(\mem2[190][19] ), .QN(n30221) );
  SDFFX1 \mem2_reg[190][18]  ( .D(n11934), .SI(\mem2[190][17] ), .SE(test_se), 
        .CLK(n1928), .Q(\mem2[190][18] ), .QN(n30222) );
  SDFFX1 \mem2_reg[190][17]  ( .D(n11933), .SI(\mem2[190][16] ), .SE(test_se), 
        .CLK(n1928), .Q(\mem2[190][17] ), .QN(n30223) );
  SDFFX1 \mem2_reg[190][16]  ( .D(n11932), .SI(\mem2[189][23] ), .SE(test_se), 
        .CLK(n1928), .Q(\mem2[190][16] ), .QN(n30224) );
  SDFFX1 \mem2_reg[189][23]  ( .D(n11931), .SI(\mem2[189][22] ), .SE(test_se), 
        .CLK(n1928), .Q(\mem2[189][23] ), .QN(n30225) );
  SDFFX1 \mem2_reg[189][22]  ( .D(n11930), .SI(\mem2[189][21] ), .SE(test_se), 
        .CLK(n1928), .Q(\mem2[189][22] ), .QN(n30226) );
  SDFFX1 \mem2_reg[189][21]  ( .D(n11929), .SI(\mem2[189][20] ), .SE(test_se), 
        .CLK(n1928), .Q(\mem2[189][21] ), .QN(n30227) );
  SDFFX1 \mem2_reg[189][20]  ( .D(n11928), .SI(\mem2[189][19] ), .SE(test_se), 
        .CLK(n1928), .Q(\mem2[189][20] ), .QN(n30228) );
  SDFFX1 \mem2_reg[189][19]  ( .D(n11927), .SI(\mem2[189][18] ), .SE(test_se), 
        .CLK(n1928), .Q(\mem2[189][19] ), .QN(n30229) );
  SDFFX1 \mem2_reg[189][18]  ( .D(n11926), .SI(\mem2[189][17] ), .SE(test_se), 
        .CLK(n1928), .Q(\mem2[189][18] ), .QN(n30230) );
  SDFFX1 \mem2_reg[189][17]  ( .D(n11925), .SI(\mem2[189][16] ), .SE(test_se), 
        .CLK(n1929), .Q(\mem2[189][17] ), .QN(n30231) );
  SDFFX1 \mem2_reg[189][16]  ( .D(n11924), .SI(\mem2[188][23] ), .SE(test_se), 
        .CLK(n1929), .Q(\mem2[189][16] ), .QN(n30232) );
  SDFFX1 \mem2_reg[188][23]  ( .D(n11923), .SI(\mem2[188][22] ), .SE(test_se), 
        .CLK(n1929), .Q(\mem2[188][23] ), .QN(n30233) );
  SDFFX1 \mem2_reg[188][22]  ( .D(n11922), .SI(\mem2[188][21] ), .SE(test_se), 
        .CLK(n1929), .Q(\mem2[188][22] ), .QN(n30234) );
  SDFFX1 \mem2_reg[188][21]  ( .D(n11921), .SI(\mem2[188][20] ), .SE(test_se), 
        .CLK(n1929), .Q(\mem2[188][21] ), .QN(n30235) );
  SDFFX1 \mem2_reg[188][20]  ( .D(n11920), .SI(\mem2[188][19] ), .SE(test_se), 
        .CLK(n1929), .Q(\mem2[188][20] ), .QN(n30236) );
  SDFFX1 \mem2_reg[188][19]  ( .D(n11919), .SI(\mem2[188][18] ), .SE(test_se), 
        .CLK(n1929), .Q(\mem2[188][19] ), .QN(n30237) );
  SDFFX1 \mem2_reg[188][18]  ( .D(n11918), .SI(\mem2[188][17] ), .SE(test_se), 
        .CLK(n1929), .Q(\mem2[188][18] ), .QN(n30238) );
  SDFFX1 \mem2_reg[188][17]  ( .D(n11917), .SI(\mem2[188][16] ), .SE(test_se), 
        .CLK(n1929), .Q(\mem2[188][17] ), .QN(n30239) );
  SDFFX1 \mem2_reg[188][16]  ( .D(n11916), .SI(\mem2[187][23] ), .SE(test_se), 
        .CLK(n1929), .Q(\mem2[188][16] ), .QN(n30240) );
  SDFFX1 \mem2_reg[187][23]  ( .D(n11915), .SI(\mem2[187][22] ), .SE(test_se), 
        .CLK(n1929), .Q(\mem2[187][23] ), .QN(n30241) );
  SDFFX1 \mem2_reg[187][22]  ( .D(n11914), .SI(\mem2[187][21] ), .SE(test_se), 
        .CLK(n1929), .Q(\mem2[187][22] ), .QN(n30242) );
  SDFFX1 \mem2_reg[187][21]  ( .D(n11913), .SI(\mem2[187][20] ), .SE(test_se), 
        .CLK(n1930), .Q(\mem2[187][21] ), .QN(n30243) );
  SDFFX1 \mem2_reg[187][20]  ( .D(n11912), .SI(\mem2[187][19] ), .SE(test_se), 
        .CLK(n1930), .Q(\mem2[187][20] ), .QN(n30244) );
  SDFFX1 \mem2_reg[187][19]  ( .D(n11911), .SI(\mem2[187][18] ), .SE(test_se), 
        .CLK(n1930), .Q(\mem2[187][19] ), .QN(n30245) );
  SDFFX1 \mem2_reg[187][18]  ( .D(n11910), .SI(\mem2[187][17] ), .SE(test_se), 
        .CLK(n1930), .Q(\mem2[187][18] ), .QN(n30246) );
  SDFFX1 \mem2_reg[187][17]  ( .D(n11909), .SI(\mem2[187][16] ), .SE(test_se), 
        .CLK(n1930), .Q(\mem2[187][17] ), .QN(n30247) );
  SDFFX1 \mem2_reg[187][16]  ( .D(n11908), .SI(\mem2[186][23] ), .SE(test_se), 
        .CLK(n1930), .Q(\mem2[187][16] ), .QN(n30248) );
  SDFFX1 \mem2_reg[186][23]  ( .D(n11907), .SI(\mem2[186][22] ), .SE(test_se), 
        .CLK(n1930), .Q(\mem2[186][23] ), .QN(n30249) );
  SDFFX1 \mem2_reg[186][22]  ( .D(n11906), .SI(\mem2[186][21] ), .SE(test_se), 
        .CLK(n1930), .Q(\mem2[186][22] ), .QN(n30250) );
  SDFFX1 \mem2_reg[186][21]  ( .D(n11905), .SI(\mem2[186][20] ), .SE(test_se), 
        .CLK(n1930), .Q(\mem2[186][21] ), .QN(n30251) );
  SDFFX1 \mem2_reg[186][20]  ( .D(n11904), .SI(\mem2[186][19] ), .SE(test_se), 
        .CLK(n1930), .Q(\mem2[186][20] ), .QN(n30252) );
  SDFFX1 \mem2_reg[186][19]  ( .D(n11903), .SI(\mem2[186][18] ), .SE(test_se), 
        .CLK(n1930), .Q(\mem2[186][19] ), .QN(n30253) );
  SDFFX1 \mem2_reg[186][18]  ( .D(n11902), .SI(\mem2[186][17] ), .SE(test_se), 
        .CLK(n1930), .Q(\mem2[186][18] ), .QN(n30254) );
  SDFFX1 \mem2_reg[186][17]  ( .D(n11901), .SI(\mem2[186][16] ), .SE(test_se), 
        .CLK(n1931), .Q(\mem2[186][17] ), .QN(n30255) );
  SDFFX1 \mem2_reg[186][16]  ( .D(n11900), .SI(\mem2[185][23] ), .SE(test_se), 
        .CLK(n1931), .Q(\mem2[186][16] ), .QN(n30256) );
  SDFFX1 \mem2_reg[185][23]  ( .D(n11899), .SI(\mem2[185][22] ), .SE(test_se), 
        .CLK(n1931), .Q(\mem2[185][23] ), .QN(n30257) );
  SDFFX1 \mem2_reg[185][22]  ( .D(n11898), .SI(\mem2[185][21] ), .SE(test_se), 
        .CLK(n1931), .Q(\mem2[185][22] ), .QN(n30258) );
  SDFFX1 \mem2_reg[185][21]  ( .D(n11897), .SI(\mem2[185][20] ), .SE(test_se), 
        .CLK(n1931), .Q(\mem2[185][21] ), .QN(n30259) );
  SDFFX1 \mem2_reg[185][20]  ( .D(n11896), .SI(\mem2[185][19] ), .SE(test_se), 
        .CLK(n1931), .Q(\mem2[185][20] ), .QN(n30260) );
  SDFFX1 \mem2_reg[185][19]  ( .D(n11895), .SI(\mem2[185][18] ), .SE(test_se), 
        .CLK(n1931), .Q(\mem2[185][19] ), .QN(n30261) );
  SDFFX1 \mem2_reg[185][18]  ( .D(n11894), .SI(\mem2[185][17] ), .SE(test_se), 
        .CLK(n1931), .Q(\mem2[185][18] ), .QN(n30262) );
  SDFFX1 \mem2_reg[185][17]  ( .D(n11893), .SI(\mem2[185][16] ), .SE(test_se), 
        .CLK(n1931), .Q(\mem2[185][17] ), .QN(n30263) );
  SDFFX1 \mem2_reg[185][16]  ( .D(n11892), .SI(\mem2[184][23] ), .SE(test_se), 
        .CLK(n1931), .Q(\mem2[185][16] ), .QN(n30264) );
  SDFFX1 \mem2_reg[184][23]  ( .D(n11891), .SI(\mem2[184][22] ), .SE(test_se), 
        .CLK(n1931), .Q(\mem2[184][23] ), .QN(n30265) );
  SDFFX1 \mem2_reg[184][22]  ( .D(n11890), .SI(\mem2[184][21] ), .SE(test_se), 
        .CLK(n1931), .Q(\mem2[184][22] ), .QN(n30266) );
  SDFFX1 \mem2_reg[184][21]  ( .D(n11889), .SI(\mem2[184][20] ), .SE(test_se), 
        .CLK(n1932), .Q(\mem2[184][21] ), .QN(n30267) );
  SDFFX1 \mem2_reg[184][20]  ( .D(n11888), .SI(\mem2[184][19] ), .SE(test_se), 
        .CLK(n1932), .Q(\mem2[184][20] ), .QN(n30268) );
  SDFFX1 \mem2_reg[184][19]  ( .D(n11887), .SI(\mem2[184][18] ), .SE(test_se), 
        .CLK(n1932), .Q(\mem2[184][19] ), .QN(n30269) );
  SDFFX1 \mem2_reg[184][18]  ( .D(n11886), .SI(\mem2[184][17] ), .SE(test_se), 
        .CLK(n1932), .Q(\mem2[184][18] ), .QN(n30270) );
  SDFFX1 \mem2_reg[184][17]  ( .D(n11885), .SI(\mem2[184][16] ), .SE(test_se), 
        .CLK(n1932), .Q(\mem2[184][17] ), .QN(n30271) );
  SDFFX1 \mem2_reg[184][16]  ( .D(n11884), .SI(\mem2[183][23] ), .SE(test_se), 
        .CLK(n1932), .Q(\mem2[184][16] ), .QN(n30272) );
  SDFFX1 \mem2_reg[183][23]  ( .D(n11883), .SI(\mem2[183][22] ), .SE(test_se), 
        .CLK(n1932), .Q(\mem2[183][23] ), .QN(n30273) );
  SDFFX1 \mem2_reg[183][22]  ( .D(n11882), .SI(\mem2[183][21] ), .SE(test_se), 
        .CLK(n1932), .Q(\mem2[183][22] ), .QN(n30274) );
  SDFFX1 \mem2_reg[183][21]  ( .D(n11881), .SI(\mem2[183][20] ), .SE(test_se), 
        .CLK(n1932), .Q(\mem2[183][21] ), .QN(n30275) );
  SDFFX1 \mem2_reg[183][20]  ( .D(n11880), .SI(\mem2[183][19] ), .SE(test_se), 
        .CLK(n1932), .Q(\mem2[183][20] ), .QN(n30276) );
  SDFFX1 \mem2_reg[183][19]  ( .D(n11879), .SI(\mem2[183][18] ), .SE(test_se), 
        .CLK(n1932), .Q(\mem2[183][19] ), .QN(n30277) );
  SDFFX1 \mem2_reg[183][18]  ( .D(n11878), .SI(\mem2[183][17] ), .SE(test_se), 
        .CLK(n1932), .Q(\mem2[183][18] ), .QN(n30278) );
  SDFFX1 \mem2_reg[183][17]  ( .D(n11877), .SI(\mem2[183][16] ), .SE(test_se), 
        .CLK(n1933), .Q(\mem2[183][17] ), .QN(n30279) );
  SDFFX1 \mem2_reg[183][16]  ( .D(n11876), .SI(\mem2[182][23] ), .SE(test_se), 
        .CLK(n1933), .Q(\mem2[183][16] ), .QN(n30280) );
  SDFFX1 \mem2_reg[182][23]  ( .D(n11875), .SI(\mem2[182][22] ), .SE(test_se), 
        .CLK(n1933), .Q(\mem2[182][23] ), .QN(n30281) );
  SDFFX1 \mem2_reg[182][22]  ( .D(n11874), .SI(\mem2[182][21] ), .SE(test_se), 
        .CLK(n1933), .Q(\mem2[182][22] ), .QN(n30282) );
  SDFFX1 \mem2_reg[182][21]  ( .D(n11873), .SI(\mem2[182][20] ), .SE(test_se), 
        .CLK(n1933), .Q(\mem2[182][21] ), .QN(n30283) );
  SDFFX1 \mem2_reg[182][20]  ( .D(n11872), .SI(\mem2[182][19] ), .SE(test_se), 
        .CLK(n1933), .Q(\mem2[182][20] ), .QN(n30284) );
  SDFFX1 \mem2_reg[182][19]  ( .D(n11871), .SI(\mem2[182][18] ), .SE(test_se), 
        .CLK(n1933), .Q(\mem2[182][19] ), .QN(n30285) );
  SDFFX1 \mem2_reg[182][18]  ( .D(n11870), .SI(\mem2[182][17] ), .SE(test_se), 
        .CLK(n1933), .Q(\mem2[182][18] ), .QN(n30286) );
  SDFFX1 \mem2_reg[182][17]  ( .D(n11869), .SI(\mem2[182][16] ), .SE(test_se), 
        .CLK(n1933), .Q(\mem2[182][17] ), .QN(n30287) );
  SDFFX1 \mem2_reg[182][16]  ( .D(n11868), .SI(\mem2[181][23] ), .SE(test_se), 
        .CLK(n1933), .Q(\mem2[182][16] ), .QN(n30288) );
  SDFFX1 \mem2_reg[181][23]  ( .D(n11867), .SI(\mem2[181][22] ), .SE(test_se), 
        .CLK(n1933), .Q(\mem2[181][23] ), .QN(n30289) );
  SDFFX1 \mem2_reg[181][22]  ( .D(n11866), .SI(\mem2[181][21] ), .SE(test_se), 
        .CLK(n1933), .Q(\mem2[181][22] ), .QN(n30290) );
  SDFFX1 \mem2_reg[181][21]  ( .D(n11865), .SI(\mem2[181][20] ), .SE(test_se), 
        .CLK(n1934), .Q(\mem2[181][21] ), .QN(n30291) );
  SDFFX1 \mem2_reg[181][20]  ( .D(n11864), .SI(\mem2[181][19] ), .SE(test_se), 
        .CLK(n1934), .Q(\mem2[181][20] ), .QN(n30292) );
  SDFFX1 \mem2_reg[181][19]  ( .D(n11863), .SI(\mem2[181][18] ), .SE(test_se), 
        .CLK(n1934), .Q(\mem2[181][19] ), .QN(n30293) );
  SDFFX1 \mem2_reg[181][18]  ( .D(n11862), .SI(\mem2[181][17] ), .SE(test_se), 
        .CLK(n1934), .Q(\mem2[181][18] ), .QN(n30294) );
  SDFFX1 \mem2_reg[181][17]  ( .D(n11861), .SI(\mem2[181][16] ), .SE(test_se), 
        .CLK(n1934), .Q(\mem2[181][17] ), .QN(n30295) );
  SDFFX1 \mem2_reg[181][16]  ( .D(n11860), .SI(\mem2[180][23] ), .SE(test_se), 
        .CLK(n1934), .Q(\mem2[181][16] ), .QN(n30296) );
  SDFFX1 \mem2_reg[180][23]  ( .D(n11859), .SI(\mem2[180][22] ), .SE(test_se), 
        .CLK(n1934), .Q(\mem2[180][23] ), .QN(n30297) );
  SDFFX1 \mem2_reg[180][22]  ( .D(n11858), .SI(\mem2[180][21] ), .SE(test_se), 
        .CLK(n1934), .Q(\mem2[180][22] ), .QN(n30298) );
  SDFFX1 \mem2_reg[180][21]  ( .D(n11857), .SI(\mem2[180][20] ), .SE(test_se), 
        .CLK(n1934), .Q(\mem2[180][21] ), .QN(n30299) );
  SDFFX1 \mem2_reg[180][20]  ( .D(n11856), .SI(\mem2[180][19] ), .SE(test_se), 
        .CLK(n1934), .Q(\mem2[180][20] ), .QN(n30300) );
  SDFFX1 \mem2_reg[180][19]  ( .D(n11855), .SI(\mem2[180][18] ), .SE(test_se), 
        .CLK(n1934), .Q(\mem2[180][19] ), .QN(n30301) );
  SDFFX1 \mem2_reg[180][18]  ( .D(n11854), .SI(\mem2[180][17] ), .SE(test_se), 
        .CLK(n1934), .Q(\mem2[180][18] ), .QN(n30302) );
  SDFFX1 \mem2_reg[180][17]  ( .D(n11853), .SI(\mem2[180][16] ), .SE(test_se), 
        .CLK(n1935), .Q(\mem2[180][17] ), .QN(n30303) );
  SDFFX1 \mem2_reg[180][16]  ( .D(n11852), .SI(\mem2[179][23] ), .SE(test_se), 
        .CLK(n1935), .Q(\mem2[180][16] ), .QN(n30304) );
  SDFFX1 \mem2_reg[179][23]  ( .D(n11851), .SI(\mem2[179][22] ), .SE(test_se), 
        .CLK(n1935), .Q(\mem2[179][23] ), .QN(n30305) );
  SDFFX1 \mem2_reg[179][22]  ( .D(n11850), .SI(\mem2[179][21] ), .SE(test_se), 
        .CLK(n1935), .Q(\mem2[179][22] ), .QN(n30306) );
  SDFFX1 \mem2_reg[179][21]  ( .D(n11849), .SI(\mem2[179][20] ), .SE(test_se), 
        .CLK(n1935), .Q(\mem2[179][21] ), .QN(n30307) );
  SDFFX1 \mem2_reg[179][20]  ( .D(n11848), .SI(\mem2[179][19] ), .SE(test_se), 
        .CLK(n1935), .Q(\mem2[179][20] ), .QN(n30308) );
  SDFFX1 \mem2_reg[179][19]  ( .D(n11847), .SI(\mem2[179][18] ), .SE(test_se), 
        .CLK(n1935), .Q(\mem2[179][19] ), .QN(n30309) );
  SDFFX1 \mem2_reg[179][18]  ( .D(n11846), .SI(\mem2[179][17] ), .SE(test_se), 
        .CLK(n1935), .Q(\mem2[179][18] ), .QN(n30310) );
  SDFFX1 \mem2_reg[179][17]  ( .D(n11845), .SI(\mem2[179][16] ), .SE(test_se), 
        .CLK(n1935), .Q(\mem2[179][17] ), .QN(n30311) );
  SDFFX1 \mem2_reg[179][16]  ( .D(n11844), .SI(\mem2[178][23] ), .SE(test_se), 
        .CLK(n1935), .Q(\mem2[179][16] ), .QN(n30312) );
  SDFFX1 \mem2_reg[178][23]  ( .D(n11843), .SI(\mem2[178][22] ), .SE(test_se), 
        .CLK(n1935), .Q(\mem2[178][23] ), .QN(n30313) );
  SDFFX1 \mem2_reg[178][22]  ( .D(n11842), .SI(\mem2[178][21] ), .SE(test_se), 
        .CLK(n1935), .Q(\mem2[178][22] ), .QN(n30314) );
  SDFFX1 \mem2_reg[178][21]  ( .D(n11841), .SI(\mem2[178][20] ), .SE(test_se), 
        .CLK(n1936), .Q(\mem2[178][21] ), .QN(n30315) );
  SDFFX1 \mem2_reg[178][20]  ( .D(n11840), .SI(\mem2[178][19] ), .SE(test_se), 
        .CLK(n1936), .Q(\mem2[178][20] ), .QN(n30316) );
  SDFFX1 \mem2_reg[178][19]  ( .D(n11839), .SI(\mem2[178][18] ), .SE(test_se), 
        .CLK(n1936), .Q(\mem2[178][19] ), .QN(n30317) );
  SDFFX1 \mem2_reg[178][18]  ( .D(n11838), .SI(\mem2[178][17] ), .SE(test_se), 
        .CLK(n1936), .Q(\mem2[178][18] ), .QN(n30318) );
  SDFFX1 \mem2_reg[178][17]  ( .D(n11837), .SI(\mem2[178][16] ), .SE(test_se), 
        .CLK(n1936), .Q(\mem2[178][17] ), .QN(n30319) );
  SDFFX1 \mem2_reg[178][16]  ( .D(n11836), .SI(\mem2[177][23] ), .SE(test_se), 
        .CLK(n1936), .Q(\mem2[178][16] ), .QN(n30320) );
  SDFFX1 \mem2_reg[177][23]  ( .D(n11835), .SI(\mem2[177][22] ), .SE(test_se), 
        .CLK(n1936), .Q(\mem2[177][23] ), .QN(n30321) );
  SDFFX1 \mem2_reg[177][22]  ( .D(n11834), .SI(\mem2[177][21] ), .SE(test_se), 
        .CLK(n1936), .Q(\mem2[177][22] ), .QN(n30322) );
  SDFFX1 \mem2_reg[177][21]  ( .D(n11833), .SI(\mem2[177][20] ), .SE(test_se), 
        .CLK(n1936), .Q(\mem2[177][21] ), .QN(n30323) );
  SDFFX1 \mem2_reg[177][20]  ( .D(n11832), .SI(\mem2[177][19] ), .SE(test_se), 
        .CLK(n1936), .Q(\mem2[177][20] ), .QN(n30324) );
  SDFFX1 \mem2_reg[177][19]  ( .D(n11831), .SI(\mem2[177][18] ), .SE(test_se), 
        .CLK(n1936), .Q(\mem2[177][19] ), .QN(n30325) );
  SDFFX1 \mem2_reg[177][18]  ( .D(n11830), .SI(\mem2[177][17] ), .SE(test_se), 
        .CLK(n1936), .Q(\mem2[177][18] ), .QN(n30326) );
  SDFFX1 \mem2_reg[177][17]  ( .D(n11829), .SI(\mem2[177][16] ), .SE(test_se), 
        .CLK(n1937), .Q(\mem2[177][17] ), .QN(n30327) );
  SDFFX1 \mem2_reg[177][16]  ( .D(n11828), .SI(\mem2[176][23] ), .SE(test_se), 
        .CLK(n1937), .Q(\mem2[177][16] ), .QN(n30328) );
  SDFFX1 \mem2_reg[176][23]  ( .D(n11827), .SI(\mem2[176][22] ), .SE(test_se), 
        .CLK(n1937), .Q(\mem2[176][23] ), .QN(n30329) );
  SDFFX1 \mem2_reg[176][22]  ( .D(n11826), .SI(\mem2[176][21] ), .SE(test_se), 
        .CLK(n1937), .Q(\mem2[176][22] ), .QN(n30330) );
  SDFFX1 \mem2_reg[176][21]  ( .D(n11825), .SI(\mem2[176][20] ), .SE(test_se), 
        .CLK(n1937), .Q(\mem2[176][21] ), .QN(n30331) );
  SDFFX1 \mem2_reg[176][20]  ( .D(n11824), .SI(\mem2[176][19] ), .SE(test_se), 
        .CLK(n1937), .Q(\mem2[176][20] ), .QN(n30332) );
  SDFFX1 \mem2_reg[176][19]  ( .D(n11823), .SI(\mem2[176][18] ), .SE(test_se), 
        .CLK(n1937), .Q(\mem2[176][19] ), .QN(n30333) );
  SDFFX1 \mem2_reg[176][18]  ( .D(n11822), .SI(\mem2[176][17] ), .SE(test_se), 
        .CLK(n1937), .Q(\mem2[176][18] ), .QN(n30334) );
  SDFFX1 \mem2_reg[176][17]  ( .D(n11821), .SI(\mem2[176][16] ), .SE(test_se), 
        .CLK(n1937), .Q(\mem2[176][17] ), .QN(n30335) );
  SDFFX1 \mem2_reg[176][16]  ( .D(n11820), .SI(\mem2[175][23] ), .SE(test_se), 
        .CLK(n1937), .Q(\mem2[176][16] ), .QN(n30336) );
  SDFFX1 \mem2_reg[175][23]  ( .D(n11819), .SI(\mem2[175][22] ), .SE(test_se), 
        .CLK(n1937), .Q(\mem2[175][23] ), .QN(n30337) );
  SDFFX1 \mem2_reg[175][22]  ( .D(n11818), .SI(\mem2[175][21] ), .SE(test_se), 
        .CLK(n1937), .Q(\mem2[175][22] ), .QN(n30338) );
  SDFFX1 \mem2_reg[175][21]  ( .D(n11817), .SI(\mem2[175][20] ), .SE(test_se), 
        .CLK(n1938), .Q(\mem2[175][21] ), .QN(n30339) );
  SDFFX1 \mem2_reg[175][20]  ( .D(n11816), .SI(\mem2[175][19] ), .SE(test_se), 
        .CLK(n1938), .Q(\mem2[175][20] ), .QN(n30340) );
  SDFFX1 \mem2_reg[175][19]  ( .D(n11815), .SI(\mem2[175][18] ), .SE(test_se), 
        .CLK(n1938), .Q(\mem2[175][19] ), .QN(n30341) );
  SDFFX1 \mem2_reg[175][18]  ( .D(n11814), .SI(\mem2[175][17] ), .SE(test_se), 
        .CLK(n1938), .Q(\mem2[175][18] ), .QN(n30342) );
  SDFFX1 \mem2_reg[175][17]  ( .D(n11813), .SI(\mem2[175][16] ), .SE(test_se), 
        .CLK(n1938), .Q(\mem2[175][17] ), .QN(n30343) );
  SDFFX1 \mem2_reg[175][16]  ( .D(n11812), .SI(\mem2[174][23] ), .SE(test_se), 
        .CLK(n1938), .Q(\mem2[175][16] ), .QN(n30344) );
  SDFFX1 \mem2_reg[174][23]  ( .D(n11811), .SI(\mem2[174][22] ), .SE(test_se), 
        .CLK(n1938), .Q(\mem2[174][23] ), .QN(n30345) );
  SDFFX1 \mem2_reg[174][22]  ( .D(n11810), .SI(\mem2[174][21] ), .SE(test_se), 
        .CLK(n1938), .Q(\mem2[174][22] ), .QN(n30346) );
  SDFFX1 \mem2_reg[174][21]  ( .D(n11809), .SI(\mem2[174][20] ), .SE(test_se), 
        .CLK(n1938), .Q(\mem2[174][21] ), .QN(n30347) );
  SDFFX1 \mem2_reg[174][20]  ( .D(n11808), .SI(\mem2[174][19] ), .SE(test_se), 
        .CLK(n1938), .Q(\mem2[174][20] ), .QN(n30348) );
  SDFFX1 \mem2_reg[174][19]  ( .D(n11807), .SI(\mem2[174][18] ), .SE(test_se), 
        .CLK(n1938), .Q(\mem2[174][19] ), .QN(n30349) );
  SDFFX1 \mem2_reg[174][18]  ( .D(n11806), .SI(\mem2[174][17] ), .SE(test_se), 
        .CLK(n1938), .Q(\mem2[174][18] ), .QN(n30350) );
  SDFFX1 \mem2_reg[174][17]  ( .D(n11805), .SI(\mem2[174][16] ), .SE(test_se), 
        .CLK(n1939), .Q(\mem2[174][17] ), .QN(n30351) );
  SDFFX1 \mem2_reg[174][16]  ( .D(n11804), .SI(\mem2[173][23] ), .SE(test_se), 
        .CLK(n1939), .Q(\mem2[174][16] ), .QN(n30352) );
  SDFFX1 \mem2_reg[173][23]  ( .D(n11803), .SI(\mem2[173][22] ), .SE(test_se), 
        .CLK(n1939), .Q(\mem2[173][23] ), .QN(n30353) );
  SDFFX1 \mem2_reg[173][22]  ( .D(n11802), .SI(\mem2[173][21] ), .SE(test_se), 
        .CLK(n1939), .Q(\mem2[173][22] ), .QN(n30354) );
  SDFFX1 \mem2_reg[173][21]  ( .D(n11801), .SI(\mem2[173][20] ), .SE(test_se), 
        .CLK(n1939), .Q(\mem2[173][21] ), .QN(n30355) );
  SDFFX1 \mem2_reg[173][20]  ( .D(n11800), .SI(\mem2[173][19] ), .SE(test_se), 
        .CLK(n1939), .Q(\mem2[173][20] ), .QN(n30356) );
  SDFFX1 \mem2_reg[173][19]  ( .D(n11799), .SI(\mem2[173][18] ), .SE(test_se), 
        .CLK(n1939), .Q(\mem2[173][19] ), .QN(n30357) );
  SDFFX1 \mem2_reg[173][18]  ( .D(n11798), .SI(\mem2[173][17] ), .SE(test_se), 
        .CLK(n1939), .Q(\mem2[173][18] ), .QN(n30358) );
  SDFFX1 \mem2_reg[173][17]  ( .D(n11797), .SI(\mem2[173][16] ), .SE(test_se), 
        .CLK(n1939), .Q(\mem2[173][17] ), .QN(n30359) );
  SDFFX1 \mem2_reg[173][16]  ( .D(n11796), .SI(\mem2[172][23] ), .SE(test_se), 
        .CLK(n1939), .Q(\mem2[173][16] ), .QN(n30360) );
  SDFFX1 \mem2_reg[172][23]  ( .D(n11795), .SI(\mem2[172][22] ), .SE(test_se), 
        .CLK(n1939), .Q(\mem2[172][23] ), .QN(n30361) );
  SDFFX1 \mem2_reg[172][22]  ( .D(n11794), .SI(\mem2[172][21] ), .SE(test_se), 
        .CLK(n1939), .Q(\mem2[172][22] ), .QN(n30362) );
  SDFFX1 \mem2_reg[172][21]  ( .D(n11793), .SI(\mem2[172][20] ), .SE(test_se), 
        .CLK(n1940), .Q(\mem2[172][21] ), .QN(n30363) );
  SDFFX1 \mem2_reg[172][20]  ( .D(n11792), .SI(\mem2[172][19] ), .SE(test_se), 
        .CLK(n1940), .Q(\mem2[172][20] ), .QN(n30364) );
  SDFFX1 \mem2_reg[172][19]  ( .D(n11791), .SI(\mem2[172][18] ), .SE(test_se), 
        .CLK(n1940), .Q(\mem2[172][19] ), .QN(n30365) );
  SDFFX1 \mem2_reg[172][18]  ( .D(n11790), .SI(\mem2[172][17] ), .SE(test_se), 
        .CLK(n1940), .Q(\mem2[172][18] ), .QN(n30366) );
  SDFFX1 \mem2_reg[172][17]  ( .D(n11789), .SI(\mem2[172][16] ), .SE(test_se), 
        .CLK(n1940), .Q(\mem2[172][17] ), .QN(n30367) );
  SDFFX1 \mem2_reg[172][16]  ( .D(n11788), .SI(\mem2[171][23] ), .SE(test_se), 
        .CLK(n1940), .Q(\mem2[172][16] ), .QN(n30368) );
  SDFFX1 \mem2_reg[171][23]  ( .D(n11787), .SI(\mem2[171][22] ), .SE(test_se), 
        .CLK(n2072), .Q(\mem2[171][23] ), .QN(n30369) );
  SDFFX1 \mem2_reg[171][22]  ( .D(n11786), .SI(\mem2[171][21] ), .SE(test_se), 
        .CLK(n2072), .Q(\mem2[171][22] ), .QN(n30370) );
  SDFFX1 \mem2_reg[171][21]  ( .D(n11785), .SI(\mem2[171][20] ), .SE(test_se), 
        .CLK(n2072), .Q(\mem2[171][21] ), .QN(n30371) );
  SDFFX1 \mem2_reg[171][20]  ( .D(n11784), .SI(\mem2[171][19] ), .SE(test_se), 
        .CLK(n2072), .Q(\mem2[171][20] ), .QN(n30372) );
  SDFFX1 \mem2_reg[171][19]  ( .D(n11783), .SI(\mem2[171][18] ), .SE(test_se), 
        .CLK(n2072), .Q(\mem2[171][19] ), .QN(n30373) );
  SDFFX1 \mem2_reg[171][18]  ( .D(n11782), .SI(\mem2[171][17] ), .SE(test_se), 
        .CLK(n2072), .Q(\mem2[171][18] ), .QN(n30374) );
  SDFFX1 \mem2_reg[171][17]  ( .D(n11781), .SI(\mem2[171][16] ), .SE(test_se), 
        .CLK(n2072), .Q(\mem2[171][17] ), .QN(n30375) );
  SDFFX1 \mem2_reg[171][16]  ( .D(n11780), .SI(\mem2[170][23] ), .SE(test_se), 
        .CLK(n2072), .Q(\mem2[171][16] ), .QN(n30376) );
  SDFFX1 \mem2_reg[170][23]  ( .D(n11779), .SI(\mem2[170][22] ), .SE(test_se), 
        .CLK(n2074), .Q(\mem2[170][23] ), .QN(n30377) );
  SDFFX1 \mem2_reg[170][22]  ( .D(n11778), .SI(\mem2[170][21] ), .SE(test_se), 
        .CLK(n2074), .Q(\mem2[170][22] ), .QN(n30378) );
  SDFFX1 \mem2_reg[170][21]  ( .D(n11777), .SI(\mem2[170][20] ), .SE(test_se), 
        .CLK(n2074), .Q(\mem2[170][21] ), .QN(n30379) );
  SDFFX1 \mem2_reg[170][20]  ( .D(n11776), .SI(\mem2[170][19] ), .SE(test_se), 
        .CLK(n2074), .Q(\mem2[170][20] ), .QN(n30380) );
  SDFFX1 \mem2_reg[170][19]  ( .D(n11775), .SI(\mem2[170][18] ), .SE(test_se), 
        .CLK(n2074), .Q(\mem2[170][19] ), .QN(n30381) );
  SDFFX1 \mem2_reg[170][18]  ( .D(n11774), .SI(\mem2[170][17] ), .SE(test_se), 
        .CLK(n2074), .Q(\mem2[170][18] ), .QN(n30382) );
  SDFFX1 \mem2_reg[170][17]  ( .D(n11773), .SI(\mem2[170][16] ), .SE(test_se), 
        .CLK(n2074), .Q(\mem2[170][17] ), .QN(n30383) );
  SDFFX1 \mem2_reg[170][16]  ( .D(n11772), .SI(\mem2[169][23] ), .SE(test_se), 
        .CLK(n2075), .Q(\mem2[170][16] ), .QN(n30384) );
  SDFFX1 \mem2_reg[169][23]  ( .D(n11771), .SI(\mem2[169][22] ), .SE(test_se), 
        .CLK(n2075), .Q(\mem2[169][23] ), .QN(n30385) );
  SDFFX1 \mem2_reg[169][22]  ( .D(n11770), .SI(\mem2[169][21] ), .SE(test_se), 
        .CLK(n2075), .Q(\mem2[169][22] ), .QN(n30386) );
  SDFFX1 \mem2_reg[169][21]  ( .D(n11769), .SI(\mem2[169][20] ), .SE(test_se), 
        .CLK(n2075), .Q(\mem2[169][21] ), .QN(n30387) );
  SDFFX1 \mem2_reg[169][20]  ( .D(n11768), .SI(\mem2[169][19] ), .SE(test_se), 
        .CLK(n2075), .Q(\mem2[169][20] ), .QN(n30388) );
  SDFFX1 \mem2_reg[169][19]  ( .D(n11767), .SI(\mem2[169][18] ), .SE(test_se), 
        .CLK(n2075), .Q(\mem2[169][19] ), .QN(n30389) );
  SDFFX1 \mem2_reg[169][18]  ( .D(n11766), .SI(\mem2[169][17] ), .SE(test_se), 
        .CLK(n2075), .Q(\mem2[169][18] ), .QN(n30390) );
  SDFFX1 \mem2_reg[169][17]  ( .D(n11765), .SI(\mem2[169][16] ), .SE(test_se), 
        .CLK(n2075), .Q(\mem2[169][17] ), .QN(n30391) );
  SDFFX1 \mem2_reg[169][16]  ( .D(n11764), .SI(test_si6), .SE(test_se), .CLK(
        n2075), .Q(\mem2[169][16] ), .QN(n30392) );
  SDFFX1 \mem2_reg[168][23]  ( .D(n11763), .SI(\mem2[168][22] ), .SE(test_se), 
        .CLK(n1940), .Q(\mem2[168][23] ), .QN(n30393) );
  SDFFX1 \mem2_reg[168][22]  ( .D(n11762), .SI(\mem2[168][21] ), .SE(test_se), 
        .CLK(n1940), .Q(\mem2[168][22] ), .QN(n30394) );
  SDFFX1 \mem2_reg[168][21]  ( .D(n11761), .SI(\mem2[168][20] ), .SE(test_se), 
        .CLK(n1940), .Q(\mem2[168][21] ), .QN(n30395) );
  SDFFX1 \mem2_reg[168][20]  ( .D(n11760), .SI(\mem2[168][19] ), .SE(test_se), 
        .CLK(n1940), .Q(\mem2[168][20] ), .QN(n30396) );
  SDFFX1 \mem2_reg[168][19]  ( .D(n11759), .SI(\mem2[168][18] ), .SE(test_se), 
        .CLK(n1940), .Q(\mem2[168][19] ), .QN(n30397) );
  SDFFX1 \mem2_reg[168][18]  ( .D(n11758), .SI(\mem2[168][17] ), .SE(test_se), 
        .CLK(n1940), .Q(\mem2[168][18] ), .QN(n30398) );
  SDFFX1 \mem2_reg[168][17]  ( .D(n11757), .SI(\mem2[168][16] ), .SE(test_se), 
        .CLK(n1941), .Q(\mem2[168][17] ), .QN(n30399) );
  SDFFX1 \mem2_reg[168][16]  ( .D(n11756), .SI(\mem2[167][23] ), .SE(test_se), 
        .CLK(n1941), .Q(\mem2[168][16] ), .QN(n30400) );
  SDFFX1 \mem2_reg[167][23]  ( .D(n11755), .SI(\mem2[167][22] ), .SE(test_se), 
        .CLK(n1941), .Q(\mem2[167][23] ), .QN(n30401) );
  SDFFX1 \mem2_reg[167][22]  ( .D(n11754), .SI(\mem2[167][21] ), .SE(test_se), 
        .CLK(n1941), .Q(\mem2[167][22] ), .QN(n30402) );
  SDFFX1 \mem2_reg[167][21]  ( .D(n11753), .SI(\mem2[167][20] ), .SE(test_se), 
        .CLK(n1941), .Q(\mem2[167][21] ), .QN(n30403) );
  SDFFX1 \mem2_reg[167][20]  ( .D(n11752), .SI(\mem2[167][19] ), .SE(test_se), 
        .CLK(n1941), .Q(\mem2[167][20] ), .QN(n30404) );
  SDFFX1 \mem2_reg[167][19]  ( .D(n11751), .SI(\mem2[167][18] ), .SE(test_se), 
        .CLK(n1941), .Q(\mem2[167][19] ), .QN(n30405) );
  SDFFX1 \mem2_reg[167][18]  ( .D(n11750), .SI(\mem2[167][17] ), .SE(test_se), 
        .CLK(n1941), .Q(\mem2[167][18] ), .QN(n30406) );
  SDFFX1 \mem2_reg[167][17]  ( .D(n11749), .SI(\mem2[167][16] ), .SE(test_se), 
        .CLK(n1941), .Q(\mem2[167][17] ), .QN(n30407) );
  SDFFX1 \mem2_reg[167][16]  ( .D(n11748), .SI(\mem2[166][23] ), .SE(test_se), 
        .CLK(n1941), .Q(\mem2[167][16] ), .QN(n30408) );
  SDFFX1 \mem2_reg[166][23]  ( .D(n11747), .SI(\mem2[166][22] ), .SE(test_se), 
        .CLK(n1941), .Q(\mem2[166][23] ), .QN(n30409) );
  SDFFX1 \mem2_reg[166][22]  ( .D(n11746), .SI(\mem2[166][21] ), .SE(test_se), 
        .CLK(n1941), .Q(\mem2[166][22] ), .QN(n30410) );
  SDFFX1 \mem2_reg[166][21]  ( .D(n11745), .SI(\mem2[166][20] ), .SE(test_se), 
        .CLK(n1942), .Q(\mem2[166][21] ), .QN(n30411) );
  SDFFX1 \mem2_reg[166][20]  ( .D(n11744), .SI(\mem2[166][19] ), .SE(test_se), 
        .CLK(n1942), .Q(\mem2[166][20] ), .QN(n30412) );
  SDFFX1 \mem2_reg[166][19]  ( .D(n11743), .SI(\mem2[166][18] ), .SE(test_se), 
        .CLK(n1942), .Q(\mem2[166][19] ), .QN(n30413) );
  SDFFX1 \mem2_reg[166][18]  ( .D(n11742), .SI(\mem2[166][17] ), .SE(test_se), 
        .CLK(n1942), .Q(\mem2[166][18] ), .QN(n30414) );
  SDFFX1 \mem2_reg[166][17]  ( .D(n11741), .SI(\mem2[166][16] ), .SE(test_se), 
        .CLK(n1942), .Q(\mem2[166][17] ), .QN(n30415) );
  SDFFX1 \mem2_reg[166][16]  ( .D(n11740), .SI(\mem2[165][23] ), .SE(test_se), 
        .CLK(n1942), .Q(\mem2[166][16] ), .QN(n30416) );
  SDFFX1 \mem2_reg[165][23]  ( .D(n11739), .SI(\mem2[165][22] ), .SE(test_se), 
        .CLK(n1942), .Q(\mem2[165][23] ), .QN(n30417) );
  SDFFX1 \mem2_reg[165][22]  ( .D(n11738), .SI(\mem2[165][21] ), .SE(test_se), 
        .CLK(n1942), .Q(\mem2[165][22] ), .QN(n30418) );
  SDFFX1 \mem2_reg[165][21]  ( .D(n11737), .SI(\mem2[165][20] ), .SE(test_se), 
        .CLK(n1942), .Q(\mem2[165][21] ), .QN(n30419) );
  SDFFX1 \mem2_reg[165][20]  ( .D(n11736), .SI(\mem2[165][19] ), .SE(test_se), 
        .CLK(n1942), .Q(\mem2[165][20] ), .QN(n30420) );
  SDFFX1 \mem2_reg[165][19]  ( .D(n11735), .SI(\mem2[165][18] ), .SE(test_se), 
        .CLK(n1942), .Q(\mem2[165][19] ), .QN(n30421) );
  SDFFX1 \mem2_reg[165][18]  ( .D(n11734), .SI(\mem2[165][17] ), .SE(test_se), 
        .CLK(n1942), .Q(\mem2[165][18] ), .QN(n30422) );
  SDFFX1 \mem2_reg[165][17]  ( .D(n11733), .SI(\mem2[165][16] ), .SE(test_se), 
        .CLK(n1943), .Q(\mem2[165][17] ), .QN(n30423) );
  SDFFX1 \mem2_reg[165][16]  ( .D(n11732), .SI(\mem2[164][23] ), .SE(test_se), 
        .CLK(n1943), .Q(\mem2[165][16] ), .QN(n30424) );
  SDFFX1 \mem2_reg[164][23]  ( .D(n11731), .SI(\mem2[164][22] ), .SE(test_se), 
        .CLK(n1943), .Q(\mem2[164][23] ), .QN(n30425) );
  SDFFX1 \mem2_reg[164][22]  ( .D(n11730), .SI(\mem2[164][21] ), .SE(test_se), 
        .CLK(n1943), .Q(\mem2[164][22] ), .QN(n30426) );
  SDFFX1 \mem2_reg[164][21]  ( .D(n11729), .SI(\mem2[164][20] ), .SE(test_se), 
        .CLK(n1943), .Q(\mem2[164][21] ), .QN(n30427) );
  SDFFX1 \mem2_reg[164][20]  ( .D(n11728), .SI(\mem2[164][19] ), .SE(test_se), 
        .CLK(n1943), .Q(\mem2[164][20] ), .QN(n30428) );
  SDFFX1 \mem2_reg[164][19]  ( .D(n11727), .SI(\mem2[164][18] ), .SE(test_se), 
        .CLK(n1943), .Q(\mem2[164][19] ), .QN(n30429) );
  SDFFX1 \mem2_reg[164][18]  ( .D(n11726), .SI(\mem2[164][17] ), .SE(test_se), 
        .CLK(n1943), .Q(\mem2[164][18] ), .QN(n30430) );
  SDFFX1 \mem2_reg[164][17]  ( .D(n11725), .SI(\mem2[164][16] ), .SE(test_se), 
        .CLK(n1943), .Q(\mem2[164][17] ), .QN(n30431) );
  SDFFX1 \mem2_reg[164][16]  ( .D(n11724), .SI(\mem2[163][23] ), .SE(test_se), 
        .CLK(n1943), .Q(\mem2[164][16] ), .QN(n30432) );
  SDFFX1 \mem2_reg[163][23]  ( .D(n11723), .SI(\mem2[163][22] ), .SE(test_se), 
        .CLK(n1943), .Q(\mem2[163][23] ), .QN(n30433) );
  SDFFX1 \mem2_reg[163][22]  ( .D(n11722), .SI(\mem2[163][21] ), .SE(test_se), 
        .CLK(n1943), .Q(\mem2[163][22] ), .QN(n30434) );
  SDFFX1 \mem2_reg[163][21]  ( .D(n11721), .SI(\mem2[163][20] ), .SE(test_se), 
        .CLK(n1944), .Q(\mem2[163][21] ), .QN(n30435) );
  SDFFX1 \mem2_reg[163][20]  ( .D(n11720), .SI(\mem2[163][19] ), .SE(test_se), 
        .CLK(n1944), .Q(\mem2[163][20] ), .QN(n30436) );
  SDFFX1 \mem2_reg[163][19]  ( .D(n11719), .SI(\mem2[163][18] ), .SE(test_se), 
        .CLK(n1944), .Q(\mem2[163][19] ), .QN(n30437) );
  SDFFX1 \mem2_reg[163][18]  ( .D(n11718), .SI(\mem2[163][17] ), .SE(test_se), 
        .CLK(n1944), .Q(\mem2[163][18] ), .QN(n30438) );
  SDFFX1 \mem2_reg[163][17]  ( .D(n11717), .SI(\mem2[163][16] ), .SE(test_se), 
        .CLK(n1944), .Q(\mem2[163][17] ), .QN(n30439) );
  SDFFX1 \mem2_reg[163][16]  ( .D(n11716), .SI(\mem2[162][23] ), .SE(test_se), 
        .CLK(n1944), .Q(\mem2[163][16] ), .QN(n30440) );
  SDFFX1 \mem2_reg[162][23]  ( .D(n11715), .SI(\mem2[162][22] ), .SE(test_se), 
        .CLK(n1944), .Q(\mem2[162][23] ), .QN(n30441) );
  SDFFX1 \mem2_reg[162][22]  ( .D(n11714), .SI(\mem2[162][21] ), .SE(test_se), 
        .CLK(n1944), .Q(\mem2[162][22] ), .QN(n30442) );
  SDFFX1 \mem2_reg[162][21]  ( .D(n11713), .SI(\mem2[162][20] ), .SE(test_se), 
        .CLK(n1944), .Q(\mem2[162][21] ), .QN(n30443) );
  SDFFX1 \mem2_reg[162][20]  ( .D(n11712), .SI(\mem2[162][19] ), .SE(test_se), 
        .CLK(n1944), .Q(\mem2[162][20] ), .QN(n30444) );
  SDFFX1 \mem2_reg[162][19]  ( .D(n11711), .SI(\mem2[162][18] ), .SE(test_se), 
        .CLK(n1944), .Q(\mem2[162][19] ), .QN(n30445) );
  SDFFX1 \mem2_reg[162][18]  ( .D(n11710), .SI(\mem2[162][17] ), .SE(test_se), 
        .CLK(n1944), .Q(\mem2[162][18] ), .QN(n30446) );
  SDFFX1 \mem2_reg[162][17]  ( .D(n11709), .SI(\mem2[162][16] ), .SE(test_se), 
        .CLK(n1945), .Q(\mem2[162][17] ), .QN(n30447) );
  SDFFX1 \mem2_reg[162][16]  ( .D(n11708), .SI(\mem2[161][23] ), .SE(test_se), 
        .CLK(n1945), .Q(\mem2[162][16] ), .QN(n30448) );
  SDFFX1 \mem2_reg[161][23]  ( .D(n11707), .SI(\mem2[161][22] ), .SE(test_se), 
        .CLK(n1945), .Q(\mem2[161][23] ), .QN(n30449) );
  SDFFX1 \mem2_reg[161][22]  ( .D(n11706), .SI(\mem2[161][21] ), .SE(test_se), 
        .CLK(n1945), .Q(\mem2[161][22] ), .QN(n30450) );
  SDFFX1 \mem2_reg[161][21]  ( .D(n11705), .SI(\mem2[161][20] ), .SE(test_se), 
        .CLK(n1945), .Q(\mem2[161][21] ), .QN(n30451) );
  SDFFX1 \mem2_reg[161][20]  ( .D(n11704), .SI(\mem2[161][19] ), .SE(test_se), 
        .CLK(n1945), .Q(\mem2[161][20] ), .QN(n30452) );
  SDFFX1 \mem2_reg[161][19]  ( .D(n11703), .SI(\mem2[161][18] ), .SE(test_se), 
        .CLK(n1945), .Q(\mem2[161][19] ), .QN(n30453) );
  SDFFX1 \mem2_reg[161][18]  ( .D(n11702), .SI(\mem2[161][17] ), .SE(test_se), 
        .CLK(n1945), .Q(\mem2[161][18] ), .QN(n30454) );
  SDFFX1 \mem2_reg[161][17]  ( .D(n11701), .SI(\mem2[161][16] ), .SE(test_se), 
        .CLK(n1945), .Q(\mem2[161][17] ), .QN(n30455) );
  SDFFX1 \mem2_reg[161][16]  ( .D(n11700), .SI(\mem2[160][23] ), .SE(test_se), 
        .CLK(n1945), .Q(\mem2[161][16] ), .QN(n30456) );
  SDFFX1 \mem2_reg[160][23]  ( .D(n11699), .SI(\mem2[160][22] ), .SE(test_se), 
        .CLK(n1945), .Q(\mem2[160][23] ), .QN(n30457) );
  SDFFX1 \mem2_reg[160][22]  ( .D(n11698), .SI(\mem2[160][21] ), .SE(test_se), 
        .CLK(n1945), .Q(\mem2[160][22] ), .QN(n30458) );
  SDFFX1 \mem2_reg[160][21]  ( .D(n11697), .SI(\mem2[160][20] ), .SE(test_se), 
        .CLK(n1946), .Q(\mem2[160][21] ), .QN(n30459) );
  SDFFX1 \mem2_reg[160][20]  ( .D(n11696), .SI(\mem2[160][19] ), .SE(test_se), 
        .CLK(n1946), .Q(\mem2[160][20] ), .QN(n30460) );
  SDFFX1 \mem2_reg[160][19]  ( .D(n11695), .SI(\mem2[160][18] ), .SE(test_se), 
        .CLK(n1946), .Q(\mem2[160][19] ), .QN(n30461) );
  SDFFX1 \mem2_reg[160][18]  ( .D(n11694), .SI(\mem2[160][17] ), .SE(test_se), 
        .CLK(n1946), .Q(\mem2[160][18] ), .QN(n30462) );
  SDFFX1 \mem2_reg[160][17]  ( .D(n11693), .SI(\mem2[160][16] ), .SE(test_se), 
        .CLK(n1946), .Q(\mem2[160][17] ), .QN(n30463) );
  SDFFX1 \mem2_reg[160][16]  ( .D(n11692), .SI(\mem2[159][23] ), .SE(test_se), 
        .CLK(n1946), .Q(\mem2[160][16] ), .QN(n30464) );
  SDFFX1 \mem2_reg[159][23]  ( .D(n11691), .SI(\mem2[159][22] ), .SE(test_se), 
        .CLK(n1946), .Q(\mem2[159][23] ), .QN(n30465) );
  SDFFX1 \mem2_reg[159][22]  ( .D(n11690), .SI(\mem2[159][21] ), .SE(test_se), 
        .CLK(n1946), .Q(\mem2[159][22] ), .QN(n30466) );
  SDFFX1 \mem2_reg[159][21]  ( .D(n11689), .SI(\mem2[159][20] ), .SE(test_se), 
        .CLK(n1946), .Q(\mem2[159][21] ), .QN(n30467) );
  SDFFX1 \mem2_reg[159][20]  ( .D(n11688), .SI(\mem2[159][19] ), .SE(test_se), 
        .CLK(n1946), .Q(\mem2[159][20] ), .QN(n30468) );
  SDFFX1 \mem2_reg[159][19]  ( .D(n11687), .SI(\mem2[159][18] ), .SE(test_se), 
        .CLK(n1946), .Q(\mem2[159][19] ), .QN(n30469) );
  SDFFX1 \mem2_reg[159][18]  ( .D(n11686), .SI(\mem2[159][17] ), .SE(test_se), 
        .CLK(n1946), .Q(\mem2[159][18] ), .QN(n30470) );
  SDFFX1 \mem2_reg[159][17]  ( .D(n11685), .SI(\mem2[159][16] ), .SE(test_se), 
        .CLK(n1947), .Q(\mem2[159][17] ), .QN(n30471) );
  SDFFX1 \mem2_reg[159][16]  ( .D(n11684), .SI(\mem2[158][23] ), .SE(test_se), 
        .CLK(n1947), .Q(\mem2[159][16] ), .QN(n30472) );
  SDFFX1 \mem2_reg[158][23]  ( .D(n11683), .SI(\mem2[158][22] ), .SE(test_se), 
        .CLK(n1947), .Q(\mem2[158][23] ), .QN(n30473) );
  SDFFX1 \mem2_reg[158][22]  ( .D(n11682), .SI(\mem2[158][21] ), .SE(test_se), 
        .CLK(n1947), .Q(\mem2[158][22] ), .QN(n30474) );
  SDFFX1 \mem2_reg[158][21]  ( .D(n11681), .SI(\mem2[158][20] ), .SE(test_se), 
        .CLK(n1947), .Q(\mem2[158][21] ), .QN(n30475) );
  SDFFX1 \mem2_reg[158][20]  ( .D(n11680), .SI(\mem2[158][19] ), .SE(test_se), 
        .CLK(n1947), .Q(\mem2[158][20] ), .QN(n30476) );
  SDFFX1 \mem2_reg[158][19]  ( .D(n11679), .SI(\mem2[158][18] ), .SE(test_se), 
        .CLK(n1947), .Q(\mem2[158][19] ), .QN(n30477) );
  SDFFX1 \mem2_reg[158][18]  ( .D(n11678), .SI(\mem2[158][17] ), .SE(test_se), 
        .CLK(n1947), .Q(\mem2[158][18] ), .QN(n30478) );
  SDFFX1 \mem2_reg[158][17]  ( .D(n11677), .SI(\mem2[158][16] ), .SE(test_se), 
        .CLK(n1947), .Q(\mem2[158][17] ), .QN(n30479) );
  SDFFX1 \mem2_reg[158][16]  ( .D(n11676), .SI(\mem2[157][23] ), .SE(test_se), 
        .CLK(n1947), .Q(\mem2[158][16] ), .QN(n30480) );
  SDFFX1 \mem2_reg[157][23]  ( .D(n11675), .SI(\mem2[157][22] ), .SE(test_se), 
        .CLK(n1947), .Q(\mem2[157][23] ), .QN(n30481) );
  SDFFX1 \mem2_reg[157][22]  ( .D(n11674), .SI(\mem2[157][21] ), .SE(test_se), 
        .CLK(n1947), .Q(\mem2[157][22] ), .QN(n30482) );
  SDFFX1 \mem2_reg[157][21]  ( .D(n11673), .SI(\mem2[157][20] ), .SE(test_se), 
        .CLK(n1948), .Q(\mem2[157][21] ), .QN(n30483) );
  SDFFX1 \mem2_reg[157][20]  ( .D(n11672), .SI(\mem2[157][19] ), .SE(test_se), 
        .CLK(n1948), .Q(\mem2[157][20] ), .QN(n30484) );
  SDFFX1 \mem2_reg[157][19]  ( .D(n11671), .SI(\mem2[157][18] ), .SE(test_se), 
        .CLK(n1948), .Q(\mem2[157][19] ), .QN(n30485) );
  SDFFX1 \mem2_reg[157][18]  ( .D(n11670), .SI(\mem2[157][17] ), .SE(test_se), 
        .CLK(n1948), .Q(\mem2[157][18] ), .QN(n30486) );
  SDFFX1 \mem2_reg[157][17]  ( .D(n11669), .SI(\mem2[157][16] ), .SE(test_se), 
        .CLK(n1948), .Q(\mem2[157][17] ), .QN(n30487) );
  SDFFX1 \mem2_reg[157][16]  ( .D(n11668), .SI(\mem2[156][23] ), .SE(test_se), 
        .CLK(n1948), .Q(\mem2[157][16] ), .QN(n30488) );
  SDFFX1 \mem2_reg[156][23]  ( .D(n11667), .SI(\mem2[156][22] ), .SE(test_se), 
        .CLK(n1948), .Q(\mem2[156][23] ), .QN(n30489) );
  SDFFX1 \mem2_reg[156][22]  ( .D(n11666), .SI(\mem2[156][21] ), .SE(test_se), 
        .CLK(n1948), .Q(\mem2[156][22] ), .QN(n30490) );
  SDFFX1 \mem2_reg[156][21]  ( .D(n11665), .SI(\mem2[156][20] ), .SE(test_se), 
        .CLK(n1948), .Q(\mem2[156][21] ), .QN(n30491) );
  SDFFX1 \mem2_reg[156][20]  ( .D(n11664), .SI(\mem2[156][19] ), .SE(test_se), 
        .CLK(n1948), .Q(\mem2[156][20] ), .QN(n30492) );
  SDFFX1 \mem2_reg[156][19]  ( .D(n11663), .SI(\mem2[156][18] ), .SE(test_se), 
        .CLK(n1948), .Q(\mem2[156][19] ), .QN(n30493) );
  SDFFX1 \mem2_reg[156][18]  ( .D(n11662), .SI(\mem2[156][17] ), .SE(test_se), 
        .CLK(n1948), .Q(\mem2[156][18] ), .QN(n30494) );
  SDFFX1 \mem2_reg[156][17]  ( .D(n11661), .SI(\mem2[156][16] ), .SE(test_se), 
        .CLK(n1949), .Q(\mem2[156][17] ), .QN(n30495) );
  SDFFX1 \mem2_reg[156][16]  ( .D(n11660), .SI(\mem2[155][23] ), .SE(test_se), 
        .CLK(n1949), .Q(\mem2[156][16] ), .QN(n30496) );
  SDFFX1 \mem2_reg[155][23]  ( .D(n11659), .SI(\mem2[155][22] ), .SE(test_se), 
        .CLK(n1949), .Q(\mem2[155][23] ), .QN(n30497) );
  SDFFX1 \mem2_reg[155][22]  ( .D(n11658), .SI(\mem2[155][21] ), .SE(test_se), 
        .CLK(n1949), .Q(\mem2[155][22] ), .QN(n30498) );
  SDFFX1 \mem2_reg[155][21]  ( .D(n11657), .SI(\mem2[155][20] ), .SE(test_se), 
        .CLK(n1949), .Q(\mem2[155][21] ), .QN(n30499) );
  SDFFX1 \mem2_reg[155][20]  ( .D(n11656), .SI(\mem2[155][19] ), .SE(test_se), 
        .CLK(n1949), .Q(\mem2[155][20] ), .QN(n30500) );
  SDFFX1 \mem2_reg[155][19]  ( .D(n11655), .SI(\mem2[155][18] ), .SE(test_se), 
        .CLK(n1949), .Q(\mem2[155][19] ), .QN(n30501) );
  SDFFX1 \mem2_reg[155][18]  ( .D(n11654), .SI(\mem2[155][17] ), .SE(test_se), 
        .CLK(n1949), .Q(\mem2[155][18] ), .QN(n30502) );
  SDFFX1 \mem2_reg[155][17]  ( .D(n11653), .SI(\mem2[155][16] ), .SE(test_se), 
        .CLK(n1949), .Q(\mem2[155][17] ), .QN(n30503) );
  SDFFX1 \mem2_reg[155][16]  ( .D(n11652), .SI(\mem2[154][23] ), .SE(test_se), 
        .CLK(n1949), .Q(\mem2[155][16] ), .QN(n30504) );
  SDFFX1 \mem2_reg[154][23]  ( .D(n11651), .SI(\mem2[154][22] ), .SE(test_se), 
        .CLK(n1949), .Q(\mem2[154][23] ), .QN(n30505) );
  SDFFX1 \mem2_reg[154][22]  ( .D(n11650), .SI(\mem2[154][21] ), .SE(test_se), 
        .CLK(n1949), .Q(\mem2[154][22] ), .QN(n30506) );
  SDFFX1 \mem2_reg[154][21]  ( .D(n11649), .SI(\mem2[154][20] ), .SE(test_se), 
        .CLK(n1950), .Q(\mem2[154][21] ), .QN(n30507) );
  SDFFX1 \mem2_reg[154][20]  ( .D(n11648), .SI(\mem2[154][19] ), .SE(test_se), 
        .CLK(n1950), .Q(\mem2[154][20] ), .QN(n30508) );
  SDFFX1 \mem2_reg[154][19]  ( .D(n11647), .SI(\mem2[154][18] ), .SE(test_se), 
        .CLK(n1950), .Q(\mem2[154][19] ), .QN(n30509) );
  SDFFX1 \mem2_reg[154][18]  ( .D(n11646), .SI(\mem2[154][17] ), .SE(test_se), 
        .CLK(n1950), .Q(\mem2[154][18] ), .QN(n30510) );
  SDFFX1 \mem2_reg[154][17]  ( .D(n11645), .SI(\mem2[154][16] ), .SE(test_se), 
        .CLK(n1950), .Q(\mem2[154][17] ), .QN(n30511) );
  SDFFX1 \mem2_reg[154][16]  ( .D(n11644), .SI(\mem2[153][23] ), .SE(test_se), 
        .CLK(n1950), .Q(\mem2[154][16] ), .QN(n30512) );
  SDFFX1 \mem2_reg[153][23]  ( .D(n11643), .SI(\mem2[153][22] ), .SE(test_se), 
        .CLK(n1950), .Q(\mem2[153][23] ), .QN(n30513) );
  SDFFX1 \mem2_reg[153][22]  ( .D(n11642), .SI(\mem2[153][21] ), .SE(test_se), 
        .CLK(n1950), .Q(\mem2[153][22] ), .QN(n30514) );
  SDFFX1 \mem2_reg[153][21]  ( .D(n11641), .SI(\mem2[153][20] ), .SE(test_se), 
        .CLK(n1950), .Q(\mem2[153][21] ), .QN(n30515) );
  SDFFX1 \mem2_reg[153][20]  ( .D(n11640), .SI(\mem2[153][19] ), .SE(test_se), 
        .CLK(n1950), .Q(\mem2[153][20] ), .QN(n30516) );
  SDFFX1 \mem2_reg[153][19]  ( .D(n11639), .SI(\mem2[153][18] ), .SE(test_se), 
        .CLK(n1950), .Q(\mem2[153][19] ), .QN(n30517) );
  SDFFX1 \mem2_reg[153][18]  ( .D(n11638), .SI(\mem2[153][17] ), .SE(test_se), 
        .CLK(n1950), .Q(\mem2[153][18] ), .QN(n30518) );
  SDFFX1 \mem2_reg[153][17]  ( .D(n11637), .SI(\mem2[153][16] ), .SE(test_se), 
        .CLK(n1951), .Q(\mem2[153][17] ), .QN(n30519) );
  SDFFX1 \mem2_reg[153][16]  ( .D(n11636), .SI(\mem2[152][23] ), .SE(test_se), 
        .CLK(n1951), .Q(\mem2[153][16] ), .QN(n30520) );
  SDFFX1 \mem2_reg[152][23]  ( .D(n11635), .SI(\mem2[152][22] ), .SE(test_se), 
        .CLK(n1951), .Q(\mem2[152][23] ), .QN(n30521) );
  SDFFX1 \mem2_reg[152][22]  ( .D(n11634), .SI(\mem2[152][21] ), .SE(test_se), 
        .CLK(n1951), .Q(\mem2[152][22] ), .QN(n30522) );
  SDFFX1 \mem2_reg[152][21]  ( .D(n11633), .SI(\mem2[152][20] ), .SE(test_se), 
        .CLK(n1951), .Q(\mem2[152][21] ), .QN(n30523) );
  SDFFX1 \mem2_reg[152][20]  ( .D(n11632), .SI(\mem2[152][19] ), .SE(test_se), 
        .CLK(n1951), .Q(\mem2[152][20] ), .QN(n30524) );
  SDFFX1 \mem2_reg[152][19]  ( .D(n11631), .SI(\mem2[152][18] ), .SE(test_se), 
        .CLK(n1951), .Q(\mem2[152][19] ), .QN(n30525) );
  SDFFX1 \mem2_reg[152][18]  ( .D(n11630), .SI(\mem2[152][17] ), .SE(test_se), 
        .CLK(n1951), .Q(\mem2[152][18] ), .QN(n30526) );
  SDFFX1 \mem2_reg[152][17]  ( .D(n11629), .SI(\mem2[152][16] ), .SE(test_se), 
        .CLK(n1951), .Q(\mem2[152][17] ), .QN(n30527) );
  SDFFX1 \mem2_reg[152][16]  ( .D(n11628), .SI(\mem2[151][23] ), .SE(test_se), 
        .CLK(n1951), .Q(\mem2[152][16] ), .QN(n30528) );
  SDFFX1 \mem2_reg[151][23]  ( .D(n11627), .SI(\mem2[151][22] ), .SE(test_se), 
        .CLK(n1951), .Q(\mem2[151][23] ), .QN(n30529) );
  SDFFX1 \mem2_reg[151][22]  ( .D(n11626), .SI(\mem2[151][21] ), .SE(test_se), 
        .CLK(n1951), .Q(\mem2[151][22] ), .QN(n30530) );
  SDFFX1 \mem2_reg[151][21]  ( .D(n11625), .SI(\mem2[151][20] ), .SE(test_se), 
        .CLK(n1952), .Q(\mem2[151][21] ), .QN(n30531) );
  SDFFX1 \mem2_reg[151][20]  ( .D(n11624), .SI(\mem2[151][19] ), .SE(test_se), 
        .CLK(n1952), .Q(\mem2[151][20] ), .QN(n30532) );
  SDFFX1 \mem2_reg[151][19]  ( .D(n11623), .SI(\mem2[151][18] ), .SE(test_se), 
        .CLK(n1952), .Q(\mem2[151][19] ), .QN(n30533) );
  SDFFX1 \mem2_reg[151][18]  ( .D(n11622), .SI(\mem2[151][17] ), .SE(test_se), 
        .CLK(n1952), .Q(\mem2[151][18] ), .QN(n30534) );
  SDFFX1 \mem2_reg[151][17]  ( .D(n11621), .SI(\mem2[151][16] ), .SE(test_se), 
        .CLK(n1952), .Q(\mem2[151][17] ), .QN(n30535) );
  SDFFX1 \mem2_reg[151][16]  ( .D(n11620), .SI(\mem2[150][23] ), .SE(test_se), 
        .CLK(n1952), .Q(\mem2[151][16] ), .QN(n30536) );
  SDFFX1 \mem2_reg[150][23]  ( .D(n11619), .SI(\mem2[150][22] ), .SE(test_se), 
        .CLK(n1952), .Q(\mem2[150][23] ), .QN(n30537) );
  SDFFX1 \mem2_reg[150][22]  ( .D(n11618), .SI(\mem2[150][21] ), .SE(test_se), 
        .CLK(n1952), .Q(\mem2[150][22] ), .QN(n30538) );
  SDFFX1 \mem2_reg[150][21]  ( .D(n11617), .SI(\mem2[150][20] ), .SE(test_se), 
        .CLK(n1952), .Q(\mem2[150][21] ), .QN(n30539) );
  SDFFX1 \mem2_reg[150][20]  ( .D(n11616), .SI(\mem2[150][19] ), .SE(test_se), 
        .CLK(n1952), .Q(\mem2[150][20] ), .QN(n30540) );
  SDFFX1 \mem2_reg[150][19]  ( .D(n11615), .SI(\mem2[150][18] ), .SE(test_se), 
        .CLK(n1952), .Q(\mem2[150][19] ), .QN(n30541) );
  SDFFX1 \mem2_reg[150][18]  ( .D(n11614), .SI(\mem2[150][17] ), .SE(test_se), 
        .CLK(n1952), .Q(\mem2[150][18] ), .QN(n30542) );
  SDFFX1 \mem2_reg[150][17]  ( .D(n11613), .SI(\mem2[150][16] ), .SE(test_se), 
        .CLK(n1953), .Q(\mem2[150][17] ), .QN(n30543) );
  SDFFX1 \mem2_reg[150][16]  ( .D(n11612), .SI(\mem2[149][23] ), .SE(test_se), 
        .CLK(n1953), .Q(\mem2[150][16] ), .QN(n30544) );
  SDFFX1 \mem2_reg[149][23]  ( .D(n11611), .SI(\mem2[149][22] ), .SE(test_se), 
        .CLK(n1953), .Q(\mem2[149][23] ), .QN(n30545) );
  SDFFX1 \mem2_reg[149][22]  ( .D(n11610), .SI(\mem2[149][21] ), .SE(test_se), 
        .CLK(n1953), .Q(\mem2[149][22] ), .QN(n30546) );
  SDFFX1 \mem2_reg[149][21]  ( .D(n11609), .SI(\mem2[149][20] ), .SE(test_se), 
        .CLK(n1953), .Q(\mem2[149][21] ), .QN(n30547) );
  SDFFX1 \mem2_reg[149][20]  ( .D(n11608), .SI(\mem2[149][19] ), .SE(test_se), 
        .CLK(n1953), .Q(\mem2[149][20] ), .QN(n30548) );
  SDFFX1 \mem2_reg[149][19]  ( .D(n11607), .SI(\mem2[149][18] ), .SE(test_se), 
        .CLK(n1953), .Q(\mem2[149][19] ), .QN(n30549) );
  SDFFX1 \mem2_reg[149][18]  ( .D(n11606), .SI(\mem2[149][17] ), .SE(test_se), 
        .CLK(n1953), .Q(\mem2[149][18] ), .QN(n30550) );
  SDFFX1 \mem2_reg[149][17]  ( .D(n11605), .SI(\mem2[149][16] ), .SE(test_se), 
        .CLK(n1953), .Q(\mem2[149][17] ), .QN(n30551) );
  SDFFX1 \mem2_reg[149][16]  ( .D(n11604), .SI(\mem2[148][23] ), .SE(test_se), 
        .CLK(n1953), .Q(\mem2[149][16] ), .QN(n30552) );
  SDFFX1 \mem2_reg[148][23]  ( .D(n11603), .SI(\mem2[148][22] ), .SE(test_se), 
        .CLK(n1953), .Q(\mem2[148][23] ), .QN(n30553) );
  SDFFX1 \mem2_reg[148][22]  ( .D(n11602), .SI(\mem2[148][21] ), .SE(test_se), 
        .CLK(n1953), .Q(\mem2[148][22] ), .QN(n30554) );
  SDFFX1 \mem2_reg[148][21]  ( .D(n11601), .SI(\mem2[148][20] ), .SE(test_se), 
        .CLK(n1954), .Q(\mem2[148][21] ), .QN(n30555) );
  SDFFX1 \mem2_reg[148][20]  ( .D(n11600), .SI(\mem2[148][19] ), .SE(test_se), 
        .CLK(n1954), .Q(\mem2[148][20] ), .QN(n30556) );
  SDFFX1 \mem2_reg[148][19]  ( .D(n11599), .SI(\mem2[148][18] ), .SE(test_se), 
        .CLK(n1954), .Q(\mem2[148][19] ), .QN(n30557) );
  SDFFX1 \mem2_reg[148][18]  ( .D(n11598), .SI(\mem2[148][17] ), .SE(test_se), 
        .CLK(n1954), .Q(\mem2[148][18] ), .QN(n30558) );
  SDFFX1 \mem2_reg[148][17]  ( .D(n11597), .SI(\mem2[148][16] ), .SE(test_se), 
        .CLK(n1954), .Q(\mem2[148][17] ), .QN(n30559) );
  SDFFX1 \mem2_reg[148][16]  ( .D(n11596), .SI(\mem2[147][23] ), .SE(test_se), 
        .CLK(n1954), .Q(\mem2[148][16] ), .QN(n30560) );
  SDFFX1 \mem2_reg[147][23]  ( .D(n11595), .SI(\mem2[147][22] ), .SE(test_se), 
        .CLK(n1954), .Q(\mem2[147][23] ), .QN(n30561) );
  SDFFX1 \mem2_reg[147][22]  ( .D(n11594), .SI(\mem2[147][21] ), .SE(test_se), 
        .CLK(n1954), .Q(\mem2[147][22] ), .QN(n30562) );
  SDFFX1 \mem2_reg[147][21]  ( .D(n11593), .SI(\mem2[147][20] ), .SE(test_se), 
        .CLK(n1954), .Q(\mem2[147][21] ), .QN(n30563) );
  SDFFX1 \mem2_reg[147][20]  ( .D(n11592), .SI(\mem2[147][19] ), .SE(test_se), 
        .CLK(n1954), .Q(\mem2[147][20] ), .QN(n30564) );
  SDFFX1 \mem2_reg[147][19]  ( .D(n11591), .SI(\mem2[147][18] ), .SE(test_se), 
        .CLK(n1954), .Q(\mem2[147][19] ), .QN(n30565) );
  SDFFX1 \mem2_reg[147][18]  ( .D(n11590), .SI(\mem2[147][17] ), .SE(test_se), 
        .CLK(n1954), .Q(\mem2[147][18] ), .QN(n30566) );
  SDFFX1 \mem2_reg[147][17]  ( .D(n11589), .SI(\mem2[147][16] ), .SE(test_se), 
        .CLK(n1955), .Q(\mem2[147][17] ), .QN(n30567) );
  SDFFX1 \mem2_reg[147][16]  ( .D(n11588), .SI(\mem2[146][23] ), .SE(test_se), 
        .CLK(n1955), .Q(\mem2[147][16] ), .QN(n30568) );
  SDFFX1 \mem2_reg[146][23]  ( .D(n11587), .SI(\mem2[146][22] ), .SE(test_se), 
        .CLK(n1955), .Q(\mem2[146][23] ), .QN(n30569) );
  SDFFX1 \mem2_reg[146][22]  ( .D(n11586), .SI(\mem2[146][21] ), .SE(test_se), 
        .CLK(n1955), .Q(\mem2[146][22] ), .QN(n30570) );
  SDFFX1 \mem2_reg[146][21]  ( .D(n11585), .SI(\mem2[146][20] ), .SE(test_se), 
        .CLK(n1955), .Q(\mem2[146][21] ), .QN(n30571) );
  SDFFX1 \mem2_reg[146][20]  ( .D(n11584), .SI(\mem2[146][19] ), .SE(test_se), 
        .CLK(n1955), .Q(\mem2[146][20] ), .QN(n30572) );
  SDFFX1 \mem2_reg[146][19]  ( .D(n11583), .SI(\mem2[146][18] ), .SE(test_se), 
        .CLK(n1955), .Q(\mem2[146][19] ), .QN(n30573) );
  SDFFX1 \mem2_reg[146][18]  ( .D(n11582), .SI(\mem2[146][17] ), .SE(test_se), 
        .CLK(n1955), .Q(\mem2[146][18] ), .QN(n30574) );
  SDFFX1 \mem2_reg[146][17]  ( .D(n11581), .SI(\mem2[146][16] ), .SE(test_se), 
        .CLK(n1955), .Q(\mem2[146][17] ), .QN(n30575) );
  SDFFX1 \mem2_reg[146][16]  ( .D(n11580), .SI(\mem2[145][23] ), .SE(test_se), 
        .CLK(n1955), .Q(\mem2[146][16] ), .QN(n30576) );
  SDFFX1 \mem2_reg[145][23]  ( .D(n11579), .SI(\mem2[145][22] ), .SE(test_se), 
        .CLK(n1955), .Q(\mem2[145][23] ), .QN(n30577) );
  SDFFX1 \mem2_reg[145][22]  ( .D(n11578), .SI(\mem2[145][21] ), .SE(test_se), 
        .CLK(n1955), .Q(\mem2[145][22] ), .QN(n30578) );
  SDFFX1 \mem2_reg[145][21]  ( .D(n11577), .SI(\mem2[145][20] ), .SE(test_se), 
        .CLK(n1956), .Q(\mem2[145][21] ), .QN(n30579) );
  SDFFX1 \mem2_reg[145][20]  ( .D(n11576), .SI(\mem2[145][19] ), .SE(test_se), 
        .CLK(n1956), .Q(\mem2[145][20] ), .QN(n30580) );
  SDFFX1 \mem2_reg[145][19]  ( .D(n11575), .SI(\mem2[145][18] ), .SE(test_se), 
        .CLK(n1956), .Q(\mem2[145][19] ), .QN(n30581) );
  SDFFX1 \mem2_reg[145][18]  ( .D(n11574), .SI(\mem2[145][17] ), .SE(test_se), 
        .CLK(n1956), .Q(\mem2[145][18] ), .QN(n30582) );
  SDFFX1 \mem2_reg[145][17]  ( .D(n11573), .SI(\mem2[145][16] ), .SE(test_se), 
        .CLK(n1956), .Q(\mem2[145][17] ), .QN(n30583) );
  SDFFX1 \mem2_reg[145][16]  ( .D(n11572), .SI(\mem2[144][23] ), .SE(test_se), 
        .CLK(n1956), .Q(\mem2[145][16] ), .QN(n30584) );
  SDFFX1 \mem2_reg[144][23]  ( .D(n11571), .SI(\mem2[144][22] ), .SE(test_se), 
        .CLK(n1956), .Q(\mem2[144][23] ), .QN(n30585) );
  SDFFX1 \mem2_reg[144][22]  ( .D(n11570), .SI(\mem2[144][21] ), .SE(test_se), 
        .CLK(n1956), .Q(\mem2[144][22] ), .QN(n30586) );
  SDFFX1 \mem2_reg[144][21]  ( .D(n11569), .SI(\mem2[144][20] ), .SE(test_se), 
        .CLK(n1956), .Q(\mem2[144][21] ), .QN(n30587) );
  SDFFX1 \mem2_reg[144][20]  ( .D(n11568), .SI(\mem2[144][19] ), .SE(test_se), 
        .CLK(n1956), .Q(\mem2[144][20] ), .QN(n30588) );
  SDFFX1 \mem2_reg[144][19]  ( .D(n11567), .SI(\mem2[144][18] ), .SE(test_se), 
        .CLK(n1956), .Q(\mem2[144][19] ), .QN(n30589) );
  SDFFX1 \mem2_reg[144][18]  ( .D(n11566), .SI(\mem2[144][17] ), .SE(test_se), 
        .CLK(n1956), .Q(\mem2[144][18] ), .QN(n30590) );
  SDFFX1 \mem2_reg[144][17]  ( .D(n11565), .SI(\mem2[144][16] ), .SE(test_se), 
        .CLK(n1957), .Q(\mem2[144][17] ), .QN(n30591) );
  SDFFX1 \mem2_reg[144][16]  ( .D(n11564), .SI(\mem2[143][23] ), .SE(test_se), 
        .CLK(n1957), .Q(\mem2[144][16] ), .QN(n30592) );
  SDFFX1 \mem2_reg[143][23]  ( .D(n11563), .SI(\mem2[143][22] ), .SE(test_se), 
        .CLK(n1957), .Q(\mem2[143][23] ), .QN(n30593) );
  SDFFX1 \mem2_reg[143][22]  ( .D(n11562), .SI(\mem2[143][21] ), .SE(test_se), 
        .CLK(n1957), .Q(\mem2[143][22] ), .QN(n30594) );
  SDFFX1 \mem2_reg[143][21]  ( .D(n11561), .SI(\mem2[143][20] ), .SE(test_se), 
        .CLK(n1957), .Q(\mem2[143][21] ), .QN(n30595) );
  SDFFX1 \mem2_reg[143][20]  ( .D(n11560), .SI(\mem2[143][19] ), .SE(test_se), 
        .CLK(n1957), .Q(\mem2[143][20] ), .QN(n30596) );
  SDFFX1 \mem2_reg[143][19]  ( .D(n11559), .SI(\mem2[143][18] ), .SE(test_se), 
        .CLK(n1957), .Q(\mem2[143][19] ), .QN(n30597) );
  SDFFX1 \mem2_reg[143][18]  ( .D(n11558), .SI(\mem2[143][17] ), .SE(test_se), 
        .CLK(n1957), .Q(\mem2[143][18] ), .QN(n30598) );
  SDFFX1 \mem2_reg[143][17]  ( .D(n11557), .SI(\mem2[143][16] ), .SE(test_se), 
        .CLK(n1957), .Q(\mem2[143][17] ), .QN(n30599) );
  SDFFX1 \mem2_reg[143][16]  ( .D(n11556), .SI(\mem2[142][23] ), .SE(test_se), 
        .CLK(n1957), .Q(\mem2[143][16] ), .QN(n30600) );
  SDFFX1 \mem2_reg[142][23]  ( .D(n11555), .SI(\mem2[142][22] ), .SE(test_se), 
        .CLK(n1957), .Q(\mem2[142][23] ), .QN(n30601) );
  SDFFX1 \mem2_reg[142][22]  ( .D(n11554), .SI(\mem2[142][21] ), .SE(test_se), 
        .CLK(n1957), .Q(\mem2[142][22] ), .QN(n30602) );
  SDFFX1 \mem2_reg[142][21]  ( .D(n11553), .SI(\mem2[142][20] ), .SE(test_se), 
        .CLK(n1958), .Q(\mem2[142][21] ), .QN(n30603) );
  SDFFX1 \mem2_reg[142][20]  ( .D(n11552), .SI(\mem2[142][19] ), .SE(test_se), 
        .CLK(n1958), .Q(\mem2[142][20] ), .QN(n30604) );
  SDFFX1 \mem2_reg[142][19]  ( .D(n11551), .SI(\mem2[142][18] ), .SE(test_se), 
        .CLK(n1958), .Q(\mem2[142][19] ), .QN(n30605) );
  SDFFX1 \mem2_reg[142][18]  ( .D(n11550), .SI(\mem2[142][17] ), .SE(test_se), 
        .CLK(n1958), .Q(\mem2[142][18] ), .QN(n30606) );
  SDFFX1 \mem2_reg[142][17]  ( .D(n11549), .SI(\mem2[142][16] ), .SE(test_se), 
        .CLK(n1958), .Q(\mem2[142][17] ), .QN(n30607) );
  SDFFX1 \mem2_reg[142][16]  ( .D(n11548), .SI(\mem2[141][23] ), .SE(test_se), 
        .CLK(n1958), .Q(\mem2[142][16] ), .QN(n30608) );
  SDFFX1 \mem2_reg[141][23]  ( .D(n11547), .SI(\mem2[141][22] ), .SE(test_se), 
        .CLK(n1958), .Q(\mem2[141][23] ), .QN(n30609) );
  SDFFX1 \mem2_reg[141][22]  ( .D(n11546), .SI(\mem2[141][21] ), .SE(test_se), 
        .CLK(n1958), .Q(\mem2[141][22] ), .QN(n30610) );
  SDFFX1 \mem2_reg[141][21]  ( .D(n11545), .SI(\mem2[141][20] ), .SE(test_se), 
        .CLK(n1958), .Q(\mem2[141][21] ), .QN(n30611) );
  SDFFX1 \mem2_reg[141][20]  ( .D(n11544), .SI(\mem2[141][19] ), .SE(test_se), 
        .CLK(n1958), .Q(\mem2[141][20] ), .QN(n30612) );
  SDFFX1 \mem2_reg[141][19]  ( .D(n11543), .SI(\mem2[141][18] ), .SE(test_se), 
        .CLK(n1958), .Q(\mem2[141][19] ), .QN(n30613) );
  SDFFX1 \mem2_reg[141][18]  ( .D(n11542), .SI(\mem2[141][17] ), .SE(test_se), 
        .CLK(n1958), .Q(\mem2[141][18] ), .QN(n30614) );
  SDFFX1 \mem2_reg[141][17]  ( .D(n11541), .SI(\mem2[141][16] ), .SE(test_se), 
        .CLK(n1959), .Q(\mem2[141][17] ), .QN(n30615) );
  SDFFX1 \mem2_reg[141][16]  ( .D(n11540), .SI(\mem2[140][23] ), .SE(test_se), 
        .CLK(n1959), .Q(\mem2[141][16] ), .QN(n30616) );
  SDFFX1 \mem2_reg[140][23]  ( .D(n11539), .SI(\mem2[140][22] ), .SE(test_se), 
        .CLK(n1959), .Q(\mem2[140][23] ), .QN(n30617) );
  SDFFX1 \mem2_reg[140][22]  ( .D(n11538), .SI(\mem2[140][21] ), .SE(test_se), 
        .CLK(n1959), .Q(\mem2[140][22] ), .QN(n30618) );
  SDFFX1 \mem2_reg[140][21]  ( .D(n11537), .SI(\mem2[140][20] ), .SE(test_se), 
        .CLK(n1959), .Q(\mem2[140][21] ), .QN(n30619) );
  SDFFX1 \mem2_reg[140][20]  ( .D(n11536), .SI(\mem2[140][19] ), .SE(test_se), 
        .CLK(n1959), .Q(\mem2[140][20] ), .QN(n30620) );
  SDFFX1 \mem2_reg[140][19]  ( .D(n11535), .SI(\mem2[140][18] ), .SE(test_se), 
        .CLK(n1959), .Q(\mem2[140][19] ), .QN(n30621) );
  SDFFX1 \mem2_reg[140][18]  ( .D(n11534), .SI(\mem2[140][17] ), .SE(test_se), 
        .CLK(n1959), .Q(\mem2[140][18] ), .QN(n30622) );
  SDFFX1 \mem2_reg[140][17]  ( .D(n11533), .SI(\mem2[140][16] ), .SE(test_se), 
        .CLK(n1959), .Q(\mem2[140][17] ), .QN(n30623) );
  SDFFX1 \mem2_reg[140][16]  ( .D(n11532), .SI(\mem2[139][23] ), .SE(test_se), 
        .CLK(n1959), .Q(\mem2[140][16] ), .QN(n30624) );
  SDFFX1 \mem2_reg[139][23]  ( .D(n11531), .SI(\mem2[139][22] ), .SE(test_se), 
        .CLK(n1959), .Q(\mem2[139][23] ), .QN(n30625) );
  SDFFX1 \mem2_reg[139][22]  ( .D(n11530), .SI(\mem2[139][21] ), .SE(test_se), 
        .CLK(n1959), .Q(\mem2[139][22] ), .QN(n30626) );
  SDFFX1 \mem2_reg[139][21]  ( .D(n11529), .SI(\mem2[139][20] ), .SE(test_se), 
        .CLK(n1960), .Q(\mem2[139][21] ), .QN(n30627) );
  SDFFX1 \mem2_reg[139][20]  ( .D(n11528), .SI(\mem2[139][19] ), .SE(test_se), 
        .CLK(n1960), .Q(\mem2[139][20] ), .QN(n30628) );
  SDFFX1 \mem2_reg[139][19]  ( .D(n11527), .SI(\mem2[139][18] ), .SE(test_se), 
        .CLK(n1960), .Q(\mem2[139][19] ), .QN(n30629) );
  SDFFX1 \mem2_reg[139][18]  ( .D(n11526), .SI(\mem2[139][17] ), .SE(test_se), 
        .CLK(n1960), .Q(\mem2[139][18] ), .QN(n30630) );
  SDFFX1 \mem2_reg[139][17]  ( .D(n11525), .SI(\mem2[139][16] ), .SE(test_se), 
        .CLK(n1960), .Q(\mem2[139][17] ), .QN(n30631) );
  SDFFX1 \mem2_reg[139][16]  ( .D(n11524), .SI(\mem2[138][23] ), .SE(test_se), 
        .CLK(n1960), .Q(\mem2[139][16] ), .QN(n30632) );
  SDFFX1 \mem2_reg[138][23]  ( .D(n11523), .SI(\mem2[138][22] ), .SE(test_se), 
        .CLK(n1960), .Q(\mem2[138][23] ), .QN(n30633) );
  SDFFX1 \mem2_reg[138][22]  ( .D(n11522), .SI(\mem2[138][21] ), .SE(test_se), 
        .CLK(n1960), .Q(\mem2[138][22] ), .QN(n30634) );
  SDFFX1 \mem2_reg[138][21]  ( .D(n11521), .SI(\mem2[138][20] ), .SE(test_se), 
        .CLK(n1960), .Q(\mem2[138][21] ), .QN(n30635) );
  SDFFX1 \mem2_reg[138][20]  ( .D(n11520), .SI(\mem2[138][19] ), .SE(test_se), 
        .CLK(n1960), .Q(\mem2[138][20] ), .QN(n30636) );
  SDFFX1 \mem2_reg[138][19]  ( .D(n11519), .SI(\mem2[138][18] ), .SE(test_se), 
        .CLK(n1960), .Q(\mem2[138][19] ), .QN(n30637) );
  SDFFX1 \mem2_reg[138][18]  ( .D(n11518), .SI(\mem2[138][17] ), .SE(test_se), 
        .CLK(n1960), .Q(\mem2[138][18] ), .QN(n30638) );
  SDFFX1 \mem2_reg[138][17]  ( .D(n11517), .SI(\mem2[138][16] ), .SE(test_se), 
        .CLK(n1961), .Q(\mem2[138][17] ), .QN(n30639) );
  SDFFX1 \mem2_reg[138][16]  ( .D(n11516), .SI(\mem2[137][23] ), .SE(test_se), 
        .CLK(n1961), .Q(\mem2[138][16] ), .QN(n30640) );
  SDFFX1 \mem2_reg[137][23]  ( .D(n11515), .SI(\mem2[137][22] ), .SE(test_se), 
        .CLK(n1961), .Q(\mem2[137][23] ), .QN(n30641) );
  SDFFX1 \mem2_reg[137][22]  ( .D(n11514), .SI(\mem2[137][21] ), .SE(test_se), 
        .CLK(n1961), .Q(\mem2[137][22] ), .QN(n30642) );
  SDFFX1 \mem2_reg[137][21]  ( .D(n11513), .SI(\mem2[137][20] ), .SE(test_se), 
        .CLK(n1961), .Q(\mem2[137][21] ), .QN(n30643) );
  SDFFX1 \mem2_reg[137][20]  ( .D(n11512), .SI(\mem2[137][19] ), .SE(test_se), 
        .CLK(n1961), .Q(\mem2[137][20] ), .QN(n30644) );
  SDFFX1 \mem2_reg[137][19]  ( .D(n11511), .SI(\mem2[137][18] ), .SE(test_se), 
        .CLK(n1961), .Q(\mem2[137][19] ), .QN(n30645) );
  SDFFX1 \mem2_reg[137][18]  ( .D(n11510), .SI(\mem2[137][17] ), .SE(test_se), 
        .CLK(n1961), .Q(\mem2[137][18] ), .QN(n30646) );
  SDFFX1 \mem2_reg[137][17]  ( .D(n11509), .SI(\mem2[137][16] ), .SE(test_se), 
        .CLK(n1961), .Q(\mem2[137][17] ), .QN(n30647) );
  SDFFX1 \mem2_reg[137][16]  ( .D(n11508), .SI(\mem2[136][23] ), .SE(test_se), 
        .CLK(n1961), .Q(\mem2[137][16] ), .QN(n30648) );
  SDFFX1 \mem2_reg[136][23]  ( .D(n11507), .SI(\mem2[136][22] ), .SE(test_se), 
        .CLK(n1961), .Q(\mem2[136][23] ), .QN(n30649) );
  SDFFX1 \mem2_reg[136][22]  ( .D(n11506), .SI(\mem2[136][21] ), .SE(test_se), 
        .CLK(n1961), .Q(\mem2[136][22] ), .QN(n30650) );
  SDFFX1 \mem2_reg[136][21]  ( .D(n11505), .SI(\mem2[136][20] ), .SE(test_se), 
        .CLK(n1962), .Q(\mem2[136][21] ), .QN(n30651) );
  SDFFX1 \mem2_reg[136][20]  ( .D(n11504), .SI(\mem2[136][19] ), .SE(test_se), 
        .CLK(n1962), .Q(\mem2[136][20] ), .QN(n30652) );
  SDFFX1 \mem2_reg[136][19]  ( .D(n11503), .SI(\mem2[136][18] ), .SE(test_se), 
        .CLK(n1962), .Q(\mem2[136][19] ), .QN(n30653) );
  SDFFX1 \mem2_reg[136][18]  ( .D(n11502), .SI(\mem2[136][17] ), .SE(test_se), 
        .CLK(n1962), .Q(\mem2[136][18] ), .QN(n30654) );
  SDFFX1 \mem2_reg[136][17]  ( .D(n11501), .SI(\mem2[136][16] ), .SE(test_se), 
        .CLK(n1962), .Q(\mem2[136][17] ), .QN(n30655) );
  SDFFX1 \mem2_reg[136][16]  ( .D(n11500), .SI(\mem2[135][23] ), .SE(test_se), 
        .CLK(n1962), .Q(\mem2[136][16] ), .QN(n30656) );
  SDFFX1 \mem2_reg[135][23]  ( .D(n11499), .SI(\mem2[135][22] ), .SE(test_se), 
        .CLK(n1962), .Q(\mem2[135][23] ), .QN(n30657) );
  SDFFX1 \mem2_reg[135][22]  ( .D(n11498), .SI(\mem2[135][21] ), .SE(test_se), 
        .CLK(n1962), .Q(\mem2[135][22] ), .QN(n30658) );
  SDFFX1 \mem2_reg[135][21]  ( .D(n11497), .SI(\mem2[135][20] ), .SE(test_se), 
        .CLK(n1962), .Q(\mem2[135][21] ), .QN(n30659) );
  SDFFX1 \mem2_reg[135][20]  ( .D(n11496), .SI(\mem2[135][19] ), .SE(test_se), 
        .CLK(n1962), .Q(\mem2[135][20] ), .QN(n30660) );
  SDFFX1 \mem2_reg[135][19]  ( .D(n11495), .SI(\mem2[135][18] ), .SE(test_se), 
        .CLK(n1962), .Q(\mem2[135][19] ), .QN(n30661) );
  SDFFX1 \mem2_reg[135][18]  ( .D(n11494), .SI(\mem2[135][17] ), .SE(test_se), 
        .CLK(n1962), .Q(\mem2[135][18] ), .QN(n30662) );
  SDFFX1 \mem2_reg[135][17]  ( .D(n11493), .SI(\mem2[135][16] ), .SE(test_se), 
        .CLK(n1963), .Q(\mem2[135][17] ), .QN(n30663) );
  SDFFX1 \mem2_reg[135][16]  ( .D(n11492), .SI(\mem2[134][23] ), .SE(test_se), 
        .CLK(n1963), .Q(\mem2[135][16] ), .QN(n30664) );
  SDFFX1 \mem2_reg[134][23]  ( .D(n11491), .SI(\mem2[134][22] ), .SE(test_se), 
        .CLK(n1963), .Q(\mem2[134][23] ), .QN(n30665) );
  SDFFX1 \mem2_reg[134][22]  ( .D(n11490), .SI(\mem2[134][21] ), .SE(test_se), 
        .CLK(n1963), .Q(\mem2[134][22] ), .QN(n30666) );
  SDFFX1 \mem2_reg[134][21]  ( .D(n11489), .SI(\mem2[134][20] ), .SE(test_se), 
        .CLK(n1963), .Q(\mem2[134][21] ), .QN(n30667) );
  SDFFX1 \mem2_reg[134][20]  ( .D(n11488), .SI(\mem2[134][19] ), .SE(test_se), 
        .CLK(n1963), .Q(\mem2[134][20] ), .QN(n30668) );
  SDFFX1 \mem2_reg[134][19]  ( .D(n11487), .SI(\mem2[134][18] ), .SE(test_se), 
        .CLK(n1963), .Q(\mem2[134][19] ), .QN(n30669) );
  SDFFX1 \mem2_reg[134][18]  ( .D(n11486), .SI(\mem2[134][17] ), .SE(test_se), 
        .CLK(n1963), .Q(\mem2[134][18] ), .QN(n30670) );
  SDFFX1 \mem2_reg[134][17]  ( .D(n11485), .SI(\mem2[134][16] ), .SE(test_se), 
        .CLK(n1963), .Q(\mem2[134][17] ), .QN(n30671) );
  SDFFX1 \mem2_reg[134][16]  ( .D(n11484), .SI(\mem2[133][23] ), .SE(test_se), 
        .CLK(n1963), .Q(\mem2[134][16] ), .QN(n30672) );
  SDFFX1 \mem2_reg[133][23]  ( .D(n11483), .SI(\mem2[133][22] ), .SE(test_se), 
        .CLK(n1963), .Q(\mem2[133][23] ), .QN(n30673) );
  SDFFX1 \mem2_reg[133][22]  ( .D(n11482), .SI(\mem2[133][21] ), .SE(test_se), 
        .CLK(n1963), .Q(\mem2[133][22] ), .QN(n30674) );
  SDFFX1 \mem2_reg[133][21]  ( .D(n11481), .SI(\mem2[133][20] ), .SE(test_se), 
        .CLK(n1964), .Q(\mem2[133][21] ), .QN(n30675) );
  SDFFX1 \mem2_reg[133][20]  ( .D(n11480), .SI(\mem2[133][19] ), .SE(test_se), 
        .CLK(n1964), .Q(\mem2[133][20] ), .QN(n30676) );
  SDFFX1 \mem2_reg[133][19]  ( .D(n11479), .SI(\mem2[133][18] ), .SE(test_se), 
        .CLK(n1964), .Q(\mem2[133][19] ), .QN(n30677) );
  SDFFX1 \mem2_reg[133][18]  ( .D(n11478), .SI(\mem2[133][17] ), .SE(test_se), 
        .CLK(n1964), .Q(\mem2[133][18] ), .QN(n30678) );
  SDFFX1 \mem2_reg[133][17]  ( .D(n11477), .SI(\mem2[133][16] ), .SE(test_se), 
        .CLK(n1964), .Q(\mem2[133][17] ), .QN(n30679) );
  SDFFX1 \mem2_reg[133][16]  ( .D(n11476), .SI(\mem2[132][23] ), .SE(test_se), 
        .CLK(n1964), .Q(\mem2[133][16] ), .QN(n30680) );
  SDFFX1 \mem2_reg[132][23]  ( .D(n11475), .SI(\mem2[132][22] ), .SE(test_se), 
        .CLK(n1964), .Q(\mem2[132][23] ), .QN(n30681) );
  SDFFX1 \mem2_reg[132][22]  ( .D(n11474), .SI(\mem2[132][21] ), .SE(test_se), 
        .CLK(n1964), .Q(\mem2[132][22] ), .QN(n30682) );
  SDFFX1 \mem2_reg[132][21]  ( .D(n11473), .SI(\mem2[132][20] ), .SE(test_se), 
        .CLK(n1964), .Q(\mem2[132][21] ), .QN(n30683) );
  SDFFX1 \mem2_reg[132][20]  ( .D(n11472), .SI(\mem2[132][19] ), .SE(test_se), 
        .CLK(n1964), .Q(\mem2[132][20] ), .QN(n30684) );
  SDFFX1 \mem2_reg[132][19]  ( .D(n11471), .SI(\mem2[132][18] ), .SE(test_se), 
        .CLK(n1964), .Q(\mem2[132][19] ), .QN(n30685) );
  SDFFX1 \mem2_reg[132][18]  ( .D(n11470), .SI(\mem2[132][17] ), .SE(test_se), 
        .CLK(n1964), .Q(\mem2[132][18] ), .QN(n30686) );
  SDFFX1 \mem2_reg[132][17]  ( .D(n11469), .SI(\mem2[132][16] ), .SE(test_se), 
        .CLK(n1965), .Q(\mem2[132][17] ), .QN(n30687) );
  SDFFX1 \mem2_reg[132][16]  ( .D(n11468), .SI(\mem2[131][23] ), .SE(test_se), 
        .CLK(n1965), .Q(\mem2[132][16] ), .QN(n30688) );
  SDFFX1 \mem2_reg[131][23]  ( .D(n11467), .SI(\mem2[131][22] ), .SE(test_se), 
        .CLK(n1965), .Q(\mem2[131][23] ), .QN(n30689) );
  SDFFX1 \mem2_reg[131][22]  ( .D(n11466), .SI(\mem2[131][21] ), .SE(test_se), 
        .CLK(n1965), .Q(\mem2[131][22] ), .QN(n30690) );
  SDFFX1 \mem2_reg[131][21]  ( .D(n11465), .SI(\mem2[131][20] ), .SE(test_se), 
        .CLK(n1965), .Q(\mem2[131][21] ), .QN(n30691) );
  SDFFX1 \mem2_reg[131][20]  ( .D(n11464), .SI(\mem2[131][19] ), .SE(test_se), 
        .CLK(n1965), .Q(\mem2[131][20] ), .QN(n30692) );
  SDFFX1 \mem2_reg[131][19]  ( .D(n11463), .SI(\mem2[131][18] ), .SE(test_se), 
        .CLK(n1965), .Q(\mem2[131][19] ), .QN(n30693) );
  SDFFX1 \mem2_reg[131][18]  ( .D(n11462), .SI(\mem2[131][17] ), .SE(test_se), 
        .CLK(n1965), .Q(\mem2[131][18] ), .QN(n30694) );
  SDFFX1 \mem2_reg[131][17]  ( .D(n11461), .SI(\mem2[131][16] ), .SE(test_se), 
        .CLK(n1965), .Q(\mem2[131][17] ), .QN(n30695) );
  SDFFX1 \mem2_reg[131][16]  ( .D(n11460), .SI(\mem2[130][23] ), .SE(test_se), 
        .CLK(n1965), .Q(\mem2[131][16] ), .QN(n30696) );
  SDFFX1 \mem2_reg[130][23]  ( .D(n11459), .SI(\mem2[130][22] ), .SE(test_se), 
        .CLK(n1965), .Q(\mem2[130][23] ), .QN(n30697) );
  SDFFX1 \mem2_reg[130][22]  ( .D(n11458), .SI(\mem2[130][21] ), .SE(test_se), 
        .CLK(n1965), .Q(\mem2[130][22] ), .QN(n30698) );
  SDFFX1 \mem2_reg[130][21]  ( .D(n11457), .SI(\mem2[130][20] ), .SE(test_se), 
        .CLK(n1966), .Q(\mem2[130][21] ), .QN(n30699) );
  SDFFX1 \mem2_reg[130][20]  ( .D(n11456), .SI(\mem2[130][19] ), .SE(test_se), 
        .CLK(n1966), .Q(\mem2[130][20] ), .QN(n30700) );
  SDFFX1 \mem2_reg[130][19]  ( .D(n11455), .SI(\mem2[130][18] ), .SE(test_se), 
        .CLK(n1966), .Q(\mem2[130][19] ), .QN(n30701) );
  SDFFX1 \mem2_reg[130][18]  ( .D(n11454), .SI(\mem2[130][17] ), .SE(test_se), 
        .CLK(n1966), .Q(\mem2[130][18] ), .QN(n30702) );
  SDFFX1 \mem2_reg[130][17]  ( .D(n11453), .SI(\mem2[130][16] ), .SE(test_se), 
        .CLK(n1966), .Q(\mem2[130][17] ), .QN(n30703) );
  SDFFX1 \mem2_reg[130][16]  ( .D(n11452), .SI(\mem2[129][23] ), .SE(test_se), 
        .CLK(n1966), .Q(\mem2[130][16] ), .QN(n30704) );
  SDFFX1 \mem2_reg[129][23]  ( .D(n11451), .SI(\mem2[129][22] ), .SE(test_se), 
        .CLK(n1966), .Q(\mem2[129][23] ), .QN(n30705) );
  SDFFX1 \mem2_reg[129][22]  ( .D(n11450), .SI(\mem2[129][21] ), .SE(test_se), 
        .CLK(n1966), .Q(\mem2[129][22] ), .QN(n30706) );
  SDFFX1 \mem2_reg[129][21]  ( .D(n11449), .SI(\mem2[129][20] ), .SE(test_se), 
        .CLK(n1966), .Q(\mem2[129][21] ), .QN(n30707) );
  SDFFX1 \mem2_reg[129][20]  ( .D(n11448), .SI(\mem2[129][19] ), .SE(test_se), 
        .CLK(n1966), .Q(\mem2[129][20] ), .QN(n30708) );
  SDFFX1 \mem2_reg[129][19]  ( .D(n11447), .SI(\mem2[129][18] ), .SE(test_se), 
        .CLK(n1966), .Q(\mem2[129][19] ), .QN(n30709) );
  SDFFX1 \mem2_reg[129][18]  ( .D(n11446), .SI(\mem2[129][17] ), .SE(test_se), 
        .CLK(n1966), .Q(\mem2[129][18] ), .QN(n30710) );
  SDFFX1 \mem2_reg[129][17]  ( .D(n11445), .SI(\mem2[129][16] ), .SE(test_se), 
        .CLK(n1967), .Q(\mem2[129][17] ), .QN(n30711) );
  SDFFX1 \mem2_reg[129][16]  ( .D(n11444), .SI(\mem2[128][23] ), .SE(test_se), 
        .CLK(n1967), .Q(\mem2[129][16] ), .QN(n30712) );
  SDFFX1 \mem2_reg[128][23]  ( .D(n11443), .SI(\mem2[128][22] ), .SE(test_se), 
        .CLK(n1967), .Q(\mem2[128][23] ), .QN(n30713) );
  SDFFX1 \mem2_reg[128][22]  ( .D(n11442), .SI(\mem2[128][21] ), .SE(test_se), 
        .CLK(n1967), .Q(\mem2[128][22] ), .QN(n30714) );
  SDFFX1 \mem2_reg[128][21]  ( .D(n11441), .SI(\mem2[128][20] ), .SE(test_se), 
        .CLK(n1967), .Q(\mem2[128][21] ), .QN(n30715) );
  SDFFX1 \mem2_reg[128][20]  ( .D(n11440), .SI(\mem2[128][19] ), .SE(test_se), 
        .CLK(n1967), .Q(\mem2[128][20] ), .QN(n30716) );
  SDFFX1 \mem2_reg[128][19]  ( .D(n11439), .SI(\mem2[128][18] ), .SE(test_se), 
        .CLK(n1967), .Q(\mem2[128][19] ), .QN(n30717) );
  SDFFX1 \mem2_reg[128][18]  ( .D(n11438), .SI(\mem2[128][17] ), .SE(test_se), 
        .CLK(n1967), .Q(\mem2[128][18] ), .QN(n30718) );
  SDFFX1 \mem2_reg[128][17]  ( .D(n11437), .SI(\mem2[128][16] ), .SE(test_se), 
        .CLK(n1967), .Q(\mem2[128][17] ), .QN(n30719) );
  SDFFX1 \mem2_reg[128][16]  ( .D(n11436), .SI(\mem2[127][23] ), .SE(test_se), 
        .CLK(n1967), .Q(\mem2[128][16] ), .QN(n30720) );
  SDFFX1 \mem2_reg[127][23]  ( .D(n11435), .SI(\mem2[127][22] ), .SE(test_se), 
        .CLK(n1967), .Q(\mem2[127][23] ), .QN(n30721) );
  SDFFX1 \mem2_reg[127][22]  ( .D(n11434), .SI(\mem2[127][21] ), .SE(test_se), 
        .CLK(n1967), .Q(\mem2[127][22] ), .QN(n30722) );
  SDFFX1 \mem2_reg[127][21]  ( .D(n11433), .SI(\mem2[127][20] ), .SE(test_se), 
        .CLK(n1968), .Q(\mem2[127][21] ), .QN(n30723) );
  SDFFX1 \mem2_reg[127][20]  ( .D(n11432), .SI(\mem2[127][19] ), .SE(test_se), 
        .CLK(n1968), .Q(\mem2[127][20] ), .QN(n30724) );
  SDFFX1 \mem2_reg[127][19]  ( .D(n11431), .SI(\mem2[127][18] ), .SE(test_se), 
        .CLK(n1968), .Q(\mem2[127][19] ), .QN(n30725) );
  SDFFX1 \mem2_reg[127][18]  ( .D(n11430), .SI(\mem2[127][17] ), .SE(test_se), 
        .CLK(n1968), .Q(\mem2[127][18] ), .QN(n30726) );
  SDFFX1 \mem2_reg[127][17]  ( .D(n11429), .SI(\mem2[127][16] ), .SE(test_se), 
        .CLK(n1968), .Q(\mem2[127][17] ), .QN(n30727) );
  SDFFX1 \mem2_reg[127][16]  ( .D(n11428), .SI(\mem2[126][23] ), .SE(test_se), 
        .CLK(n1968), .Q(\mem2[127][16] ), .QN(n30728) );
  SDFFX1 \mem2_reg[126][23]  ( .D(n11427), .SI(\mem2[126][22] ), .SE(test_se), 
        .CLK(n1968), .Q(\mem2[126][23] ), .QN(n30729) );
  SDFFX1 \mem2_reg[126][22]  ( .D(n11426), .SI(\mem2[126][21] ), .SE(test_se), 
        .CLK(n1968), .Q(\mem2[126][22] ), .QN(n30730) );
  SDFFX1 \mem2_reg[126][21]  ( .D(n11425), .SI(\mem2[126][20] ), .SE(test_se), 
        .CLK(n1968), .Q(\mem2[126][21] ), .QN(n30731) );
  SDFFX1 \mem2_reg[126][20]  ( .D(n11424), .SI(\mem2[126][19] ), .SE(test_se), 
        .CLK(n1968), .Q(\mem2[126][20] ), .QN(n30732) );
  SDFFX1 \mem2_reg[126][19]  ( .D(n11423), .SI(\mem2[126][18] ), .SE(test_se), 
        .CLK(n1968), .Q(\mem2[126][19] ), .QN(n30733) );
  SDFFX1 \mem2_reg[126][18]  ( .D(n11422), .SI(\mem2[126][17] ), .SE(test_se), 
        .CLK(n1968), .Q(\mem2[126][18] ), .QN(n30734) );
  SDFFX1 \mem2_reg[126][17]  ( .D(n11421), .SI(\mem2[126][16] ), .SE(test_se), 
        .CLK(n1969), .Q(\mem2[126][17] ), .QN(n30735) );
  SDFFX1 \mem2_reg[126][16]  ( .D(n11420), .SI(\mem2[125][23] ), .SE(test_se), 
        .CLK(n1969), .Q(\mem2[126][16] ), .QN(n30736) );
  SDFFX1 \mem2_reg[125][23]  ( .D(n11419), .SI(\mem2[125][22] ), .SE(test_se), 
        .CLK(n1969), .Q(\mem2[125][23] ), .QN(n30737) );
  SDFFX1 \mem2_reg[125][22]  ( .D(n11418), .SI(\mem2[125][21] ), .SE(test_se), 
        .CLK(n1969), .Q(\mem2[125][22] ), .QN(n30738) );
  SDFFX1 \mem2_reg[125][21]  ( .D(n11417), .SI(\mem2[125][20] ), .SE(test_se), 
        .CLK(n1969), .Q(\mem2[125][21] ), .QN(n30739) );
  SDFFX1 \mem2_reg[125][20]  ( .D(n11416), .SI(\mem2[125][19] ), .SE(test_se), 
        .CLK(n1969), .Q(\mem2[125][20] ), .QN(n30740) );
  SDFFX1 \mem2_reg[125][19]  ( .D(n11415), .SI(\mem2[125][18] ), .SE(test_se), 
        .CLK(n1969), .Q(\mem2[125][19] ), .QN(n30741) );
  SDFFX1 \mem2_reg[125][18]  ( .D(n11414), .SI(\mem2[125][17] ), .SE(test_se), 
        .CLK(n1969), .Q(\mem2[125][18] ), .QN(n30742) );
  SDFFX1 \mem2_reg[125][17]  ( .D(n11413), .SI(\mem2[125][16] ), .SE(test_se), 
        .CLK(n1969), .Q(\mem2[125][17] ), .QN(n30743) );
  SDFFX1 \mem2_reg[125][16]  ( .D(n11412), .SI(\mem2[124][23] ), .SE(test_se), 
        .CLK(n1969), .Q(\mem2[125][16] ), .QN(n30744) );
  SDFFX1 \mem2_reg[124][23]  ( .D(n11411), .SI(\mem2[124][22] ), .SE(test_se), 
        .CLK(n1969), .Q(\mem2[124][23] ), .QN(n30745) );
  SDFFX1 \mem2_reg[124][22]  ( .D(n11410), .SI(\mem2[124][21] ), .SE(test_se), 
        .CLK(n1969), .Q(\mem2[124][22] ), .QN(n30746) );
  SDFFX1 \mem2_reg[124][21]  ( .D(n11409), .SI(\mem2[124][20] ), .SE(test_se), 
        .CLK(n1970), .Q(\mem2[124][21] ), .QN(n30747) );
  SDFFX1 \mem2_reg[124][20]  ( .D(n11408), .SI(\mem2[124][19] ), .SE(test_se), 
        .CLK(n1970), .Q(\mem2[124][20] ), .QN(n30748) );
  SDFFX1 \mem2_reg[124][19]  ( .D(n11407), .SI(\mem2[124][18] ), .SE(test_se), 
        .CLK(n1970), .Q(\mem2[124][19] ), .QN(n30749) );
  SDFFX1 \mem2_reg[124][18]  ( .D(n11406), .SI(\mem2[124][17] ), .SE(test_se), 
        .CLK(n1970), .Q(\mem2[124][18] ), .QN(n30750) );
  SDFFX1 \mem2_reg[124][17]  ( .D(n11405), .SI(\mem2[124][16] ), .SE(test_se), 
        .CLK(n1970), .Q(\mem2[124][17] ), .QN(n30751) );
  SDFFX1 \mem2_reg[124][16]  ( .D(n11404), .SI(\mem2[123][23] ), .SE(test_se), 
        .CLK(n1970), .Q(\mem2[124][16] ), .QN(n30752) );
  SDFFX1 \mem2_reg[123][23]  ( .D(n11403), .SI(\mem2[123][22] ), .SE(test_se), 
        .CLK(n1970), .Q(\mem2[123][23] ), .QN(n30753) );
  SDFFX1 \mem2_reg[123][22]  ( .D(n11402), .SI(\mem2[123][21] ), .SE(test_se), 
        .CLK(n1970), .Q(\mem2[123][22] ), .QN(n30754) );
  SDFFX1 \mem2_reg[123][21]  ( .D(n11401), .SI(\mem2[123][20] ), .SE(test_se), 
        .CLK(n1970), .Q(\mem2[123][21] ), .QN(n30755) );
  SDFFX1 \mem2_reg[123][20]  ( .D(n11400), .SI(\mem2[123][19] ), .SE(test_se), 
        .CLK(n1970), .Q(\mem2[123][20] ), .QN(n30756) );
  SDFFX1 \mem2_reg[123][19]  ( .D(n11399), .SI(\mem2[123][18] ), .SE(test_se), 
        .CLK(n1970), .Q(\mem2[123][19] ), .QN(n30757) );
  SDFFX1 \mem2_reg[123][18]  ( .D(n11398), .SI(\mem2[123][17] ), .SE(test_se), 
        .CLK(n1970), .Q(\mem2[123][18] ), .QN(n30758) );
  SDFFX1 \mem2_reg[123][17]  ( .D(n11397), .SI(\mem2[123][16] ), .SE(test_se), 
        .CLK(n1971), .Q(\mem2[123][17] ), .QN(n30759) );
  SDFFX1 \mem2_reg[123][16]  ( .D(n11396), .SI(\mem2[122][23] ), .SE(test_se), 
        .CLK(n1971), .Q(\mem2[123][16] ), .QN(n30760) );
  SDFFX1 \mem2_reg[122][23]  ( .D(n11395), .SI(\mem2[122][22] ), .SE(test_se), 
        .CLK(n1971), .Q(\mem2[122][23] ), .QN(n30761) );
  SDFFX1 \mem2_reg[122][22]  ( .D(n11394), .SI(\mem2[122][21] ), .SE(test_se), 
        .CLK(n1971), .Q(\mem2[122][22] ), .QN(n30762) );
  SDFFX1 \mem2_reg[122][21]  ( .D(n11393), .SI(\mem2[122][20] ), .SE(test_se), 
        .CLK(n1971), .Q(\mem2[122][21] ), .QN(n30763) );
  SDFFX1 \mem2_reg[122][20]  ( .D(n11392), .SI(\mem2[122][19] ), .SE(test_se), 
        .CLK(n1971), .Q(\mem2[122][20] ), .QN(n30764) );
  SDFFX1 \mem2_reg[122][19]  ( .D(n11391), .SI(\mem2[122][18] ), .SE(test_se), 
        .CLK(n1971), .Q(\mem2[122][19] ), .QN(n30765) );
  SDFFX1 \mem2_reg[122][18]  ( .D(n11390), .SI(\mem2[122][17] ), .SE(test_se), 
        .CLK(n1971), .Q(\mem2[122][18] ), .QN(n30766) );
  SDFFX1 \mem2_reg[122][17]  ( .D(n11389), .SI(\mem2[122][16] ), .SE(test_se), 
        .CLK(n1971), .Q(\mem2[122][17] ), .QN(n30767) );
  SDFFX1 \mem2_reg[122][16]  ( .D(n11388), .SI(\mem2[121][23] ), .SE(test_se), 
        .CLK(n1971), .Q(\mem2[122][16] ), .QN(n30768) );
  SDFFX1 \mem2_reg[121][23]  ( .D(n11387), .SI(\mem2[121][22] ), .SE(test_se), 
        .CLK(n1971), .Q(\mem2[121][23] ), .QN(n30769) );
  SDFFX1 \mem2_reg[121][22]  ( .D(n11386), .SI(\mem2[121][21] ), .SE(test_se), 
        .CLK(n1971), .Q(\mem2[121][22] ), .QN(n30770) );
  SDFFX1 \mem2_reg[121][21]  ( .D(n11385), .SI(\mem2[121][20] ), .SE(test_se), 
        .CLK(n1972), .Q(\mem2[121][21] ), .QN(n30771) );
  SDFFX1 \mem2_reg[121][20]  ( .D(n11384), .SI(\mem2[121][19] ), .SE(test_se), 
        .CLK(n1972), .Q(\mem2[121][20] ), .QN(n30772) );
  SDFFX1 \mem2_reg[121][19]  ( .D(n11383), .SI(\mem2[121][18] ), .SE(test_se), 
        .CLK(n1972), .Q(\mem2[121][19] ), .QN(n30773) );
  SDFFX1 \mem2_reg[121][18]  ( .D(n11382), .SI(\mem2[121][17] ), .SE(test_se), 
        .CLK(n1972), .Q(\mem2[121][18] ), .QN(n30774) );
  SDFFX1 \mem2_reg[121][17]  ( .D(n11381), .SI(\mem2[121][16] ), .SE(test_se), 
        .CLK(n1972), .Q(\mem2[121][17] ), .QN(n30775) );
  SDFFX1 \mem2_reg[121][16]  ( .D(n11380), .SI(\mem2[120][23] ), .SE(test_se), 
        .CLK(n1972), .Q(\mem2[121][16] ), .QN(n30776) );
  SDFFX1 \mem2_reg[120][23]  ( .D(n11379), .SI(\mem2[120][22] ), .SE(test_se), 
        .CLK(n1972), .Q(\mem2[120][23] ), .QN(n30777) );
  SDFFX1 \mem2_reg[120][22]  ( .D(n11378), .SI(\mem2[120][21] ), .SE(test_se), 
        .CLK(n1972), .Q(\mem2[120][22] ), .QN(n30778) );
  SDFFX1 \mem2_reg[120][21]  ( .D(n11377), .SI(\mem2[120][20] ), .SE(test_se), 
        .CLK(n1972), .Q(\mem2[120][21] ), .QN(n30779) );
  SDFFX1 \mem2_reg[120][20]  ( .D(n11376), .SI(\mem2[120][19] ), .SE(test_se), 
        .CLK(n1972), .Q(\mem2[120][20] ), .QN(n30780) );
  SDFFX1 \mem2_reg[120][19]  ( .D(n11375), .SI(\mem2[120][18] ), .SE(test_se), 
        .CLK(n1972), .Q(\mem2[120][19] ), .QN(n30781) );
  SDFFX1 \mem2_reg[120][18]  ( .D(n11374), .SI(\mem2[120][17] ), .SE(test_se), 
        .CLK(n1972), .Q(\mem2[120][18] ), .QN(n30782) );
  SDFFX1 \mem2_reg[120][17]  ( .D(n11373), .SI(\mem2[120][16] ), .SE(test_se), 
        .CLK(n1973), .Q(\mem2[120][17] ), .QN(n30783) );
  SDFFX1 \mem2_reg[120][16]  ( .D(n11372), .SI(\mem2[119][23] ), .SE(test_se), 
        .CLK(n1973), .Q(\mem2[120][16] ), .QN(n30784) );
  SDFFX1 \mem2_reg[119][23]  ( .D(n11371), .SI(\mem2[119][22] ), .SE(test_se), 
        .CLK(n1973), .Q(\mem2[119][23] ), .QN(n30785) );
  SDFFX1 \mem2_reg[119][22]  ( .D(n11370), .SI(\mem2[119][21] ), .SE(test_se), 
        .CLK(n1973), .Q(\mem2[119][22] ), .QN(n30786) );
  SDFFX1 \mem2_reg[119][21]  ( .D(n11369), .SI(\mem2[119][20] ), .SE(test_se), 
        .CLK(n1973), .Q(\mem2[119][21] ), .QN(n30787) );
  SDFFX1 \mem2_reg[119][20]  ( .D(n11368), .SI(\mem2[119][19] ), .SE(test_se), 
        .CLK(n1973), .Q(\mem2[119][20] ), .QN(n30788) );
  SDFFX1 \mem2_reg[119][19]  ( .D(n11367), .SI(\mem2[119][18] ), .SE(test_se), 
        .CLK(n1973), .Q(\mem2[119][19] ), .QN(n30789) );
  SDFFX1 \mem2_reg[119][18]  ( .D(n11366), .SI(\mem2[119][17] ), .SE(test_se), 
        .CLK(n1973), .Q(\mem2[119][18] ), .QN(n30790) );
  SDFFX1 \mem2_reg[119][17]  ( .D(n11365), .SI(\mem2[119][16] ), .SE(test_se), 
        .CLK(n1973), .Q(\mem2[119][17] ), .QN(n30791) );
  SDFFX1 \mem2_reg[119][16]  ( .D(n11364), .SI(\mem2[118][23] ), .SE(test_se), 
        .CLK(n1973), .Q(\mem2[119][16] ), .QN(n30792) );
  SDFFX1 \mem2_reg[118][23]  ( .D(n11363), .SI(\mem2[118][22] ), .SE(test_se), 
        .CLK(n1973), .Q(\mem2[118][23] ), .QN(n30793) );
  SDFFX1 \mem2_reg[118][22]  ( .D(n11362), .SI(\mem2[118][21] ), .SE(test_se), 
        .CLK(n1973), .Q(\mem2[118][22] ), .QN(n30794) );
  SDFFX1 \mem2_reg[118][21]  ( .D(n11361), .SI(\mem2[118][20] ), .SE(test_se), 
        .CLK(n1974), .Q(\mem2[118][21] ), .QN(n30795) );
  SDFFX1 \mem2_reg[118][20]  ( .D(n11360), .SI(\mem2[118][19] ), .SE(test_se), 
        .CLK(n1974), .Q(\mem2[118][20] ), .QN(n30796) );
  SDFFX1 \mem2_reg[118][19]  ( .D(n11359), .SI(\mem2[118][18] ), .SE(test_se), 
        .CLK(n1974), .Q(\mem2[118][19] ), .QN(n30797) );
  SDFFX1 \mem2_reg[118][18]  ( .D(n11358), .SI(\mem2[118][17] ), .SE(test_se), 
        .CLK(n1974), .Q(\mem2[118][18] ), .QN(n30798) );
  SDFFX1 \mem2_reg[118][17]  ( .D(n11357), .SI(\mem2[118][16] ), .SE(test_se), 
        .CLK(n1974), .Q(\mem2[118][17] ), .QN(n30799) );
  SDFFX1 \mem2_reg[118][16]  ( .D(n11356), .SI(\mem2[117][23] ), .SE(test_se), 
        .CLK(n1974), .Q(\mem2[118][16] ), .QN(n30800) );
  SDFFX1 \mem2_reg[117][23]  ( .D(n11355), .SI(\mem2[117][22] ), .SE(test_se), 
        .CLK(n1974), .Q(\mem2[117][23] ), .QN(n30801) );
  SDFFX1 \mem2_reg[117][22]  ( .D(n11354), .SI(\mem2[117][21] ), .SE(test_se), 
        .CLK(n1974), .Q(\mem2[117][22] ), .QN(n30802) );
  SDFFX1 \mem2_reg[117][21]  ( .D(n11353), .SI(\mem2[117][20] ), .SE(test_se), 
        .CLK(n1974), .Q(\mem2[117][21] ), .QN(n30803) );
  SDFFX1 \mem2_reg[117][20]  ( .D(n11352), .SI(\mem2[117][19] ), .SE(test_se), 
        .CLK(n1974), .Q(\mem2[117][20] ), .QN(n30804) );
  SDFFX1 \mem2_reg[117][19]  ( .D(n11351), .SI(\mem2[117][18] ), .SE(test_se), 
        .CLK(n1974), .Q(\mem2[117][19] ), .QN(n30805) );
  SDFFX1 \mem2_reg[117][18]  ( .D(n11350), .SI(\mem2[117][17] ), .SE(test_se), 
        .CLK(n1974), .Q(\mem2[117][18] ), .QN(n30806) );
  SDFFX1 \mem2_reg[117][17]  ( .D(n11349), .SI(\mem2[117][16] ), .SE(test_se), 
        .CLK(n1975), .Q(\mem2[117][17] ), .QN(n30807) );
  SDFFX1 \mem2_reg[117][16]  ( .D(n11348), .SI(\mem2[116][23] ), .SE(test_se), 
        .CLK(n1975), .Q(\mem2[117][16] ), .QN(n30808) );
  SDFFX1 \mem2_reg[116][23]  ( .D(n11347), .SI(\mem2[116][22] ), .SE(test_se), 
        .CLK(n1975), .Q(\mem2[116][23] ), .QN(n30809) );
  SDFFX1 \mem2_reg[116][22]  ( .D(n11346), .SI(\mem2[116][21] ), .SE(test_se), 
        .CLK(n1975), .Q(\mem2[116][22] ), .QN(n30810) );
  SDFFX1 \mem2_reg[116][21]  ( .D(n11345), .SI(\mem2[116][20] ), .SE(test_se), 
        .CLK(n1975), .Q(\mem2[116][21] ), .QN(n30811) );
  SDFFX1 \mem2_reg[116][20]  ( .D(n11344), .SI(\mem2[116][19] ), .SE(test_se), 
        .CLK(n1975), .Q(\mem2[116][20] ), .QN(n30812) );
  SDFFX1 \mem2_reg[116][19]  ( .D(n11343), .SI(\mem2[116][18] ), .SE(test_se), 
        .CLK(n1975), .Q(\mem2[116][19] ), .QN(n30813) );
  SDFFX1 \mem2_reg[116][18]  ( .D(n11342), .SI(\mem2[116][17] ), .SE(test_se), 
        .CLK(n1975), .Q(\mem2[116][18] ), .QN(n30814) );
  SDFFX1 \mem2_reg[116][17]  ( .D(n11341), .SI(\mem2[116][16] ), .SE(test_se), 
        .CLK(n1975), .Q(\mem2[116][17] ), .QN(n30815) );
  SDFFX1 \mem2_reg[116][16]  ( .D(n11340), .SI(\mem2[115][23] ), .SE(test_se), 
        .CLK(n1975), .Q(\mem2[116][16] ), .QN(n30816) );
  SDFFX1 \mem2_reg[115][23]  ( .D(n11339), .SI(\mem2[115][22] ), .SE(test_se), 
        .CLK(n1975), .Q(\mem2[115][23] ), .QN(n30817) );
  SDFFX1 \mem2_reg[115][22]  ( .D(n11338), .SI(\mem2[115][21] ), .SE(test_se), 
        .CLK(n1975), .Q(\mem2[115][22] ), .QN(n30818) );
  SDFFX1 \mem2_reg[115][21]  ( .D(n11337), .SI(\mem2[115][20] ), .SE(test_se), 
        .CLK(n1976), .Q(\mem2[115][21] ), .QN(n30819) );
  SDFFX1 \mem2_reg[115][20]  ( .D(n11336), .SI(\mem2[115][19] ), .SE(test_se), 
        .CLK(n1976), .Q(\mem2[115][20] ), .QN(n30820) );
  SDFFX1 \mem2_reg[115][19]  ( .D(n11335), .SI(\mem2[115][18] ), .SE(test_se), 
        .CLK(n1976), .Q(\mem2[115][19] ), .QN(n30821) );
  SDFFX1 \mem2_reg[115][18]  ( .D(n11334), .SI(\mem2[115][17] ), .SE(test_se), 
        .CLK(n1976), .Q(\mem2[115][18] ), .QN(n30822) );
  SDFFX1 \mem2_reg[115][17]  ( .D(n11333), .SI(\mem2[115][16] ), .SE(test_se), 
        .CLK(n1976), .Q(\mem2[115][17] ), .QN(n30823) );
  SDFFX1 \mem2_reg[115][16]  ( .D(n11332), .SI(\mem2[114][23] ), .SE(test_se), 
        .CLK(n1976), .Q(\mem2[115][16] ), .QN(n30824) );
  SDFFX1 \mem2_reg[114][23]  ( .D(n11331), .SI(\mem2[114][22] ), .SE(test_se), 
        .CLK(n1976), .Q(\mem2[114][23] ), .QN(n30825) );
  SDFFX1 \mem2_reg[114][22]  ( .D(n11330), .SI(\mem2[114][21] ), .SE(test_se), 
        .CLK(n1976), .Q(\mem2[114][22] ), .QN(n30826) );
  SDFFX1 \mem2_reg[114][21]  ( .D(n11329), .SI(\mem2[114][20] ), .SE(test_se), 
        .CLK(n1976), .Q(\mem2[114][21] ), .QN(n30827) );
  SDFFX1 \mem2_reg[114][20]  ( .D(n11328), .SI(\mem2[114][19] ), .SE(test_se), 
        .CLK(n1976), .Q(\mem2[114][20] ), .QN(n30828) );
  SDFFX1 \mem2_reg[114][19]  ( .D(n11327), .SI(\mem2[114][18] ), .SE(test_se), 
        .CLK(n1976), .Q(\mem2[114][19] ), .QN(n30829) );
  SDFFX1 \mem2_reg[114][18]  ( .D(n11326), .SI(\mem2[114][17] ), .SE(test_se), 
        .CLK(n1976), .Q(\mem2[114][18] ), .QN(n30830) );
  SDFFX1 \mem2_reg[114][17]  ( .D(n11325), .SI(\mem2[114][16] ), .SE(test_se), 
        .CLK(n1977), .Q(\mem2[114][17] ), .QN(n30831) );
  SDFFX1 \mem2_reg[114][16]  ( .D(n11324), .SI(\mem2[113][23] ), .SE(test_se), 
        .CLK(n1977), .Q(\mem2[114][16] ), .QN(n30832) );
  SDFFX1 \mem2_reg[113][23]  ( .D(n11323), .SI(\mem2[113][22] ), .SE(test_se), 
        .CLK(n1977), .Q(\mem2[113][23] ), .QN(n30833) );
  SDFFX1 \mem2_reg[113][22]  ( .D(n11322), .SI(\mem2[113][21] ), .SE(test_se), 
        .CLK(n1977), .Q(\mem2[113][22] ), .QN(n30834) );
  SDFFX1 \mem2_reg[113][21]  ( .D(n11321), .SI(\mem2[113][20] ), .SE(test_se), 
        .CLK(n1977), .Q(\mem2[113][21] ), .QN(n30835) );
  SDFFX1 \mem2_reg[113][20]  ( .D(n11320), .SI(\mem2[113][19] ), .SE(test_se), 
        .CLK(n1977), .Q(\mem2[113][20] ), .QN(n30836) );
  SDFFX1 \mem2_reg[113][19]  ( .D(n11319), .SI(\mem2[113][18] ), .SE(test_se), 
        .CLK(n1977), .Q(\mem2[113][19] ), .QN(n30837) );
  SDFFX1 \mem2_reg[113][18]  ( .D(n11318), .SI(\mem2[113][17] ), .SE(test_se), 
        .CLK(n1977), .Q(\mem2[113][18] ), .QN(n30838) );
  SDFFX1 \mem2_reg[113][17]  ( .D(n11317), .SI(\mem2[113][16] ), .SE(test_se), 
        .CLK(n1977), .Q(\mem2[113][17] ), .QN(n30839) );
  SDFFX1 \mem2_reg[113][16]  ( .D(n11316), .SI(\mem2[112][23] ), .SE(test_se), 
        .CLK(n1977), .Q(\mem2[113][16] ), .QN(n30840) );
  SDFFX1 \mem2_reg[112][23]  ( .D(n11315), .SI(\mem2[112][22] ), .SE(test_se), 
        .CLK(n1977), .Q(\mem2[112][23] ), .QN(n30841) );
  SDFFX1 \mem2_reg[112][22]  ( .D(n11314), .SI(\mem2[112][21] ), .SE(test_se), 
        .CLK(n1977), .Q(\mem2[112][22] ), .QN(n30842) );
  SDFFX1 \mem2_reg[112][21]  ( .D(n11313), .SI(\mem2[112][20] ), .SE(test_se), 
        .CLK(n1978), .Q(\mem2[112][21] ), .QN(n30843) );
  SDFFX1 \mem2_reg[112][20]  ( .D(n11312), .SI(\mem2[112][19] ), .SE(test_se), 
        .CLK(n1978), .Q(\mem2[112][20] ), .QN(n30844) );
  SDFFX1 \mem2_reg[112][19]  ( .D(n11311), .SI(\mem2[112][18] ), .SE(test_se), 
        .CLK(n1978), .Q(\mem2[112][19] ), .QN(n30845) );
  SDFFX1 \mem2_reg[112][18]  ( .D(n11310), .SI(\mem2[112][17] ), .SE(test_se), 
        .CLK(n1978), .Q(\mem2[112][18] ), .QN(n30846) );
  SDFFX1 \mem2_reg[112][17]  ( .D(n11309), .SI(\mem2[112][16] ), .SE(test_se), 
        .CLK(n1978), .Q(\mem2[112][17] ), .QN(n30847) );
  SDFFX1 \mem2_reg[112][16]  ( .D(n11308), .SI(\mem2[111][23] ), .SE(test_se), 
        .CLK(n1978), .Q(\mem2[112][16] ), .QN(n30848) );
  SDFFX1 \mem2_reg[111][23]  ( .D(n11307), .SI(\mem2[111][22] ), .SE(test_se), 
        .CLK(n1978), .Q(\mem2[111][23] ), .QN(n30849) );
  SDFFX1 \mem2_reg[111][22]  ( .D(n11306), .SI(\mem2[111][21] ), .SE(test_se), 
        .CLK(n1978), .Q(\mem2[111][22] ), .QN(n30850) );
  SDFFX1 \mem2_reg[111][21]  ( .D(n11305), .SI(\mem2[111][20] ), .SE(test_se), 
        .CLK(n1978), .Q(\mem2[111][21] ), .QN(n30851) );
  SDFFX1 \mem2_reg[111][20]  ( .D(n11304), .SI(\mem2[111][19] ), .SE(test_se), 
        .CLK(n1978), .Q(\mem2[111][20] ), .QN(n30852) );
  SDFFX1 \mem2_reg[111][19]  ( .D(n11303), .SI(\mem2[111][18] ), .SE(test_se), 
        .CLK(n1978), .Q(\mem2[111][19] ), .QN(n30853) );
  SDFFX1 \mem2_reg[111][18]  ( .D(n11302), .SI(\mem2[111][17] ), .SE(test_se), 
        .CLK(n1978), .Q(\mem2[111][18] ), .QN(n30854) );
  SDFFX1 \mem2_reg[111][17]  ( .D(n11301), .SI(\mem2[111][16] ), .SE(test_se), 
        .CLK(n1979), .Q(\mem2[111][17] ), .QN(n30855) );
  SDFFX1 \mem2_reg[111][16]  ( .D(n11300), .SI(\mem2[110][23] ), .SE(test_se), 
        .CLK(n1979), .Q(\mem2[111][16] ), .QN(n30856) );
  SDFFX1 \mem2_reg[110][23]  ( .D(n11299), .SI(\mem2[110][22] ), .SE(test_se), 
        .CLK(n1979), .Q(\mem2[110][23] ), .QN(n30857) );
  SDFFX1 \mem2_reg[110][22]  ( .D(n11298), .SI(\mem2[110][21] ), .SE(test_se), 
        .CLK(n1979), .Q(\mem2[110][22] ), .QN(n30858) );
  SDFFX1 \mem2_reg[110][21]  ( .D(n11297), .SI(\mem2[110][20] ), .SE(test_se), 
        .CLK(n1979), .Q(\mem2[110][21] ), .QN(n30859) );
  SDFFX1 \mem2_reg[110][20]  ( .D(n11296), .SI(\mem2[110][19] ), .SE(test_se), 
        .CLK(n1979), .Q(\mem2[110][20] ), .QN(n30860) );
  SDFFX1 \mem2_reg[110][19]  ( .D(n11295), .SI(\mem2[110][18] ), .SE(test_se), 
        .CLK(n1979), .Q(\mem2[110][19] ), .QN(n30861) );
  SDFFX1 \mem2_reg[110][18]  ( .D(n11294), .SI(\mem2[110][17] ), .SE(test_se), 
        .CLK(n1979), .Q(\mem2[110][18] ), .QN(n30862) );
  SDFFX1 \mem2_reg[110][17]  ( .D(n11293), .SI(\mem2[110][16] ), .SE(test_se), 
        .CLK(n1979), .Q(\mem2[110][17] ), .QN(n30863) );
  SDFFX1 \mem2_reg[110][16]  ( .D(n11292), .SI(\mem2[109][23] ), .SE(test_se), 
        .CLK(n1979), .Q(\mem2[110][16] ), .QN(n30864) );
  SDFFX1 \mem2_reg[109][23]  ( .D(n11291), .SI(\mem2[109][22] ), .SE(test_se), 
        .CLK(n1979), .Q(\mem2[109][23] ), .QN(n30865) );
  SDFFX1 \mem2_reg[109][22]  ( .D(n11290), .SI(\mem2[109][21] ), .SE(test_se), 
        .CLK(n1979), .Q(\mem2[109][22] ), .QN(n30866) );
  SDFFX1 \mem2_reg[109][21]  ( .D(n11289), .SI(\mem2[109][20] ), .SE(test_se), 
        .CLK(n1980), .Q(\mem2[109][21] ), .QN(n30867) );
  SDFFX1 \mem2_reg[109][20]  ( .D(n11288), .SI(\mem2[109][19] ), .SE(test_se), 
        .CLK(n1980), .Q(\mem2[109][20] ), .QN(n30868) );
  SDFFX1 \mem2_reg[109][19]  ( .D(n11287), .SI(\mem2[109][18] ), .SE(test_se), 
        .CLK(n1980), .Q(\mem2[109][19] ), .QN(n30869) );
  SDFFX1 \mem2_reg[109][18]  ( .D(n11286), .SI(\mem2[109][17] ), .SE(test_se), 
        .CLK(n1980), .Q(\mem2[109][18] ), .QN(n30870) );
  SDFFX1 \mem2_reg[109][17]  ( .D(n11285), .SI(\mem2[109][16] ), .SE(test_se), 
        .CLK(n1980), .Q(\mem2[109][17] ), .QN(n30871) );
  SDFFX1 \mem2_reg[109][16]  ( .D(n11284), .SI(\mem2[108][23] ), .SE(test_se), 
        .CLK(n1980), .Q(\mem2[109][16] ), .QN(n30872) );
  SDFFX1 \mem2_reg[108][23]  ( .D(n11283), .SI(\mem2[108][22] ), .SE(test_se), 
        .CLK(n1980), .Q(\mem2[108][23] ), .QN(n30873) );
  SDFFX1 \mem2_reg[108][22]  ( .D(n11282), .SI(\mem2[108][21] ), .SE(test_se), 
        .CLK(n1980), .Q(\mem2[108][22] ), .QN(n30874) );
  SDFFX1 \mem2_reg[108][21]  ( .D(n11281), .SI(\mem2[108][20] ), .SE(test_se), 
        .CLK(n1980), .Q(\mem2[108][21] ), .QN(n30875) );
  SDFFX1 \mem2_reg[108][20]  ( .D(n11280), .SI(\mem2[108][19] ), .SE(test_se), 
        .CLK(n1980), .Q(\mem2[108][20] ), .QN(n30876) );
  SDFFX1 \mem2_reg[108][19]  ( .D(n11279), .SI(\mem2[108][18] ), .SE(test_se), 
        .CLK(n1980), .Q(\mem2[108][19] ), .QN(n30877) );
  SDFFX1 \mem2_reg[108][18]  ( .D(n11278), .SI(\mem2[108][17] ), .SE(test_se), 
        .CLK(n1980), .Q(\mem2[108][18] ), .QN(n30878) );
  SDFFX1 \mem2_reg[108][17]  ( .D(n11277), .SI(\mem2[108][16] ), .SE(test_se), 
        .CLK(n1981), .Q(\mem2[108][17] ), .QN(n30879) );
  SDFFX1 \mem2_reg[108][16]  ( .D(n11276), .SI(\mem2[107][23] ), .SE(test_se), 
        .CLK(n1981), .Q(\mem2[108][16] ), .QN(n30880) );
  SDFFX1 \mem2_reg[107][23]  ( .D(n11275), .SI(\mem2[107][22] ), .SE(test_se), 
        .CLK(n1981), .Q(\mem2[107][23] ), .QN(n30881) );
  SDFFX1 \mem2_reg[107][22]  ( .D(n11274), .SI(\mem2[107][21] ), .SE(test_se), 
        .CLK(n1981), .Q(\mem2[107][22] ), .QN(n30882) );
  SDFFX1 \mem2_reg[107][21]  ( .D(n11273), .SI(\mem2[107][20] ), .SE(test_se), 
        .CLK(n1981), .Q(\mem2[107][21] ), .QN(n30883) );
  SDFFX1 \mem2_reg[107][20]  ( .D(n11272), .SI(\mem2[107][19] ), .SE(test_se), 
        .CLK(n1981), .Q(\mem2[107][20] ), .QN(n30884) );
  SDFFX1 \mem2_reg[107][19]  ( .D(n11271), .SI(\mem2[107][18] ), .SE(test_se), 
        .CLK(n1981), .Q(\mem2[107][19] ), .QN(n30885) );
  SDFFX1 \mem2_reg[107][18]  ( .D(n11270), .SI(\mem2[107][17] ), .SE(test_se), 
        .CLK(n1981), .Q(\mem2[107][18] ), .QN(n30886) );
  SDFFX1 \mem2_reg[107][17]  ( .D(n11269), .SI(\mem2[107][16] ), .SE(test_se), 
        .CLK(n1981), .Q(\mem2[107][17] ), .QN(n30887) );
  SDFFX1 \mem2_reg[107][16]  ( .D(n11268), .SI(\mem2[106][23] ), .SE(test_se), 
        .CLK(n1981), .Q(\mem2[107][16] ), .QN(n30888) );
  SDFFX1 \mem2_reg[106][23]  ( .D(n11267), .SI(\mem2[106][22] ), .SE(test_se), 
        .CLK(n1981), .Q(\mem2[106][23] ), .QN(n30889) );
  SDFFX1 \mem2_reg[106][22]  ( .D(n11266), .SI(\mem2[106][21] ), .SE(test_se), 
        .CLK(n1981), .Q(\mem2[106][22] ), .QN(n30890) );
  SDFFX1 \mem2_reg[106][21]  ( .D(n11265), .SI(\mem2[106][20] ), .SE(test_se), 
        .CLK(n1982), .Q(\mem2[106][21] ), .QN(n30891) );
  SDFFX1 \mem2_reg[106][20]  ( .D(n11264), .SI(\mem2[106][19] ), .SE(test_se), 
        .CLK(n1982), .Q(\mem2[106][20] ), .QN(n30892) );
  SDFFX1 \mem2_reg[106][19]  ( .D(n11263), .SI(\mem2[106][18] ), .SE(test_se), 
        .CLK(n1982), .Q(\mem2[106][19] ), .QN(n30893) );
  SDFFX1 \mem2_reg[106][18]  ( .D(n11262), .SI(\mem2[106][17] ), .SE(test_se), 
        .CLK(n1982), .Q(\mem2[106][18] ), .QN(n30894) );
  SDFFX1 \mem2_reg[106][17]  ( .D(n11261), .SI(\mem2[106][16] ), .SE(test_se), 
        .CLK(n1982), .Q(\mem2[106][17] ), .QN(n30895) );
  SDFFX1 \mem2_reg[106][16]  ( .D(n11260), .SI(\mem2[105][23] ), .SE(test_se), 
        .CLK(n1982), .Q(\mem2[106][16] ), .QN(n30896) );
  SDFFX1 \mem2_reg[105][23]  ( .D(n11259), .SI(\mem2[105][22] ), .SE(test_se), 
        .CLK(n1982), .Q(\mem2[105][23] ), .QN(n30897) );
  SDFFX1 \mem2_reg[105][22]  ( .D(n11258), .SI(\mem2[105][21] ), .SE(test_se), 
        .CLK(n1982), .Q(\mem2[105][22] ), .QN(n30898) );
  SDFFX1 \mem2_reg[105][21]  ( .D(n11257), .SI(\mem2[105][20] ), .SE(test_se), 
        .CLK(n1982), .Q(\mem2[105][21] ), .QN(n30899) );
  SDFFX1 \mem2_reg[105][20]  ( .D(n11256), .SI(\mem2[105][19] ), .SE(test_se), 
        .CLK(n1982), .Q(\mem2[105][20] ), .QN(n30900) );
  SDFFX1 \mem2_reg[105][19]  ( .D(n11255), .SI(\mem2[105][18] ), .SE(test_se), 
        .CLK(n1982), .Q(\mem2[105][19] ), .QN(n30901) );
  SDFFX1 \mem2_reg[105][18]  ( .D(n11254), .SI(\mem2[105][17] ), .SE(test_se), 
        .CLK(n1982), .Q(\mem2[105][18] ), .QN(n30902) );
  SDFFX1 \mem2_reg[105][17]  ( .D(n11253), .SI(\mem2[105][16] ), .SE(test_se), 
        .CLK(n1983), .Q(\mem2[105][17] ), .QN(n30903) );
  SDFFX1 \mem2_reg[105][16]  ( .D(n11252), .SI(\mem2[104][23] ), .SE(test_se), 
        .CLK(n1983), .Q(\mem2[105][16] ), .QN(n30904) );
  SDFFX1 \mem2_reg[104][23]  ( .D(n11251), .SI(\mem2[104][22] ), .SE(test_se), 
        .CLK(n1983), .Q(\mem2[104][23] ), .QN(n30905) );
  SDFFX1 \mem2_reg[104][22]  ( .D(n11250), .SI(\mem2[104][21] ), .SE(test_se), 
        .CLK(n1983), .Q(\mem2[104][22] ), .QN(n30906) );
  SDFFX1 \mem2_reg[104][21]  ( .D(n11249), .SI(\mem2[104][20] ), .SE(test_se), 
        .CLK(n1983), .Q(\mem2[104][21] ), .QN(n30907) );
  SDFFX1 \mem2_reg[104][20]  ( .D(n11248), .SI(\mem2[104][19] ), .SE(test_se), 
        .CLK(n1983), .Q(\mem2[104][20] ), .QN(n30908) );
  SDFFX1 \mem2_reg[104][19]  ( .D(n11247), .SI(\mem2[104][18] ), .SE(test_se), 
        .CLK(n1983), .Q(\mem2[104][19] ), .QN(n30909) );
  SDFFX1 \mem2_reg[104][18]  ( .D(n11246), .SI(\mem2[104][17] ), .SE(test_se), 
        .CLK(n1983), .Q(\mem2[104][18] ), .QN(n30910) );
  SDFFX1 \mem2_reg[104][17]  ( .D(n11245), .SI(\mem2[104][16] ), .SE(test_se), 
        .CLK(n1983), .Q(\mem2[104][17] ), .QN(n30911) );
  SDFFX1 \mem2_reg[104][16]  ( .D(n11244), .SI(\mem2[103][23] ), .SE(test_se), 
        .CLK(n1983), .Q(\mem2[104][16] ), .QN(n30912) );
  SDFFX1 \mem2_reg[103][23]  ( .D(n11243), .SI(\mem2[103][22] ), .SE(test_se), 
        .CLK(n1983), .Q(\mem2[103][23] ), .QN(n30913) );
  SDFFX1 \mem2_reg[103][22]  ( .D(n11242), .SI(\mem2[103][21] ), .SE(test_se), 
        .CLK(n1983), .Q(\mem2[103][22] ), .QN(n30914) );
  SDFFX1 \mem2_reg[103][21]  ( .D(n11241), .SI(\mem2[103][20] ), .SE(test_se), 
        .CLK(n1984), .Q(\mem2[103][21] ), .QN(n30915) );
  SDFFX1 \mem2_reg[103][20]  ( .D(n11240), .SI(\mem2[103][19] ), .SE(test_se), 
        .CLK(n1984), .Q(\mem2[103][20] ), .QN(n30916) );
  SDFFX1 \mem2_reg[103][19]  ( .D(n11239), .SI(\mem2[103][18] ), .SE(test_se), 
        .CLK(n1984), .Q(\mem2[103][19] ), .QN(n30917) );
  SDFFX1 \mem2_reg[103][18]  ( .D(n11238), .SI(\mem2[103][17] ), .SE(test_se), 
        .CLK(n1984), .Q(\mem2[103][18] ), .QN(n30918) );
  SDFFX1 \mem2_reg[103][17]  ( .D(n11237), .SI(\mem2[103][16] ), .SE(test_se), 
        .CLK(n1984), .Q(\mem2[103][17] ), .QN(n30919) );
  SDFFX1 \mem2_reg[103][16]  ( .D(n11236), .SI(\mem2[102][23] ), .SE(test_se), 
        .CLK(n1984), .Q(\mem2[103][16] ), .QN(n30920) );
  SDFFX1 \mem2_reg[102][23]  ( .D(n11235), .SI(\mem2[102][22] ), .SE(test_se), 
        .CLK(n1984), .Q(\mem2[102][23] ), .QN(n30921) );
  SDFFX1 \mem2_reg[102][22]  ( .D(n11234), .SI(\mem2[102][21] ), .SE(test_se), 
        .CLK(n1984), .Q(\mem2[102][22] ), .QN(n30922) );
  SDFFX1 \mem2_reg[102][21]  ( .D(n11233), .SI(\mem2[102][20] ), .SE(test_se), 
        .CLK(n1984), .Q(\mem2[102][21] ), .QN(n30923) );
  SDFFX1 \mem2_reg[102][20]  ( .D(n11232), .SI(\mem2[102][19] ), .SE(test_se), 
        .CLK(n1984), .Q(\mem2[102][20] ), .QN(n30924) );
  SDFFX1 \mem2_reg[102][19]  ( .D(n11231), .SI(\mem2[102][18] ), .SE(test_se), 
        .CLK(n1984), .Q(\mem2[102][19] ), .QN(n30925) );
  SDFFX1 \mem2_reg[102][18]  ( .D(n11230), .SI(\mem2[102][17] ), .SE(test_se), 
        .CLK(n1984), .Q(\mem2[102][18] ), .QN(n30926) );
  SDFFX1 \mem2_reg[102][17]  ( .D(n11229), .SI(\mem2[102][16] ), .SE(test_se), 
        .CLK(n1985), .Q(\mem2[102][17] ), .QN(n30927) );
  SDFFX1 \mem2_reg[102][16]  ( .D(n11228), .SI(\mem2[101][23] ), .SE(test_se), 
        .CLK(n1985), .Q(\mem2[102][16] ), .QN(n30928) );
  SDFFX1 \mem2_reg[101][23]  ( .D(n11227), .SI(\mem2[101][22] ), .SE(test_se), 
        .CLK(n1985), .Q(\mem2[101][23] ), .QN(n30929) );
  SDFFX1 \mem2_reg[101][22]  ( .D(n11226), .SI(\mem2[101][21] ), .SE(test_se), 
        .CLK(n1985), .Q(\mem2[101][22] ), .QN(n30930) );
  SDFFX1 \mem2_reg[101][21]  ( .D(n11225), .SI(\mem2[101][20] ), .SE(test_se), 
        .CLK(n1985), .Q(\mem2[101][21] ), .QN(n30931) );
  SDFFX1 \mem2_reg[101][20]  ( .D(n11224), .SI(\mem2[101][19] ), .SE(test_se), 
        .CLK(n1985), .Q(\mem2[101][20] ), .QN(n30932) );
  SDFFX1 \mem2_reg[101][19]  ( .D(n11223), .SI(\mem2[101][18] ), .SE(test_se), 
        .CLK(n1985), .Q(\mem2[101][19] ), .QN(n30933) );
  SDFFX1 \mem2_reg[101][18]  ( .D(n11222), .SI(\mem2[101][17] ), .SE(test_se), 
        .CLK(n1985), .Q(\mem2[101][18] ), .QN(n30934) );
  SDFFX1 \mem2_reg[101][17]  ( .D(n11221), .SI(\mem2[101][16] ), .SE(test_se), 
        .CLK(n1985), .Q(\mem2[101][17] ), .QN(n30935) );
  SDFFX1 \mem2_reg[101][16]  ( .D(n11220), .SI(\mem2[100][23] ), .SE(test_se), 
        .CLK(n1985), .Q(\mem2[101][16] ), .QN(n30936) );
  SDFFX1 \mem2_reg[100][23]  ( .D(n11219), .SI(\mem2[100][22] ), .SE(test_se), 
        .CLK(n1985), .Q(\mem2[100][23] ), .QN(n30937) );
  SDFFX1 \mem2_reg[100][22]  ( .D(n11218), .SI(\mem2[100][21] ), .SE(test_se), 
        .CLK(n1985), .Q(\mem2[100][22] ), .QN(n30938) );
  SDFFX1 \mem2_reg[100][21]  ( .D(n11217), .SI(\mem2[100][20] ), .SE(test_se), 
        .CLK(n1986), .Q(\mem2[100][21] ), .QN(n30939) );
  SDFFX1 \mem2_reg[100][20]  ( .D(n11216), .SI(\mem2[100][19] ), .SE(test_se), 
        .CLK(n1986), .Q(\mem2[100][20] ), .QN(n30940) );
  SDFFX1 \mem2_reg[100][19]  ( .D(n11215), .SI(\mem2[100][18] ), .SE(test_se), 
        .CLK(n1986), .Q(\mem2[100][19] ), .QN(n30941) );
  SDFFX1 \mem2_reg[100][18]  ( .D(n11214), .SI(\mem2[100][17] ), .SE(test_se), 
        .CLK(n1986), .Q(\mem2[100][18] ), .QN(n30942) );
  SDFFX1 \mem2_reg[100][17]  ( .D(n11213), .SI(\mem2[100][16] ), .SE(test_se), 
        .CLK(n1986), .Q(\mem2[100][17] ), .QN(n30943) );
  SDFFX1 \mem2_reg[100][16]  ( .D(n11212), .SI(\mem2[99][23] ), .SE(test_se), 
        .CLK(n1986), .Q(\mem2[100][16] ), .QN(n30944) );
  SDFFX1 \mem2_reg[99][23]  ( .D(n11211), .SI(\mem2[99][22] ), .SE(test_se), 
        .CLK(n1986), .Q(\mem2[99][23] ), .QN(n30945) );
  SDFFX1 \mem2_reg[99][22]  ( .D(n11210), .SI(\mem2[99][21] ), .SE(test_se), 
        .CLK(n1986), .Q(\mem2[99][22] ), .QN(n30946) );
  SDFFX1 \mem2_reg[99][21]  ( .D(n11209), .SI(\mem2[99][20] ), .SE(test_se), 
        .CLK(n1986), .Q(\mem2[99][21] ), .QN(n30947) );
  SDFFX1 \mem2_reg[99][20]  ( .D(n11208), .SI(\mem2[99][19] ), .SE(test_se), 
        .CLK(n1986), .Q(\mem2[99][20] ), .QN(n30948) );
  SDFFX1 \mem2_reg[99][19]  ( .D(n11207), .SI(\mem2[99][18] ), .SE(test_se), 
        .CLK(n1986), .Q(\mem2[99][19] ), .QN(n30949) );
  SDFFX1 \mem2_reg[99][18]  ( .D(n11206), .SI(\mem2[99][17] ), .SE(test_se), 
        .CLK(n1986), .Q(\mem2[99][18] ), .QN(n30950) );
  SDFFX1 \mem2_reg[99][17]  ( .D(n11205), .SI(\mem2[99][16] ), .SE(test_se), 
        .CLK(n1987), .Q(\mem2[99][17] ), .QN(n30951) );
  SDFFX1 \mem2_reg[99][16]  ( .D(n11204), .SI(\mem2[98][23] ), .SE(test_se), 
        .CLK(n1987), .Q(\mem2[99][16] ), .QN(n30952) );
  SDFFX1 \mem2_reg[98][23]  ( .D(n11203), .SI(\mem2[98][22] ), .SE(test_se), 
        .CLK(n1987), .Q(\mem2[98][23] ), .QN(n30953) );
  SDFFX1 \mem2_reg[98][22]  ( .D(n11202), .SI(\mem2[98][21] ), .SE(test_se), 
        .CLK(n1987), .Q(\mem2[98][22] ), .QN(n30954) );
  SDFFX1 \mem2_reg[98][21]  ( .D(n11201), .SI(\mem2[98][20] ), .SE(test_se), 
        .CLK(n1987), .Q(\mem2[98][21] ), .QN(n30955) );
  SDFFX1 \mem2_reg[98][20]  ( .D(n11200), .SI(\mem2[98][19] ), .SE(test_se), 
        .CLK(n1987), .Q(\mem2[98][20] ), .QN(n30956) );
  SDFFX1 \mem2_reg[98][19]  ( .D(n11199), .SI(\mem2[98][18] ), .SE(test_se), 
        .CLK(n1987), .Q(\mem2[98][19] ), .QN(n30957) );
  SDFFX1 \mem2_reg[98][18]  ( .D(n11198), .SI(\mem2[98][17] ), .SE(test_se), 
        .CLK(n1987), .Q(\mem2[98][18] ), .QN(n30958) );
  SDFFX1 \mem2_reg[98][17]  ( .D(n11197), .SI(\mem2[98][16] ), .SE(test_se), 
        .CLK(n1987), .Q(\mem2[98][17] ), .QN(n30959) );
  SDFFX1 \mem2_reg[98][16]  ( .D(n11196), .SI(\mem2[97][23] ), .SE(test_se), 
        .CLK(n1987), .Q(\mem2[98][16] ), .QN(n30960) );
  SDFFX1 \mem2_reg[97][23]  ( .D(n11195), .SI(\mem2[97][22] ), .SE(test_se), 
        .CLK(n1987), .Q(\mem2[97][23] ), .QN(n30961) );
  SDFFX1 \mem2_reg[97][22]  ( .D(n11194), .SI(\mem2[97][21] ), .SE(test_se), 
        .CLK(n1987), .Q(\mem2[97][22] ), .QN(n30962) );
  SDFFX1 \mem2_reg[97][21]  ( .D(n11193), .SI(\mem2[97][20] ), .SE(test_se), 
        .CLK(n1988), .Q(\mem2[97][21] ), .QN(n30963) );
  SDFFX1 \mem2_reg[97][20]  ( .D(n11192), .SI(\mem2[97][19] ), .SE(test_se), 
        .CLK(n1988), .Q(\mem2[97][20] ), .QN(n30964) );
  SDFFX1 \mem2_reg[97][19]  ( .D(n11191), .SI(\mem2[97][18] ), .SE(test_se), 
        .CLK(n1988), .Q(\mem2[97][19] ), .QN(n30965) );
  SDFFX1 \mem2_reg[97][18]  ( .D(n11190), .SI(\mem2[97][17] ), .SE(test_se), 
        .CLK(n1988), .Q(\mem2[97][18] ), .QN(n30966) );
  SDFFX1 \mem2_reg[97][17]  ( .D(n11189), .SI(\mem2[97][16] ), .SE(test_se), 
        .CLK(n1988), .Q(\mem2[97][17] ), .QN(n30967) );
  SDFFX1 \mem2_reg[97][16]  ( .D(n11188), .SI(\mem2[96][23] ), .SE(test_se), 
        .CLK(n1988), .Q(\mem2[97][16] ), .QN(n30968) );
  SDFFX1 \mem2_reg[96][23]  ( .D(n11187), .SI(\mem2[96][22] ), .SE(test_se), 
        .CLK(n1988), .Q(\mem2[96][23] ), .QN(n30969) );
  SDFFX1 \mem2_reg[96][22]  ( .D(n11186), .SI(\mem2[96][21] ), .SE(test_se), 
        .CLK(n1988), .Q(\mem2[96][22] ), .QN(n30970) );
  SDFFX1 \mem2_reg[96][21]  ( .D(n11185), .SI(\mem2[96][20] ), .SE(test_se), 
        .CLK(n1988), .Q(\mem2[96][21] ), .QN(n30971) );
  SDFFX1 \mem2_reg[96][20]  ( .D(n11184), .SI(\mem2[96][19] ), .SE(test_se), 
        .CLK(n1988), .Q(\mem2[96][20] ), .QN(n30972) );
  SDFFX1 \mem2_reg[96][19]  ( .D(n11183), .SI(\mem2[96][18] ), .SE(test_se), 
        .CLK(n1988), .Q(\mem2[96][19] ), .QN(n30973) );
  SDFFX1 \mem2_reg[96][18]  ( .D(n11182), .SI(\mem2[96][17] ), .SE(test_se), 
        .CLK(n1988), .Q(\mem2[96][18] ), .QN(n30974) );
  SDFFX1 \mem2_reg[96][17]  ( .D(n11181), .SI(\mem2[96][16] ), .SE(test_se), 
        .CLK(n1989), .Q(\mem2[96][17] ), .QN(n30975) );
  SDFFX1 \mem2_reg[96][16]  ( .D(n11180), .SI(\mem2[95][23] ), .SE(test_se), 
        .CLK(n1989), .Q(\mem2[96][16] ), .QN(n30976) );
  SDFFX1 \mem2_reg[95][23]  ( .D(n11179), .SI(\mem2[95][22] ), .SE(test_se), 
        .CLK(n1989), .Q(\mem2[95][23] ), .QN(n30977) );
  SDFFX1 \mem2_reg[95][22]  ( .D(n11178), .SI(\mem2[95][21] ), .SE(test_se), 
        .CLK(n1989), .Q(\mem2[95][22] ), .QN(n30978) );
  SDFFX1 \mem2_reg[95][21]  ( .D(n11177), .SI(\mem2[95][20] ), .SE(test_se), 
        .CLK(n1989), .Q(\mem2[95][21] ), .QN(n30979) );
  SDFFX1 \mem2_reg[95][20]  ( .D(n11176), .SI(\mem2[95][19] ), .SE(test_se), 
        .CLK(n1989), .Q(\mem2[95][20] ), .QN(n30980) );
  SDFFX1 \mem2_reg[95][19]  ( .D(n11175), .SI(\mem2[95][18] ), .SE(test_se), 
        .CLK(n1989), .Q(\mem2[95][19] ), .QN(n30981) );
  SDFFX1 \mem2_reg[95][18]  ( .D(n11174), .SI(\mem2[95][17] ), .SE(test_se), 
        .CLK(n1989), .Q(\mem2[95][18] ), .QN(n30982) );
  SDFFX1 \mem2_reg[95][17]  ( .D(n11173), .SI(\mem2[95][16] ), .SE(test_se), 
        .CLK(n1989), .Q(\mem2[95][17] ), .QN(n30983) );
  SDFFX1 \mem2_reg[95][16]  ( .D(n11172), .SI(\mem2[94][23] ), .SE(test_se), 
        .CLK(n1989), .Q(\mem2[95][16] ), .QN(n30984) );
  SDFFX1 \mem2_reg[94][23]  ( .D(n11171), .SI(\mem2[94][22] ), .SE(test_se), 
        .CLK(n1989), .Q(\mem2[94][23] ), .QN(n30985) );
  SDFFX1 \mem2_reg[94][22]  ( .D(n11170), .SI(\mem2[94][21] ), .SE(test_se), 
        .CLK(n1989), .Q(\mem2[94][22] ), .QN(n30986) );
  SDFFX1 \mem2_reg[94][21]  ( .D(n11169), .SI(\mem2[94][20] ), .SE(test_se), 
        .CLK(n1990), .Q(\mem2[94][21] ), .QN(n30987) );
  SDFFX1 \mem2_reg[94][20]  ( .D(n11168), .SI(\mem2[94][19] ), .SE(test_se), 
        .CLK(n1990), .Q(\mem2[94][20] ), .QN(n30988) );
  SDFFX1 \mem2_reg[94][19]  ( .D(n11167), .SI(\mem2[94][18] ), .SE(test_se), 
        .CLK(n1990), .Q(\mem2[94][19] ), .QN(n30989) );
  SDFFX1 \mem2_reg[94][18]  ( .D(n11166), .SI(\mem2[94][17] ), .SE(test_se), 
        .CLK(n1990), .Q(\mem2[94][18] ), .QN(n30990) );
  SDFFX1 \mem2_reg[94][17]  ( .D(n11165), .SI(\mem2[94][16] ), .SE(test_se), 
        .CLK(n1990), .Q(\mem2[94][17] ), .QN(n30991) );
  SDFFX1 \mem2_reg[94][16]  ( .D(n11164), .SI(\mem2[93][23] ), .SE(test_se), 
        .CLK(n1990), .Q(\mem2[94][16] ), .QN(n30992) );
  SDFFX1 \mem2_reg[93][23]  ( .D(n11163), .SI(\mem2[93][22] ), .SE(test_se), 
        .CLK(n1990), .Q(\mem2[93][23] ), .QN(n30993) );
  SDFFX1 \mem2_reg[93][22]  ( .D(n11162), .SI(\mem2[93][21] ), .SE(test_se), 
        .CLK(n1990), .Q(\mem2[93][22] ), .QN(n30994) );
  SDFFX1 \mem2_reg[93][21]  ( .D(n11161), .SI(\mem2[93][20] ), .SE(test_se), 
        .CLK(n1990), .Q(\mem2[93][21] ), .QN(n30995) );
  SDFFX1 \mem2_reg[93][20]  ( .D(n11160), .SI(\mem2[93][19] ), .SE(test_se), 
        .CLK(n1990), .Q(\mem2[93][20] ), .QN(n30996) );
  SDFFX1 \mem2_reg[93][19]  ( .D(n11159), .SI(\mem2[93][18] ), .SE(test_se), 
        .CLK(n1990), .Q(\mem2[93][19] ), .QN(n30997) );
  SDFFX1 \mem2_reg[93][18]  ( .D(n11158), .SI(\mem2[93][17] ), .SE(test_se), 
        .CLK(n1990), .Q(\mem2[93][18] ), .QN(n30998) );
  SDFFX1 \mem2_reg[93][17]  ( .D(n11157), .SI(\mem2[93][16] ), .SE(test_se), 
        .CLK(n1991), .Q(\mem2[93][17] ), .QN(n30999) );
  SDFFX1 \mem2_reg[93][16]  ( .D(n11156), .SI(\mem2[92][23] ), .SE(test_se), 
        .CLK(n1991), .Q(\mem2[93][16] ), .QN(n31000) );
  SDFFX1 \mem2_reg[92][23]  ( .D(n11155), .SI(\mem2[92][22] ), .SE(test_se), 
        .CLK(n1991), .Q(\mem2[92][23] ), .QN(n31001) );
  SDFFX1 \mem2_reg[92][22]  ( .D(n11154), .SI(\mem2[92][21] ), .SE(test_se), 
        .CLK(n1991), .Q(\mem2[92][22] ), .QN(n31002) );
  SDFFX1 \mem2_reg[92][21]  ( .D(n11153), .SI(\mem2[92][20] ), .SE(test_se), 
        .CLK(n1991), .Q(\mem2[92][21] ), .QN(n31003) );
  SDFFX1 \mem2_reg[92][20]  ( .D(n11152), .SI(\mem2[92][19] ), .SE(test_se), 
        .CLK(n1991), .Q(\mem2[92][20] ), .QN(n31004) );
  SDFFX1 \mem2_reg[92][19]  ( .D(n11151), .SI(\mem2[92][18] ), .SE(test_se), 
        .CLK(n1991), .Q(\mem2[92][19] ), .QN(n31005) );
  SDFFX1 \mem2_reg[92][18]  ( .D(n11150), .SI(\mem2[92][17] ), .SE(test_se), 
        .CLK(n1991), .Q(\mem2[92][18] ), .QN(n31006) );
  SDFFX1 \mem2_reg[92][17]  ( .D(n11149), .SI(\mem2[92][16] ), .SE(test_se), 
        .CLK(n1991), .Q(\mem2[92][17] ), .QN(n31007) );
  SDFFX1 \mem2_reg[92][16]  ( .D(n11148), .SI(\mem2[91][23] ), .SE(test_se), 
        .CLK(n1991), .Q(\mem2[92][16] ), .QN(n31008) );
  SDFFX1 \mem2_reg[91][23]  ( .D(n11147), .SI(\mem2[91][22] ), .SE(test_se), 
        .CLK(n1991), .Q(\mem2[91][23] ), .QN(n31009) );
  SDFFX1 \mem2_reg[91][22]  ( .D(n11146), .SI(\mem2[91][21] ), .SE(test_se), 
        .CLK(n1991), .Q(\mem2[91][22] ), .QN(n31010) );
  SDFFX1 \mem2_reg[91][21]  ( .D(n11145), .SI(\mem2[91][20] ), .SE(test_se), 
        .CLK(n1992), .Q(\mem2[91][21] ), .QN(n31011) );
  SDFFX1 \mem2_reg[91][20]  ( .D(n11144), .SI(\mem2[91][19] ), .SE(test_se), 
        .CLK(n1992), .Q(\mem2[91][20] ), .QN(n31012) );
  SDFFX1 \mem2_reg[91][19]  ( .D(n11143), .SI(\mem2[91][18] ), .SE(test_se), 
        .CLK(n1992), .Q(\mem2[91][19] ), .QN(n31013) );
  SDFFX1 \mem2_reg[91][18]  ( .D(n11142), .SI(\mem2[91][17] ), .SE(test_se), 
        .CLK(n1992), .Q(\mem2[91][18] ), .QN(n31014) );
  SDFFX1 \mem2_reg[91][17]  ( .D(n11141), .SI(\mem2[91][16] ), .SE(test_se), 
        .CLK(n1992), .Q(\mem2[91][17] ), .QN(n31015) );
  SDFFX1 \mem2_reg[91][16]  ( .D(n11140), .SI(\mem2[90][23] ), .SE(test_se), 
        .CLK(n1992), .Q(\mem2[91][16] ), .QN(n31016) );
  SDFFX1 \mem2_reg[90][23]  ( .D(n11139), .SI(\mem2[90][22] ), .SE(test_se), 
        .CLK(n1992), .Q(\mem2[90][23] ), .QN(n31017) );
  SDFFX1 \mem2_reg[90][22]  ( .D(n11138), .SI(\mem2[90][21] ), .SE(test_se), 
        .CLK(n1992), .Q(\mem2[90][22] ), .QN(n31018) );
  SDFFX1 \mem2_reg[90][21]  ( .D(n11137), .SI(\mem2[90][20] ), .SE(test_se), 
        .CLK(n1992), .Q(\mem2[90][21] ), .QN(n31019) );
  SDFFX1 \mem2_reg[90][20]  ( .D(n11136), .SI(\mem2[90][19] ), .SE(test_se), 
        .CLK(n1992), .Q(\mem2[90][20] ), .QN(n31020) );
  SDFFX1 \mem2_reg[90][19]  ( .D(n11135), .SI(\mem2[90][18] ), .SE(test_se), 
        .CLK(n1992), .Q(\mem2[90][19] ), .QN(n31021) );
  SDFFX1 \mem2_reg[90][18]  ( .D(n11134), .SI(\mem2[90][17] ), .SE(test_se), 
        .CLK(n1992), .Q(\mem2[90][18] ), .QN(n31022) );
  SDFFX1 \mem2_reg[90][17]  ( .D(n11133), .SI(\mem2[90][16] ), .SE(test_se), 
        .CLK(n1993), .Q(\mem2[90][17] ), .QN(n31023) );
  SDFFX1 \mem2_reg[90][16]  ( .D(n11132), .SI(\mem2[89][23] ), .SE(test_se), 
        .CLK(n1993), .Q(\mem2[90][16] ), .QN(n31024) );
  SDFFX1 \mem2_reg[89][23]  ( .D(n11131), .SI(\mem2[89][22] ), .SE(test_se), 
        .CLK(n1993), .Q(\mem2[89][23] ), .QN(n31025) );
  SDFFX1 \mem2_reg[89][22]  ( .D(n11130), .SI(\mem2[89][21] ), .SE(test_se), 
        .CLK(n1993), .Q(\mem2[89][22] ), .QN(n31026) );
  SDFFX1 \mem2_reg[89][21]  ( .D(n11129), .SI(\mem2[89][20] ), .SE(test_se), 
        .CLK(n1993), .Q(\mem2[89][21] ), .QN(n31027) );
  SDFFX1 \mem2_reg[89][20]  ( .D(n11128), .SI(\mem2[89][19] ), .SE(test_se), 
        .CLK(n1993), .Q(\mem2[89][20] ), .QN(n31028) );
  SDFFX1 \mem2_reg[89][19]  ( .D(n11127), .SI(\mem2[89][18] ), .SE(test_se), 
        .CLK(n1993), .Q(\mem2[89][19] ), .QN(n31029) );
  SDFFX1 \mem2_reg[89][18]  ( .D(n11126), .SI(\mem2[89][17] ), .SE(test_se), 
        .CLK(n1993), .Q(\mem2[89][18] ), .QN(n31030) );
  SDFFX1 \mem2_reg[89][17]  ( .D(n11125), .SI(\mem2[89][16] ), .SE(test_se), 
        .CLK(n1993), .Q(\mem2[89][17] ), .QN(n31031) );
  SDFFX1 \mem2_reg[89][16]  ( .D(n11124), .SI(\mem2[88][23] ), .SE(test_se), 
        .CLK(n1993), .Q(\mem2[89][16] ), .QN(n31032) );
  SDFFX1 \mem2_reg[88][23]  ( .D(n11123), .SI(\mem2[88][22] ), .SE(test_se), 
        .CLK(n1993), .Q(\mem2[88][23] ), .QN(n31033) );
  SDFFX1 \mem2_reg[88][22]  ( .D(n11122), .SI(\mem2[88][21] ), .SE(test_se), 
        .CLK(n1993), .Q(\mem2[88][22] ), .QN(n31034) );
  SDFFX1 \mem2_reg[88][21]  ( .D(n11121), .SI(\mem2[88][20] ), .SE(test_se), 
        .CLK(n1994), .Q(\mem2[88][21] ), .QN(n31035) );
  SDFFX1 \mem2_reg[88][20]  ( .D(n11120), .SI(\mem2[88][19] ), .SE(test_se), 
        .CLK(n1994), .Q(\mem2[88][20] ), .QN(n31036) );
  SDFFX1 \mem2_reg[88][19]  ( .D(n11119), .SI(\mem2[88][18] ), .SE(test_se), 
        .CLK(n1994), .Q(\mem2[88][19] ), .QN(n31037) );
  SDFFX1 \mem2_reg[88][18]  ( .D(n11118), .SI(\mem2[88][17] ), .SE(test_se), 
        .CLK(n1994), .Q(\mem2[88][18] ), .QN(n31038) );
  SDFFX1 \mem2_reg[88][17]  ( .D(n11117), .SI(\mem2[88][16] ), .SE(test_se), 
        .CLK(n1994), .Q(\mem2[88][17] ), .QN(n31039) );
  SDFFX1 \mem2_reg[88][16]  ( .D(n11116), .SI(\mem2[87][23] ), .SE(test_se), 
        .CLK(n1994), .Q(\mem2[88][16] ), .QN(n31040) );
  SDFFX1 \mem2_reg[87][23]  ( .D(n11115), .SI(\mem2[87][22] ), .SE(test_se), 
        .CLK(n1994), .Q(\mem2[87][23] ), .QN(n31041) );
  SDFFX1 \mem2_reg[87][22]  ( .D(n11114), .SI(\mem2[87][21] ), .SE(test_se), 
        .CLK(n1994), .Q(\mem2[87][22] ), .QN(n31042) );
  SDFFX1 \mem2_reg[87][21]  ( .D(n11113), .SI(\mem2[87][20] ), .SE(test_se), 
        .CLK(n1994), .Q(\mem2[87][21] ), .QN(n31043) );
  SDFFX1 \mem2_reg[87][20]  ( .D(n11112), .SI(\mem2[87][19] ), .SE(test_se), 
        .CLK(n1994), .Q(\mem2[87][20] ), .QN(n31044) );
  SDFFX1 \mem2_reg[87][19]  ( .D(n11111), .SI(\mem2[87][18] ), .SE(test_se), 
        .CLK(n1994), .Q(\mem2[87][19] ), .QN(n31045) );
  SDFFX1 \mem2_reg[87][18]  ( .D(n11110), .SI(\mem2[87][17] ), .SE(test_se), 
        .CLK(n1994), .Q(\mem2[87][18] ), .QN(n31046) );
  SDFFX1 \mem2_reg[87][17]  ( .D(n11109), .SI(\mem2[87][16] ), .SE(test_se), 
        .CLK(n1995), .Q(\mem2[87][17] ), .QN(n31047) );
  SDFFX1 \mem2_reg[87][16]  ( .D(n11108), .SI(\mem2[86][23] ), .SE(test_se), 
        .CLK(n1995), .Q(\mem2[87][16] ), .QN(n31048) );
  SDFFX1 \mem2_reg[86][23]  ( .D(n11107), .SI(\mem2[86][22] ), .SE(test_se), 
        .CLK(n1995), .Q(\mem2[86][23] ), .QN(n31049) );
  SDFFX1 \mem2_reg[86][22]  ( .D(n11106), .SI(\mem2[86][21] ), .SE(test_se), 
        .CLK(n1995), .Q(\mem2[86][22] ), .QN(n31050) );
  SDFFX1 \mem2_reg[86][21]  ( .D(n11105), .SI(\mem2[86][20] ), .SE(test_se), 
        .CLK(n1995), .Q(\mem2[86][21] ), .QN(n31051) );
  SDFFX1 \mem2_reg[86][20]  ( .D(n11104), .SI(\mem2[86][19] ), .SE(test_se), 
        .CLK(n1995), .Q(\mem2[86][20] ), .QN(n31052) );
  SDFFX1 \mem2_reg[86][19]  ( .D(n11103), .SI(\mem2[86][18] ), .SE(test_se), 
        .CLK(n1995), .Q(\mem2[86][19] ), .QN(n31053) );
  SDFFX1 \mem2_reg[86][18]  ( .D(n11102), .SI(\mem2[86][17] ), .SE(test_se), 
        .CLK(n1995), .Q(\mem2[86][18] ), .QN(n31054) );
  SDFFX1 \mem2_reg[86][17]  ( .D(n11101), .SI(\mem2[86][16] ), .SE(test_se), 
        .CLK(n1995), .Q(\mem2[86][17] ), .QN(n31055) );
  SDFFX1 \mem2_reg[86][16]  ( .D(n11100), .SI(\mem2[85][23] ), .SE(test_se), 
        .CLK(n1995), .Q(\mem2[86][16] ), .QN(n31056) );
  SDFFX1 \mem2_reg[85][23]  ( .D(n11099), .SI(\mem2[85][22] ), .SE(test_se), 
        .CLK(n1995), .Q(\mem2[85][23] ), .QN(n31057) );
  SDFFX1 \mem2_reg[85][22]  ( .D(n11098), .SI(\mem2[85][21] ), .SE(test_se), 
        .CLK(n1995), .Q(\mem2[85][22] ), .QN(n31058) );
  SDFFX1 \mem2_reg[85][21]  ( .D(n11097), .SI(\mem2[85][20] ), .SE(test_se), 
        .CLK(n1996), .Q(\mem2[85][21] ), .QN(n31059) );
  SDFFX1 \mem2_reg[85][20]  ( .D(n11096), .SI(\mem2[85][19] ), .SE(test_se), 
        .CLK(n1996), .Q(\mem2[85][20] ), .QN(n31060) );
  SDFFX1 \mem2_reg[85][19]  ( .D(n11095), .SI(\mem2[85][18] ), .SE(test_se), 
        .CLK(n1996), .Q(\mem2[85][19] ), .QN(n31061) );
  SDFFX1 \mem2_reg[85][18]  ( .D(n11094), .SI(\mem2[85][17] ), .SE(test_se), 
        .CLK(n1996), .Q(\mem2[85][18] ), .QN(n31062) );
  SDFFX1 \mem2_reg[85][17]  ( .D(n11093), .SI(\mem2[85][16] ), .SE(test_se), 
        .CLK(n1996), .Q(\mem2[85][17] ), .QN(n31063) );
  SDFFX1 \mem2_reg[85][16]  ( .D(n11092), .SI(\mem2[84][23] ), .SE(test_se), 
        .CLK(n1996), .Q(\mem2[85][16] ), .QN(n31064) );
  SDFFX1 \mem2_reg[84][23]  ( .D(n11091), .SI(\mem2[84][22] ), .SE(test_se), 
        .CLK(n1996), .Q(\mem2[84][23] ), .QN(n31065) );
  SDFFX1 \mem2_reg[84][22]  ( .D(n11090), .SI(\mem2[84][21] ), .SE(test_se), 
        .CLK(n1996), .Q(\mem2[84][22] ), .QN(n31066) );
  SDFFX1 \mem2_reg[84][21]  ( .D(n11089), .SI(\mem2[84][20] ), .SE(test_se), 
        .CLK(n1996), .Q(\mem2[84][21] ), .QN(n31067) );
  SDFFX1 \mem2_reg[84][20]  ( .D(n11088), .SI(\mem2[84][19] ), .SE(test_se), 
        .CLK(n1996), .Q(\mem2[84][20] ), .QN(n31068) );
  SDFFX1 \mem2_reg[84][19]  ( .D(n11087), .SI(\mem2[84][18] ), .SE(test_se), 
        .CLK(n1996), .Q(\mem2[84][19] ), .QN(n31069) );
  SDFFX1 \mem2_reg[84][18]  ( .D(n11086), .SI(\mem2[84][17] ), .SE(test_se), 
        .CLK(n1996), .Q(\mem2[84][18] ), .QN(n31070) );
  SDFFX1 \mem2_reg[84][17]  ( .D(n11085), .SI(\mem2[84][16] ), .SE(test_se), 
        .CLK(n1997), .Q(\mem2[84][17] ), .QN(n31071) );
  SDFFX1 \mem2_reg[84][16]  ( .D(n11084), .SI(\mem2[83][23] ), .SE(test_se), 
        .CLK(n1997), .Q(\mem2[84][16] ), .QN(n31072) );
  SDFFX1 \mem2_reg[83][23]  ( .D(n11083), .SI(\mem2[83][22] ), .SE(test_se), 
        .CLK(n1997), .Q(\mem2[83][23] ), .QN(n31073) );
  SDFFX1 \mem2_reg[83][22]  ( .D(n11082), .SI(\mem2[83][21] ), .SE(test_se), 
        .CLK(n1997), .Q(\mem2[83][22] ), .QN(n31074) );
  SDFFX1 \mem2_reg[83][21]  ( .D(n11081), .SI(\mem2[83][20] ), .SE(test_se), 
        .CLK(n1997), .Q(\mem2[83][21] ), .QN(n31075) );
  SDFFX1 \mem2_reg[83][20]  ( .D(n11080), .SI(\mem2[83][19] ), .SE(test_se), 
        .CLK(n1997), .Q(\mem2[83][20] ), .QN(n31076) );
  SDFFX1 \mem2_reg[83][19]  ( .D(n11079), .SI(\mem2[83][18] ), .SE(test_se), 
        .CLK(n1997), .Q(\mem2[83][19] ), .QN(n31077) );
  SDFFX1 \mem2_reg[83][18]  ( .D(n11078), .SI(\mem2[83][17] ), .SE(test_se), 
        .CLK(n1997), .Q(\mem2[83][18] ), .QN(n31078) );
  SDFFX1 \mem2_reg[83][17]  ( .D(n11077), .SI(\mem2[83][16] ), .SE(test_se), 
        .CLK(n1997), .Q(\mem2[83][17] ), .QN(n31079) );
  SDFFX1 \mem2_reg[83][16]  ( .D(n11076), .SI(\mem2[82][23] ), .SE(test_se), 
        .CLK(n1997), .Q(\mem2[83][16] ), .QN(n31080) );
  SDFFX1 \mem2_reg[82][23]  ( .D(n11075), .SI(\mem2[82][22] ), .SE(test_se), 
        .CLK(n1997), .Q(\mem2[82][23] ), .QN(n31081) );
  SDFFX1 \mem2_reg[82][22]  ( .D(n11074), .SI(\mem2[82][21] ), .SE(test_se), 
        .CLK(n1997), .Q(\mem2[82][22] ), .QN(n31082) );
  SDFFX1 \mem2_reg[82][21]  ( .D(n11073), .SI(\mem2[82][20] ), .SE(test_se), 
        .CLK(n1998), .Q(\mem2[82][21] ), .QN(n31083) );
  SDFFX1 \mem2_reg[82][20]  ( .D(n11072), .SI(\mem2[82][19] ), .SE(test_se), 
        .CLK(n1998), .Q(\mem2[82][20] ), .QN(n31084) );
  SDFFX1 \mem2_reg[82][19]  ( .D(n11071), .SI(\mem2[82][18] ), .SE(test_se), 
        .CLK(n1998), .Q(\mem2[82][19] ), .QN(n31085) );
  SDFFX1 \mem2_reg[82][18]  ( .D(n11070), .SI(\mem2[82][17] ), .SE(test_se), 
        .CLK(n1998), .Q(\mem2[82][18] ), .QN(n31086) );
  SDFFX1 \mem2_reg[82][17]  ( .D(n11069), .SI(\mem2[82][16] ), .SE(test_se), 
        .CLK(n1998), .Q(\mem2[82][17] ), .QN(n31087) );
  SDFFX1 \mem2_reg[82][16]  ( .D(n11068), .SI(\mem2[81][23] ), .SE(test_se), 
        .CLK(n1998), .Q(\mem2[82][16] ), .QN(n31088) );
  SDFFX1 \mem2_reg[81][23]  ( .D(n11067), .SI(\mem2[81][22] ), .SE(test_se), 
        .CLK(n1998), .Q(\mem2[81][23] ), .QN(n31089) );
  SDFFX1 \mem2_reg[81][22]  ( .D(n11066), .SI(\mem2[81][21] ), .SE(test_se), 
        .CLK(n1998), .Q(\mem2[81][22] ), .QN(n31090) );
  SDFFX1 \mem2_reg[81][21]  ( .D(n11065), .SI(\mem2[81][20] ), .SE(test_se), 
        .CLK(n1998), .Q(\mem2[81][21] ), .QN(n31091) );
  SDFFX1 \mem2_reg[81][20]  ( .D(n11064), .SI(\mem2[81][19] ), .SE(test_se), 
        .CLK(n1998), .Q(\mem2[81][20] ), .QN(n31092) );
  SDFFX1 \mem2_reg[81][19]  ( .D(n11063), .SI(\mem2[81][18] ), .SE(test_se), 
        .CLK(n1998), .Q(\mem2[81][19] ), .QN(n31093) );
  SDFFX1 \mem2_reg[81][18]  ( .D(n11062), .SI(\mem2[81][17] ), .SE(test_se), 
        .CLK(n1998), .Q(\mem2[81][18] ), .QN(n31094) );
  SDFFX1 \mem2_reg[81][17]  ( .D(n11061), .SI(\mem2[81][16] ), .SE(test_se), 
        .CLK(n1999), .Q(\mem2[81][17] ), .QN(n31095) );
  SDFFX1 \mem2_reg[81][16]  ( .D(n11060), .SI(\mem2[80][23] ), .SE(test_se), 
        .CLK(n1999), .Q(\mem2[81][16] ), .QN(n31096) );
  SDFFX1 \mem2_reg[80][23]  ( .D(n11059), .SI(\mem2[80][22] ), .SE(test_se), 
        .CLK(n1999), .Q(\mem2[80][23] ), .QN(n31097) );
  SDFFX1 \mem2_reg[80][22]  ( .D(n11058), .SI(\mem2[80][21] ), .SE(test_se), 
        .CLK(n1999), .Q(\mem2[80][22] ), .QN(n31098) );
  SDFFX1 \mem2_reg[80][21]  ( .D(n11057), .SI(\mem2[80][20] ), .SE(test_se), 
        .CLK(n1999), .Q(\mem2[80][21] ), .QN(n31099) );
  SDFFX1 \mem2_reg[80][20]  ( .D(n11056), .SI(\mem2[80][19] ), .SE(test_se), 
        .CLK(n1999), .Q(\mem2[80][20] ), .QN(n31100) );
  SDFFX1 \mem2_reg[80][19]  ( .D(n11055), .SI(\mem2[80][18] ), .SE(test_se), 
        .CLK(n1999), .Q(\mem2[80][19] ), .QN(n31101) );
  SDFFX1 \mem2_reg[80][18]  ( .D(n11054), .SI(\mem2[80][17] ), .SE(test_se), 
        .CLK(n1999), .Q(\mem2[80][18] ), .QN(n31102) );
  SDFFX1 \mem2_reg[80][17]  ( .D(n11053), .SI(\mem2[80][16] ), .SE(test_se), 
        .CLK(n1999), .Q(\mem2[80][17] ), .QN(n31103) );
  SDFFX1 \mem2_reg[80][16]  ( .D(n11052), .SI(\mem2[79][23] ), .SE(test_se), 
        .CLK(n1999), .Q(\mem2[80][16] ), .QN(n31104) );
  SDFFX1 \mem2_reg[79][23]  ( .D(n11051), .SI(\mem2[79][22] ), .SE(test_se), 
        .CLK(n1999), .Q(\mem2[79][23] ), .QN(n31105) );
  SDFFX1 \mem2_reg[79][22]  ( .D(n11050), .SI(\mem2[79][21] ), .SE(test_se), 
        .CLK(n1999), .Q(\mem2[79][22] ), .QN(n31106) );
  SDFFX1 \mem2_reg[79][21]  ( .D(n11049), .SI(\mem2[79][20] ), .SE(test_se), 
        .CLK(n2000), .Q(\mem2[79][21] ), .QN(n31107) );
  SDFFX1 \mem2_reg[79][20]  ( .D(n11048), .SI(\mem2[79][19] ), .SE(test_se), 
        .CLK(n2000), .Q(\mem2[79][20] ), .QN(n31108) );
  SDFFX1 \mem2_reg[79][19]  ( .D(n11047), .SI(\mem2[79][18] ), .SE(test_se), 
        .CLK(n2000), .Q(\mem2[79][19] ), .QN(n31109) );
  SDFFX1 \mem2_reg[79][18]  ( .D(n11046), .SI(\mem2[79][17] ), .SE(test_se), 
        .CLK(n2000), .Q(\mem2[79][18] ), .QN(n31110) );
  SDFFX1 \mem2_reg[79][17]  ( .D(n11045), .SI(\mem2[79][16] ), .SE(test_se), 
        .CLK(n2000), .Q(\mem2[79][17] ), .QN(n31111) );
  SDFFX1 \mem2_reg[79][16]  ( .D(n11044), .SI(\mem2[78][23] ), .SE(test_se), 
        .CLK(n2000), .Q(\mem2[79][16] ), .QN(n31112) );
  SDFFX1 \mem2_reg[78][23]  ( .D(n11043), .SI(\mem2[78][22] ), .SE(test_se), 
        .CLK(n2000), .Q(\mem2[78][23] ), .QN(n31113) );
  SDFFX1 \mem2_reg[78][22]  ( .D(n11042), .SI(\mem2[78][21] ), .SE(test_se), 
        .CLK(n2000), .Q(\mem2[78][22] ), .QN(n31114) );
  SDFFX1 \mem2_reg[78][21]  ( .D(n11041), .SI(\mem2[78][20] ), .SE(test_se), 
        .CLK(n2000), .Q(\mem2[78][21] ), .QN(n31115) );
  SDFFX1 \mem2_reg[78][20]  ( .D(n11040), .SI(\mem2[78][19] ), .SE(test_se), 
        .CLK(n2000), .Q(\mem2[78][20] ), .QN(n31116) );
  SDFFX1 \mem2_reg[78][19]  ( .D(n11039), .SI(\mem2[78][18] ), .SE(test_se), 
        .CLK(n2000), .Q(\mem2[78][19] ), .QN(n31117) );
  SDFFX1 \mem2_reg[78][18]  ( .D(n11038), .SI(\mem2[78][17] ), .SE(test_se), 
        .CLK(n2000), .Q(\mem2[78][18] ), .QN(n31118) );
  SDFFX1 \mem2_reg[78][17]  ( .D(n11037), .SI(\mem2[78][16] ), .SE(test_se), 
        .CLK(n2001), .Q(\mem2[78][17] ), .QN(n31119) );
  SDFFX1 \mem2_reg[78][16]  ( .D(n11036), .SI(\mem2[77][23] ), .SE(test_se), 
        .CLK(n2001), .Q(\mem2[78][16] ), .QN(n31120) );
  SDFFX1 \mem2_reg[77][23]  ( .D(n11035), .SI(\mem2[77][22] ), .SE(test_se), 
        .CLK(n2001), .Q(\mem2[77][23] ), .QN(n31121) );
  SDFFX1 \mem2_reg[77][22]  ( .D(n11034), .SI(\mem2[77][21] ), .SE(test_se), 
        .CLK(n2001), .Q(\mem2[77][22] ), .QN(n31122) );
  SDFFX1 \mem2_reg[77][21]  ( .D(n11033), .SI(\mem2[77][20] ), .SE(test_se), 
        .CLK(n2001), .Q(\mem2[77][21] ), .QN(n31123) );
  SDFFX1 \mem2_reg[77][20]  ( .D(n11032), .SI(\mem2[77][19] ), .SE(test_se), 
        .CLK(n2001), .Q(\mem2[77][20] ), .QN(n31124) );
  SDFFX1 \mem2_reg[77][19]  ( .D(n11031), .SI(\mem2[77][18] ), .SE(test_se), 
        .CLK(n2001), .Q(\mem2[77][19] ), .QN(n31125) );
  SDFFX1 \mem2_reg[77][18]  ( .D(n11030), .SI(\mem2[77][17] ), .SE(test_se), 
        .CLK(n2001), .Q(\mem2[77][18] ), .QN(n31126) );
  SDFFX1 \mem2_reg[77][17]  ( .D(n11029), .SI(\mem2[77][16] ), .SE(test_se), 
        .CLK(n2001), .Q(\mem2[77][17] ), .QN(n31127) );
  SDFFX1 \mem2_reg[77][16]  ( .D(n11028), .SI(\mem2[76][23] ), .SE(test_se), 
        .CLK(n2001), .Q(\mem2[77][16] ), .QN(n31128) );
  SDFFX1 \mem2_reg[76][23]  ( .D(n11027), .SI(\mem2[76][22] ), .SE(test_se), 
        .CLK(n2001), .Q(\mem2[76][23] ), .QN(n31129) );
  SDFFX1 \mem2_reg[76][22]  ( .D(n11026), .SI(\mem2[76][21] ), .SE(test_se), 
        .CLK(n2001), .Q(\mem2[76][22] ), .QN(n31130) );
  SDFFX1 \mem2_reg[76][21]  ( .D(n11025), .SI(\mem2[76][20] ), .SE(test_se), 
        .CLK(n2002), .Q(\mem2[76][21] ), .QN(n31131) );
  SDFFX1 \mem2_reg[76][20]  ( .D(n11024), .SI(\mem2[76][19] ), .SE(test_se), 
        .CLK(n2002), .Q(\mem2[76][20] ), .QN(n31132) );
  SDFFX1 \mem2_reg[76][19]  ( .D(n11023), .SI(\mem2[76][18] ), .SE(test_se), 
        .CLK(n2002), .Q(\mem2[76][19] ), .QN(n31133) );
  SDFFX1 \mem2_reg[76][18]  ( .D(n11022), .SI(\mem2[76][17] ), .SE(test_se), 
        .CLK(n2002), .Q(\mem2[76][18] ), .QN(n31134) );
  SDFFX1 \mem2_reg[76][17]  ( .D(n11021), .SI(\mem2[76][16] ), .SE(test_se), 
        .CLK(n2002), .Q(\mem2[76][17] ), .QN(n31135) );
  SDFFX1 \mem2_reg[76][16]  ( .D(n11020), .SI(\mem2[75][23] ), .SE(test_se), 
        .CLK(n2002), .Q(\mem2[76][16] ), .QN(n31136) );
  SDFFX1 \mem2_reg[75][23]  ( .D(n11019), .SI(\mem2[75][22] ), .SE(test_se), 
        .CLK(n2002), .Q(\mem2[75][23] ), .QN(n31137) );
  SDFFX1 \mem2_reg[75][22]  ( .D(n11018), .SI(\mem2[75][21] ), .SE(test_se), 
        .CLK(n2002), .Q(\mem2[75][22] ), .QN(n31138) );
  SDFFX1 \mem2_reg[75][21]  ( .D(n11017), .SI(\mem2[75][20] ), .SE(test_se), 
        .CLK(n2002), .Q(\mem2[75][21] ), .QN(n31139) );
  SDFFX1 \mem2_reg[75][20]  ( .D(n11016), .SI(\mem2[75][19] ), .SE(test_se), 
        .CLK(n2002), .Q(\mem2[75][20] ), .QN(n31140) );
  SDFFX1 \mem2_reg[75][19]  ( .D(n11015), .SI(\mem2[75][18] ), .SE(test_se), 
        .CLK(n2002), .Q(\mem2[75][19] ), .QN(n31141) );
  SDFFX1 \mem2_reg[75][18]  ( .D(n11014), .SI(\mem2[75][17] ), .SE(test_se), 
        .CLK(n2002), .Q(\mem2[75][18] ), .QN(n31142) );
  SDFFX1 \mem2_reg[75][17]  ( .D(n11013), .SI(\mem2[75][16] ), .SE(test_se), 
        .CLK(n2003), .Q(\mem2[75][17] ), .QN(n31143) );
  SDFFX1 \mem2_reg[75][16]  ( .D(n11012), .SI(\mem2[74][23] ), .SE(test_se), 
        .CLK(n2003), .Q(\mem2[75][16] ), .QN(n31144) );
  SDFFX1 \mem2_reg[74][23]  ( .D(n11011), .SI(\mem2[74][22] ), .SE(test_se), 
        .CLK(n2003), .Q(\mem2[74][23] ), .QN(n31145) );
  SDFFX1 \mem2_reg[74][22]  ( .D(n11010), .SI(\mem2[74][21] ), .SE(test_se), 
        .CLK(n2003), .Q(\mem2[74][22] ), .QN(n31146) );
  SDFFX1 \mem2_reg[74][21]  ( .D(n11009), .SI(\mem2[74][20] ), .SE(test_se), 
        .CLK(n2003), .Q(\mem2[74][21] ), .QN(n31147) );
  SDFFX1 \mem2_reg[74][20]  ( .D(n11008), .SI(\mem2[74][19] ), .SE(test_se), 
        .CLK(n2003), .Q(\mem2[74][20] ), .QN(n31148) );
  SDFFX1 \mem2_reg[74][19]  ( .D(n11007), .SI(\mem2[74][18] ), .SE(test_se), 
        .CLK(n2003), .Q(\mem2[74][19] ), .QN(n31149) );
  SDFFX1 \mem2_reg[74][18]  ( .D(n11006), .SI(\mem2[74][17] ), .SE(test_se), 
        .CLK(n2003), .Q(\mem2[74][18] ), .QN(n31150) );
  SDFFX1 \mem2_reg[74][17]  ( .D(n11005), .SI(\mem2[74][16] ), .SE(test_se), 
        .CLK(n2003), .Q(\mem2[74][17] ), .QN(n31151) );
  SDFFX1 \mem2_reg[74][16]  ( .D(n11004), .SI(\mem2[73][23] ), .SE(test_se), 
        .CLK(n2003), .Q(\mem2[74][16] ), .QN(n31152) );
  SDFFX1 \mem2_reg[73][23]  ( .D(n11003), .SI(\mem2[73][22] ), .SE(test_se), 
        .CLK(n2003), .Q(\mem2[73][23] ), .QN(n31153) );
  SDFFX1 \mem2_reg[73][22]  ( .D(n11002), .SI(\mem2[73][21] ), .SE(test_se), 
        .CLK(n2003), .Q(\mem2[73][22] ), .QN(n31154) );
  SDFFX1 \mem2_reg[73][21]  ( .D(n11001), .SI(\mem2[73][20] ), .SE(test_se), 
        .CLK(n2004), .Q(\mem2[73][21] ), .QN(n31155) );
  SDFFX1 \mem2_reg[73][20]  ( .D(n11000), .SI(\mem2[73][19] ), .SE(test_se), 
        .CLK(n2004), .Q(\mem2[73][20] ), .QN(n31156) );
  SDFFX1 \mem2_reg[73][19]  ( .D(n10999), .SI(\mem2[73][18] ), .SE(test_se), 
        .CLK(n2004), .Q(\mem2[73][19] ), .QN(n31157) );
  SDFFX1 \mem2_reg[73][18]  ( .D(n10998), .SI(\mem2[73][17] ), .SE(test_se), 
        .CLK(n2004), .Q(\mem2[73][18] ), .QN(n31158) );
  SDFFX1 \mem2_reg[73][17]  ( .D(n10997), .SI(\mem2[73][16] ), .SE(test_se), 
        .CLK(n2004), .Q(\mem2[73][17] ), .QN(n31159) );
  SDFFX1 \mem2_reg[73][16]  ( .D(n10996), .SI(\mem2[72][23] ), .SE(test_se), 
        .CLK(n2004), .Q(\mem2[73][16] ), .QN(n31160) );
  SDFFX1 \mem2_reg[72][23]  ( .D(n10995), .SI(\mem2[72][22] ), .SE(test_se), 
        .CLK(n2004), .Q(\mem2[72][23] ), .QN(n31161) );
  SDFFX1 \mem2_reg[72][22]  ( .D(n10994), .SI(\mem2[72][21] ), .SE(test_se), 
        .CLK(n2004), .Q(\mem2[72][22] ), .QN(n31162) );
  SDFFX1 \mem2_reg[72][21]  ( .D(n10993), .SI(\mem2[72][20] ), .SE(test_se), 
        .CLK(n2004), .Q(\mem2[72][21] ), .QN(n31163) );
  SDFFX1 \mem2_reg[72][20]  ( .D(n10992), .SI(\mem2[72][19] ), .SE(test_se), 
        .CLK(n2004), .Q(\mem2[72][20] ), .QN(n31164) );
  SDFFX1 \mem2_reg[72][19]  ( .D(n10991), .SI(\mem2[72][18] ), .SE(test_se), 
        .CLK(n2004), .Q(\mem2[72][19] ), .QN(n31165) );
  SDFFX1 \mem2_reg[72][18]  ( .D(n10990), .SI(\mem2[72][17] ), .SE(test_se), 
        .CLK(n2004), .Q(\mem2[72][18] ), .QN(n31166) );
  SDFFX1 \mem2_reg[72][17]  ( .D(n10989), .SI(\mem2[72][16] ), .SE(test_se), 
        .CLK(n2005), .Q(\mem2[72][17] ), .QN(n31167) );
  SDFFX1 \mem2_reg[72][16]  ( .D(n10988), .SI(\mem2[71][23] ), .SE(test_se), 
        .CLK(n2005), .Q(\mem2[72][16] ), .QN(n31168) );
  SDFFX1 \mem2_reg[71][23]  ( .D(n10987), .SI(\mem2[71][22] ), .SE(test_se), 
        .CLK(n2005), .Q(\mem2[71][23] ), .QN(n31169) );
  SDFFX1 \mem2_reg[71][22]  ( .D(n10986), .SI(\mem2[71][21] ), .SE(test_se), 
        .CLK(n2005), .Q(\mem2[71][22] ), .QN(n31170) );
  SDFFX1 \mem2_reg[71][21]  ( .D(n10985), .SI(\mem2[71][20] ), .SE(test_se), 
        .CLK(n2005), .Q(\mem2[71][21] ), .QN(n31171) );
  SDFFX1 \mem2_reg[71][20]  ( .D(n10984), .SI(\mem2[71][19] ), .SE(test_se), 
        .CLK(n2005), .Q(\mem2[71][20] ), .QN(n31172) );
  SDFFX1 \mem2_reg[71][19]  ( .D(n10983), .SI(\mem2[71][18] ), .SE(test_se), 
        .CLK(n2005), .Q(\mem2[71][19] ), .QN(n31173) );
  SDFFX1 \mem2_reg[71][18]  ( .D(n10982), .SI(\mem2[71][17] ), .SE(test_se), 
        .CLK(n2005), .Q(\mem2[71][18] ), .QN(n31174) );
  SDFFX1 \mem2_reg[71][17]  ( .D(n10981), .SI(\mem2[71][16] ), .SE(test_se), 
        .CLK(n2005), .Q(\mem2[71][17] ), .QN(n31175) );
  SDFFX1 \mem2_reg[71][16]  ( .D(n10980), .SI(\mem2[70][23] ), .SE(test_se), 
        .CLK(n2005), .Q(\mem2[71][16] ), .QN(n31176) );
  SDFFX1 \mem2_reg[70][23]  ( .D(n10979), .SI(\mem2[70][22] ), .SE(test_se), 
        .CLK(n2005), .Q(\mem2[70][23] ), .QN(n31177) );
  SDFFX1 \mem2_reg[70][22]  ( .D(n10978), .SI(\mem2[70][21] ), .SE(test_se), 
        .CLK(n2005), .Q(\mem2[70][22] ), .QN(n31178) );
  SDFFX1 \mem2_reg[70][21]  ( .D(n10977), .SI(\mem2[70][20] ), .SE(test_se), 
        .CLK(n2006), .Q(\mem2[70][21] ), .QN(n31179) );
  SDFFX1 \mem2_reg[70][20]  ( .D(n10976), .SI(\mem2[70][19] ), .SE(test_se), 
        .CLK(n2006), .Q(\mem2[70][20] ), .QN(n31180) );
  SDFFX1 \mem2_reg[70][19]  ( .D(n10975), .SI(\mem2[70][18] ), .SE(test_se), 
        .CLK(n2006), .Q(\mem2[70][19] ), .QN(n31181) );
  SDFFX1 \mem2_reg[70][18]  ( .D(n10974), .SI(\mem2[70][17] ), .SE(test_se), 
        .CLK(n2006), .Q(\mem2[70][18] ), .QN(n31182) );
  SDFFX1 \mem2_reg[70][17]  ( .D(n10973), .SI(\mem2[70][16] ), .SE(test_se), 
        .CLK(n2006), .Q(\mem2[70][17] ), .QN(n31183) );
  SDFFX1 \mem2_reg[70][16]  ( .D(n10972), .SI(\mem2[69][23] ), .SE(test_se), 
        .CLK(n2006), .Q(\mem2[70][16] ), .QN(n31184) );
  SDFFX1 \mem2_reg[69][23]  ( .D(n10971), .SI(\mem2[69][22] ), .SE(test_se), 
        .CLK(n2006), .Q(\mem2[69][23] ), .QN(n31185) );
  SDFFX1 \mem2_reg[69][22]  ( .D(n10970), .SI(\mem2[69][21] ), .SE(test_se), 
        .CLK(n2006), .Q(\mem2[69][22] ), .QN(n31186) );
  SDFFX1 \mem2_reg[69][21]  ( .D(n10969), .SI(\mem2[69][20] ), .SE(test_se), 
        .CLK(n2006), .Q(\mem2[69][21] ), .QN(n31187) );
  SDFFX1 \mem2_reg[69][20]  ( .D(n10968), .SI(\mem2[69][19] ), .SE(test_se), 
        .CLK(n2006), .Q(\mem2[69][20] ), .QN(n31188) );
  SDFFX1 \mem2_reg[69][19]  ( .D(n10967), .SI(\mem2[69][18] ), .SE(test_se), 
        .CLK(n2006), .Q(\mem2[69][19] ), .QN(n31189) );
  SDFFX1 \mem2_reg[69][18]  ( .D(n10966), .SI(\mem2[69][17] ), .SE(test_se), 
        .CLK(n2006), .Q(\mem2[69][18] ), .QN(n31190) );
  SDFFX1 \mem2_reg[69][17]  ( .D(n10965), .SI(\mem2[69][16] ), .SE(test_se), 
        .CLK(n2007), .Q(\mem2[69][17] ), .QN(n31191) );
  SDFFX1 \mem2_reg[69][16]  ( .D(n10964), .SI(\mem2[68][23] ), .SE(test_se), 
        .CLK(n2007), .Q(\mem2[69][16] ), .QN(n31192) );
  SDFFX1 \mem2_reg[68][23]  ( .D(n10963), .SI(\mem2[68][22] ), .SE(test_se), 
        .CLK(n2007), .Q(\mem2[68][23] ), .QN(n31193) );
  SDFFX1 \mem2_reg[68][22]  ( .D(n10962), .SI(\mem2[68][21] ), .SE(test_se), 
        .CLK(n2007), .Q(\mem2[68][22] ), .QN(n31194) );
  SDFFX1 \mem2_reg[68][21]  ( .D(n10961), .SI(\mem2[68][20] ), .SE(test_se), 
        .CLK(n2007), .Q(\mem2[68][21] ), .QN(n31195) );
  SDFFX1 \mem2_reg[68][20]  ( .D(n10960), .SI(\mem2[68][19] ), .SE(test_se), 
        .CLK(n2007), .Q(\mem2[68][20] ), .QN(n31196) );
  SDFFX1 \mem2_reg[68][19]  ( .D(n10959), .SI(\mem2[68][18] ), .SE(test_se), 
        .CLK(n2007), .Q(\mem2[68][19] ), .QN(n31197) );
  SDFFX1 \mem2_reg[68][18]  ( .D(n10958), .SI(\mem2[68][17] ), .SE(test_se), 
        .CLK(n2007), .Q(\mem2[68][18] ), .QN(n31198) );
  SDFFX1 \mem2_reg[68][17]  ( .D(n10957), .SI(\mem2[68][16] ), .SE(test_se), 
        .CLK(n2007), .Q(\mem2[68][17] ), .QN(n31199) );
  SDFFX1 \mem2_reg[68][16]  ( .D(n10956), .SI(\mem2[67][23] ), .SE(test_se), 
        .CLK(n2007), .Q(\mem2[68][16] ), .QN(n31200) );
  SDFFX1 \mem2_reg[67][23]  ( .D(n10955), .SI(\mem2[67][22] ), .SE(test_se), 
        .CLK(n2007), .Q(\mem2[67][23] ), .QN(n31201) );
  SDFFX1 \mem2_reg[67][22]  ( .D(n10954), .SI(\mem2[67][21] ), .SE(test_se), 
        .CLK(n2007), .Q(\mem2[67][22] ), .QN(n31202) );
  SDFFX1 \mem2_reg[67][21]  ( .D(n10953), .SI(\mem2[67][20] ), .SE(test_se), 
        .CLK(n2008), .Q(\mem2[67][21] ), .QN(n31203) );
  SDFFX1 \mem2_reg[67][20]  ( .D(n10952), .SI(\mem2[67][19] ), .SE(test_se), 
        .CLK(n2008), .Q(\mem2[67][20] ), .QN(n31204) );
  SDFFX1 \mem2_reg[67][19]  ( .D(n10951), .SI(\mem2[67][18] ), .SE(test_se), 
        .CLK(n2008), .Q(\mem2[67][19] ), .QN(n31205) );
  SDFFX1 \mem2_reg[67][18]  ( .D(n10950), .SI(\mem2[67][17] ), .SE(test_se), 
        .CLK(n2008), .Q(\mem2[67][18] ), .QN(n31206) );
  SDFFX1 \mem2_reg[67][17]  ( .D(n10949), .SI(\mem2[67][16] ), .SE(test_se), 
        .CLK(n2008), .Q(\mem2[67][17] ), .QN(n31207) );
  SDFFX1 \mem2_reg[67][16]  ( .D(n10948), .SI(\mem2[66][23] ), .SE(test_se), 
        .CLK(n2008), .Q(\mem2[67][16] ), .QN(n31208) );
  SDFFX1 \mem2_reg[66][23]  ( .D(n10947), .SI(\mem2[66][22] ), .SE(test_se), 
        .CLK(n2008), .Q(\mem2[66][23] ), .QN(n31209) );
  SDFFX1 \mem2_reg[66][22]  ( .D(n10946), .SI(\mem2[66][21] ), .SE(test_se), 
        .CLK(n2008), .Q(\mem2[66][22] ), .QN(n31210) );
  SDFFX1 \mem2_reg[66][21]  ( .D(n10945), .SI(\mem2[66][20] ), .SE(test_se), 
        .CLK(n2008), .Q(\mem2[66][21] ), .QN(n31211) );
  SDFFX1 \mem2_reg[66][20]  ( .D(n10944), .SI(\mem2[66][19] ), .SE(test_se), 
        .CLK(n2008), .Q(\mem2[66][20] ), .QN(n31212) );
  SDFFX1 \mem2_reg[66][19]  ( .D(n10943), .SI(\mem2[66][18] ), .SE(test_se), 
        .CLK(n2008), .Q(\mem2[66][19] ), .QN(n31213) );
  SDFFX1 \mem2_reg[66][18]  ( .D(n10942), .SI(\mem2[66][17] ), .SE(test_se), 
        .CLK(n2008), .Q(\mem2[66][18] ), .QN(n31214) );
  SDFFX1 \mem2_reg[66][17]  ( .D(n10941), .SI(\mem2[66][16] ), .SE(test_se), 
        .CLK(n2009), .Q(\mem2[66][17] ), .QN(n31215) );
  SDFFX1 \mem2_reg[66][16]  ( .D(n10940), .SI(\mem2[65][23] ), .SE(test_se), 
        .CLK(n2009), .Q(\mem2[66][16] ), .QN(n31216) );
  SDFFX1 \mem2_reg[65][23]  ( .D(n10939), .SI(\mem2[65][22] ), .SE(test_se), 
        .CLK(n2009), .Q(\mem2[65][23] ), .QN(n31217) );
  SDFFX1 \mem2_reg[65][22]  ( .D(n10938), .SI(\mem2[65][21] ), .SE(test_se), 
        .CLK(n2009), .Q(\mem2[65][22] ), .QN(n31218) );
  SDFFX1 \mem2_reg[65][21]  ( .D(n10937), .SI(\mem2[65][20] ), .SE(test_se), 
        .CLK(n2009), .Q(\mem2[65][21] ), .QN(n31219) );
  SDFFX1 \mem2_reg[65][20]  ( .D(n10936), .SI(\mem2[65][19] ), .SE(test_se), 
        .CLK(n2009), .Q(\mem2[65][20] ), .QN(n31220) );
  SDFFX1 \mem2_reg[65][19]  ( .D(n10935), .SI(\mem2[65][18] ), .SE(test_se), 
        .CLK(n2009), .Q(\mem2[65][19] ), .QN(n31221) );
  SDFFX1 \mem2_reg[65][18]  ( .D(n10934), .SI(\mem2[65][17] ), .SE(test_se), 
        .CLK(n2009), .Q(\mem2[65][18] ), .QN(n31222) );
  SDFFX1 \mem2_reg[65][17]  ( .D(n10933), .SI(\mem2[65][16] ), .SE(test_se), 
        .CLK(n2009), .Q(\mem2[65][17] ), .QN(n31223) );
  SDFFX1 \mem2_reg[65][16]  ( .D(n10932), .SI(\mem2[64][23] ), .SE(test_se), 
        .CLK(n2009), .Q(\mem2[65][16] ), .QN(n31224) );
  SDFFX1 \mem2_reg[64][23]  ( .D(n10931), .SI(\mem2[64][22] ), .SE(test_se), 
        .CLK(n2009), .Q(\mem2[64][23] ), .QN(n31225) );
  SDFFX1 \mem2_reg[64][22]  ( .D(n10930), .SI(\mem2[64][21] ), .SE(test_se), 
        .CLK(n2009), .Q(\mem2[64][22] ), .QN(n31226) );
  SDFFX1 \mem2_reg[64][21]  ( .D(n10929), .SI(\mem2[64][20] ), .SE(test_se), 
        .CLK(n2010), .Q(\mem2[64][21] ), .QN(n31227) );
  SDFFX1 \mem2_reg[64][20]  ( .D(n10928), .SI(\mem2[64][19] ), .SE(test_se), 
        .CLK(n2010), .Q(\mem2[64][20] ), .QN(n31228) );
  SDFFX1 \mem2_reg[64][19]  ( .D(n10927), .SI(\mem2[64][18] ), .SE(test_se), 
        .CLK(n2010), .Q(\mem2[64][19] ), .QN(n31229) );
  SDFFX1 \mem2_reg[64][18]  ( .D(n10926), .SI(\mem2[64][17] ), .SE(test_se), 
        .CLK(n2010), .Q(\mem2[64][18] ), .QN(n31230) );
  SDFFX1 \mem2_reg[64][17]  ( .D(n10925), .SI(\mem2[64][16] ), .SE(test_se), 
        .CLK(n2010), .Q(\mem2[64][17] ), .QN(n31231) );
  SDFFX1 \mem2_reg[64][16]  ( .D(n10924), .SI(\mem2[63][23] ), .SE(test_se), 
        .CLK(n2010), .Q(\mem2[64][16] ), .QN(n31232) );
  SDFFX1 \mem2_reg[63][23]  ( .D(n10923), .SI(\mem2[63][22] ), .SE(test_se), 
        .CLK(n2010), .Q(\mem2[63][23] ), .QN(n31233) );
  SDFFX1 \mem2_reg[63][22]  ( .D(n10922), .SI(\mem2[63][21] ), .SE(test_se), 
        .CLK(n2010), .Q(\mem2[63][22] ), .QN(n31234) );
  SDFFX1 \mem2_reg[63][21]  ( .D(n10921), .SI(\mem2[63][20] ), .SE(test_se), 
        .CLK(n2010), .Q(\mem2[63][21] ), .QN(n31235) );
  SDFFX1 \mem2_reg[63][20]  ( .D(n10920), .SI(\mem2[63][19] ), .SE(test_se), 
        .CLK(n2010), .Q(\mem2[63][20] ), .QN(n31236) );
  SDFFX1 \mem2_reg[63][19]  ( .D(n10919), .SI(\mem2[63][18] ), .SE(test_se), 
        .CLK(n2010), .Q(\mem2[63][19] ), .QN(n31237) );
  SDFFX1 \mem2_reg[63][18]  ( .D(n10918), .SI(\mem2[63][17] ), .SE(test_se), 
        .CLK(n2010), .Q(\mem2[63][18] ), .QN(n31238) );
  SDFFX1 \mem2_reg[63][17]  ( .D(n10917), .SI(\mem2[63][16] ), .SE(test_se), 
        .CLK(n2011), .Q(\mem2[63][17] ), .QN(n31239) );
  SDFFX1 \mem2_reg[63][16]  ( .D(n10916), .SI(\mem2[62][23] ), .SE(test_se), 
        .CLK(n2011), .Q(\mem2[63][16] ), .QN(n31240) );
  SDFFX1 \mem2_reg[62][23]  ( .D(n10915), .SI(\mem2[62][22] ), .SE(test_se), 
        .CLK(n2011), .Q(\mem2[62][23] ), .QN(n31241) );
  SDFFX1 \mem2_reg[62][22]  ( .D(n10914), .SI(\mem2[62][21] ), .SE(test_se), 
        .CLK(n2011), .Q(\mem2[62][22] ), .QN(n31242) );
  SDFFX1 \mem2_reg[62][21]  ( .D(n10913), .SI(\mem2[62][20] ), .SE(test_se), 
        .CLK(n2011), .Q(\mem2[62][21] ), .QN(n31243) );
  SDFFX1 \mem2_reg[62][20]  ( .D(n10912), .SI(\mem2[62][19] ), .SE(test_se), 
        .CLK(n2011), .Q(\mem2[62][20] ), .QN(n31244) );
  SDFFX1 \mem2_reg[62][19]  ( .D(n10911), .SI(\mem2[62][18] ), .SE(test_se), 
        .CLK(n2011), .Q(\mem2[62][19] ), .QN(n31245) );
  SDFFX1 \mem2_reg[62][18]  ( .D(n10910), .SI(\mem2[62][17] ), .SE(test_se), 
        .CLK(n2011), .Q(\mem2[62][18] ), .QN(n31246) );
  SDFFX1 \mem2_reg[62][17]  ( .D(n10909), .SI(\mem2[62][16] ), .SE(test_se), 
        .CLK(n2011), .Q(\mem2[62][17] ), .QN(n31247) );
  SDFFX1 \mem2_reg[62][16]  ( .D(n10908), .SI(\mem2[61][23] ), .SE(test_se), 
        .CLK(n2011), .Q(\mem2[62][16] ), .QN(n31248) );
  SDFFX1 \mem2_reg[61][23]  ( .D(n10907), .SI(\mem2[61][22] ), .SE(test_se), 
        .CLK(n2011), .Q(\mem2[61][23] ), .QN(n31249) );
  SDFFX1 \mem2_reg[61][22]  ( .D(n10906), .SI(\mem2[61][21] ), .SE(test_se), 
        .CLK(n2011), .Q(\mem2[61][22] ), .QN(n31250) );
  SDFFX1 \mem2_reg[61][21]  ( .D(n10905), .SI(\mem2[61][20] ), .SE(test_se), 
        .CLK(n2012), .Q(\mem2[61][21] ), .QN(n31251) );
  SDFFX1 \mem2_reg[61][20]  ( .D(n10904), .SI(\mem2[61][19] ), .SE(test_se), 
        .CLK(n2012), .Q(\mem2[61][20] ), .QN(n31252) );
  SDFFX1 \mem2_reg[61][19]  ( .D(n10903), .SI(\mem2[61][18] ), .SE(test_se), 
        .CLK(n2012), .Q(\mem2[61][19] ), .QN(n31253) );
  SDFFX1 \mem2_reg[61][18]  ( .D(n10902), .SI(\mem2[61][17] ), .SE(test_se), 
        .CLK(n2012), .Q(\mem2[61][18] ), .QN(n31254) );
  SDFFX1 \mem2_reg[61][17]  ( .D(n10901), .SI(\mem2[61][16] ), .SE(test_se), 
        .CLK(n2012), .Q(\mem2[61][17] ), .QN(n31255) );
  SDFFX1 \mem2_reg[61][16]  ( .D(n10900), .SI(\mem2[60][23] ), .SE(test_se), 
        .CLK(n2012), .Q(\mem2[61][16] ), .QN(n31256) );
  SDFFX1 \mem2_reg[60][23]  ( .D(n10899), .SI(\mem2[60][22] ), .SE(test_se), 
        .CLK(n2012), .Q(\mem2[60][23] ), .QN(n31257) );
  SDFFX1 \mem2_reg[60][22]  ( .D(n10898), .SI(\mem2[60][21] ), .SE(test_se), 
        .CLK(n2012), .Q(\mem2[60][22] ), .QN(n31258) );
  SDFFX1 \mem2_reg[60][21]  ( .D(n10897), .SI(\mem2[60][20] ), .SE(test_se), 
        .CLK(n2012), .Q(\mem2[60][21] ), .QN(n31259) );
  SDFFX1 \mem2_reg[60][20]  ( .D(n10896), .SI(\mem2[60][19] ), .SE(test_se), 
        .CLK(n2012), .Q(\mem2[60][20] ), .QN(n31260) );
  SDFFX1 \mem2_reg[60][19]  ( .D(n10895), .SI(\mem2[60][18] ), .SE(test_se), 
        .CLK(n2012), .Q(\mem2[60][19] ), .QN(n31261) );
  SDFFX1 \mem2_reg[60][18]  ( .D(n10894), .SI(\mem2[60][17] ), .SE(test_se), 
        .CLK(n2012), .Q(\mem2[60][18] ), .QN(n31262) );
  SDFFX1 \mem2_reg[60][17]  ( .D(n10893), .SI(\mem2[60][16] ), .SE(test_se), 
        .CLK(n2013), .Q(\mem2[60][17] ), .QN(n31263) );
  SDFFX1 \mem2_reg[60][16]  ( .D(n10892), .SI(\mem2[59][23] ), .SE(test_se), 
        .CLK(n2013), .Q(\mem2[60][16] ), .QN(n31264) );
  SDFFX1 \mem2_reg[59][23]  ( .D(n10891), .SI(\mem2[59][22] ), .SE(test_se), 
        .CLK(n2013), .Q(\mem2[59][23] ), .QN(n31265) );
  SDFFX1 \mem2_reg[59][22]  ( .D(n10890), .SI(\mem2[59][21] ), .SE(test_se), 
        .CLK(n2013), .Q(\mem2[59][22] ), .QN(n31266) );
  SDFFX1 \mem2_reg[59][21]  ( .D(n10889), .SI(\mem2[59][20] ), .SE(test_se), 
        .CLK(n2013), .Q(\mem2[59][21] ), .QN(n31267) );
  SDFFX1 \mem2_reg[59][20]  ( .D(n10888), .SI(\mem2[59][19] ), .SE(test_se), 
        .CLK(n2013), .Q(\mem2[59][20] ), .QN(n31268) );
  SDFFX1 \mem2_reg[59][19]  ( .D(n10887), .SI(\mem2[59][18] ), .SE(test_se), 
        .CLK(n2013), .Q(\mem2[59][19] ), .QN(n31269) );
  SDFFX1 \mem2_reg[59][18]  ( .D(n10886), .SI(\mem2[59][17] ), .SE(test_se), 
        .CLK(n2013), .Q(\mem2[59][18] ), .QN(n31270) );
  SDFFX1 \mem2_reg[59][17]  ( .D(n10885), .SI(\mem2[59][16] ), .SE(test_se), 
        .CLK(n2013), .Q(\mem2[59][17] ), .QN(n31271) );
  SDFFX1 \mem2_reg[59][16]  ( .D(n10884), .SI(\mem2[58][23] ), .SE(test_se), 
        .CLK(n2013), .Q(\mem2[59][16] ), .QN(n31272) );
  SDFFX1 \mem2_reg[58][23]  ( .D(n10883), .SI(\mem2[58][22] ), .SE(test_se), 
        .CLK(n2013), .Q(\mem2[58][23] ), .QN(n31273) );
  SDFFX1 \mem2_reg[58][22]  ( .D(n10882), .SI(\mem2[58][21] ), .SE(test_se), 
        .CLK(n2013), .Q(\mem2[58][22] ), .QN(n31274) );
  SDFFX1 \mem2_reg[58][21]  ( .D(n10881), .SI(\mem2[58][20] ), .SE(test_se), 
        .CLK(n2014), .Q(\mem2[58][21] ), .QN(n31275) );
  SDFFX1 \mem2_reg[58][20]  ( .D(n10880), .SI(\mem2[58][19] ), .SE(test_se), 
        .CLK(n2014), .Q(\mem2[58][20] ), .QN(n31276) );
  SDFFX1 \mem2_reg[58][19]  ( .D(n10879), .SI(\mem2[58][18] ), .SE(test_se), 
        .CLK(n2014), .Q(\mem2[58][19] ), .QN(n31277) );
  SDFFX1 \mem2_reg[58][18]  ( .D(n10878), .SI(\mem2[58][17] ), .SE(test_se), 
        .CLK(n2014), .Q(\mem2[58][18] ), .QN(n31278) );
  SDFFX1 \mem2_reg[58][17]  ( .D(n10877), .SI(\mem2[58][16] ), .SE(test_se), 
        .CLK(n2014), .Q(\mem2[58][17] ), .QN(n31279) );
  SDFFX1 \mem2_reg[58][16]  ( .D(n10876), .SI(\mem2[57][23] ), .SE(test_se), 
        .CLK(n2014), .Q(\mem2[58][16] ), .QN(n31280) );
  SDFFX1 \mem2_reg[57][23]  ( .D(n10875), .SI(\mem2[57][22] ), .SE(test_se), 
        .CLK(n2014), .Q(\mem2[57][23] ), .QN(n31281) );
  SDFFX1 \mem2_reg[57][22]  ( .D(n10874), .SI(\mem2[57][21] ), .SE(test_se), 
        .CLK(n2014), .Q(\mem2[57][22] ), .QN(n31282) );
  SDFFX1 \mem2_reg[57][21]  ( .D(n10873), .SI(\mem2[57][20] ), .SE(test_se), 
        .CLK(n2014), .Q(\mem2[57][21] ), .QN(n31283) );
  SDFFX1 \mem2_reg[57][20]  ( .D(n10872), .SI(\mem2[57][19] ), .SE(test_se), 
        .CLK(n2014), .Q(\mem2[57][20] ), .QN(n31284) );
  SDFFX1 \mem2_reg[57][19]  ( .D(n10871), .SI(\mem2[57][18] ), .SE(test_se), 
        .CLK(n2014), .Q(\mem2[57][19] ), .QN(n31285) );
  SDFFX1 \mem2_reg[57][18]  ( .D(n10870), .SI(\mem2[57][17] ), .SE(test_se), 
        .CLK(n2014), .Q(\mem2[57][18] ), .QN(n31286) );
  SDFFX1 \mem2_reg[57][17]  ( .D(n10869), .SI(\mem2[57][16] ), .SE(test_se), 
        .CLK(n2015), .Q(\mem2[57][17] ), .QN(n31287) );
  SDFFX1 \mem2_reg[57][16]  ( .D(n10868), .SI(\mem2[56][23] ), .SE(test_se), 
        .CLK(n2015), .Q(\mem2[57][16] ), .QN(n31288) );
  SDFFX1 \mem2_reg[56][23]  ( .D(n10867), .SI(\mem2[56][22] ), .SE(test_se), 
        .CLK(n2015), .Q(\mem2[56][23] ), .QN(n31289) );
  SDFFX1 \mem2_reg[56][22]  ( .D(n10866), .SI(\mem2[56][21] ), .SE(test_se), 
        .CLK(n2015), .Q(\mem2[56][22] ), .QN(n31290) );
  SDFFX1 \mem2_reg[56][21]  ( .D(n10865), .SI(\mem2[56][20] ), .SE(test_se), 
        .CLK(n2015), .Q(\mem2[56][21] ), .QN(n31291) );
  SDFFX1 \mem2_reg[56][20]  ( .D(n10864), .SI(\mem2[56][19] ), .SE(test_se), 
        .CLK(n2015), .Q(\mem2[56][20] ), .QN(n31292) );
  SDFFX1 \mem2_reg[56][19]  ( .D(n10863), .SI(\mem2[56][18] ), .SE(test_se), 
        .CLK(n2015), .Q(\mem2[56][19] ), .QN(n31293) );
  SDFFX1 \mem2_reg[56][18]  ( .D(n10862), .SI(\mem2[56][17] ), .SE(test_se), 
        .CLK(n2015), .Q(\mem2[56][18] ), .QN(n31294) );
  SDFFX1 \mem2_reg[56][17]  ( .D(n10861), .SI(\mem2[56][16] ), .SE(test_se), 
        .CLK(n2015), .Q(\mem2[56][17] ), .QN(n31295) );
  SDFFX1 \mem2_reg[56][16]  ( .D(n10860), .SI(\mem2[55][23] ), .SE(test_se), 
        .CLK(n2015), .Q(\mem2[56][16] ), .QN(n31296) );
  SDFFX1 \mem2_reg[55][23]  ( .D(n10859), .SI(\mem2[55][22] ), .SE(test_se), 
        .CLK(n2015), .Q(\mem2[55][23] ), .QN(n31297) );
  SDFFX1 \mem2_reg[55][22]  ( .D(n10858), .SI(\mem2[55][21] ), .SE(test_se), 
        .CLK(n2015), .Q(\mem2[55][22] ), .QN(n31298) );
  SDFFX1 \mem2_reg[55][21]  ( .D(n10857), .SI(\mem2[55][20] ), .SE(test_se), 
        .CLK(n2016), .Q(\mem2[55][21] ), .QN(n31299) );
  SDFFX1 \mem2_reg[55][20]  ( .D(n10856), .SI(\mem2[55][19] ), .SE(test_se), 
        .CLK(n2016), .Q(\mem2[55][20] ), .QN(n31300) );
  SDFFX1 \mem2_reg[55][19]  ( .D(n10855), .SI(\mem2[55][18] ), .SE(test_se), 
        .CLK(n2016), .Q(\mem2[55][19] ), .QN(n31301) );
  SDFFX1 \mem2_reg[55][18]  ( .D(n10854), .SI(\mem2[55][17] ), .SE(test_se), 
        .CLK(n2016), .Q(\mem2[55][18] ), .QN(n31302) );
  SDFFX1 \mem2_reg[55][17]  ( .D(n10853), .SI(\mem2[55][16] ), .SE(test_se), 
        .CLK(n2016), .Q(\mem2[55][17] ), .QN(n31303) );
  SDFFX1 \mem2_reg[55][16]  ( .D(n10852), .SI(\mem2[54][23] ), .SE(test_se), 
        .CLK(n2016), .Q(\mem2[55][16] ), .QN(n31304) );
  SDFFX1 \mem2_reg[54][23]  ( .D(n10851), .SI(\mem2[54][22] ), .SE(test_se), 
        .CLK(n2016), .Q(\mem2[54][23] ), .QN(n31305) );
  SDFFX1 \mem2_reg[54][22]  ( .D(n10850), .SI(\mem2[54][21] ), .SE(test_se), 
        .CLK(n2016), .Q(\mem2[54][22] ), .QN(n31306) );
  SDFFX1 \mem2_reg[54][21]  ( .D(n10849), .SI(\mem2[54][20] ), .SE(test_se), 
        .CLK(n2016), .Q(\mem2[54][21] ), .QN(n31307) );
  SDFFX1 \mem2_reg[54][20]  ( .D(n10848), .SI(\mem2[54][19] ), .SE(test_se), 
        .CLK(n2016), .Q(\mem2[54][20] ), .QN(n31308) );
  SDFFX1 \mem2_reg[54][19]  ( .D(n10847), .SI(\mem2[54][18] ), .SE(test_se), 
        .CLK(n2016), .Q(\mem2[54][19] ), .QN(n31309) );
  SDFFX1 \mem2_reg[54][18]  ( .D(n10846), .SI(\mem2[54][17] ), .SE(test_se), 
        .CLK(n2016), .Q(\mem2[54][18] ), .QN(n31310) );
  SDFFX1 \mem2_reg[54][17]  ( .D(n10845), .SI(\mem2[54][16] ), .SE(test_se), 
        .CLK(n2017), .Q(\mem2[54][17] ), .QN(n31311) );
  SDFFX1 \mem2_reg[54][16]  ( .D(n10844), .SI(\mem2[53][23] ), .SE(test_se), 
        .CLK(n2017), .Q(\mem2[54][16] ), .QN(n31312) );
  SDFFX1 \mem2_reg[53][23]  ( .D(n10843), .SI(\mem2[53][22] ), .SE(test_se), 
        .CLK(n2017), .Q(\mem2[53][23] ), .QN(n31313) );
  SDFFX1 \mem2_reg[53][22]  ( .D(n10842), .SI(\mem2[53][21] ), .SE(test_se), 
        .CLK(n2017), .Q(\mem2[53][22] ), .QN(n31314) );
  SDFFX1 \mem2_reg[53][21]  ( .D(n10841), .SI(\mem2[53][20] ), .SE(test_se), 
        .CLK(n2017), .Q(\mem2[53][21] ), .QN(n31315) );
  SDFFX1 \mem2_reg[53][20]  ( .D(n10840), .SI(\mem2[53][19] ), .SE(test_se), 
        .CLK(n2017), .Q(\mem2[53][20] ), .QN(n31316) );
  SDFFX1 \mem2_reg[53][19]  ( .D(n10839), .SI(\mem2[53][18] ), .SE(test_se), 
        .CLK(n2017), .Q(\mem2[53][19] ), .QN(n31317) );
  SDFFX1 \mem2_reg[53][18]  ( .D(n10838), .SI(\mem2[53][17] ), .SE(test_se), 
        .CLK(n2017), .Q(\mem2[53][18] ), .QN(n31318) );
  SDFFX1 \mem2_reg[53][17]  ( .D(n10837), .SI(\mem2[53][16] ), .SE(test_se), 
        .CLK(n2017), .Q(\mem2[53][17] ), .QN(n31319) );
  SDFFX1 \mem2_reg[53][16]  ( .D(n10836), .SI(\mem2[52][23] ), .SE(test_se), 
        .CLK(n2017), .Q(\mem2[53][16] ), .QN(n31320) );
  SDFFX1 \mem2_reg[52][23]  ( .D(n10835), .SI(\mem2[52][22] ), .SE(test_se), 
        .CLK(n2017), .Q(\mem2[52][23] ), .QN(n31321) );
  SDFFX1 \mem2_reg[52][22]  ( .D(n10834), .SI(\mem2[52][21] ), .SE(test_se), 
        .CLK(n2017), .Q(\mem2[52][22] ), .QN(n31322) );
  SDFFX1 \mem2_reg[52][21]  ( .D(n10833), .SI(\mem2[52][20] ), .SE(test_se), 
        .CLK(n2018), .Q(\mem2[52][21] ), .QN(n31323) );
  SDFFX1 \mem2_reg[52][20]  ( .D(n10832), .SI(\mem2[52][19] ), .SE(test_se), 
        .CLK(n2018), .Q(\mem2[52][20] ), .QN(n31324) );
  SDFFX1 \mem2_reg[52][19]  ( .D(n10831), .SI(\mem2[52][18] ), .SE(test_se), 
        .CLK(n2018), .Q(\mem2[52][19] ), .QN(n31325) );
  SDFFX1 \mem2_reg[52][18]  ( .D(n10830), .SI(\mem2[52][17] ), .SE(test_se), 
        .CLK(n2018), .Q(\mem2[52][18] ), .QN(n31326) );
  SDFFX1 \mem2_reg[52][17]  ( .D(n10829), .SI(\mem2[52][16] ), .SE(test_se), 
        .CLK(n2018), .Q(\mem2[52][17] ), .QN(n31327) );
  SDFFX1 \mem2_reg[52][16]  ( .D(n10828), .SI(\mem2[51][23] ), .SE(test_se), 
        .CLK(n2018), .Q(\mem2[52][16] ), .QN(n31328) );
  SDFFX1 \mem2_reg[51][23]  ( .D(n10827), .SI(\mem2[51][22] ), .SE(test_se), 
        .CLK(n2018), .Q(\mem2[51][23] ), .QN(n31329) );
  SDFFX1 \mem2_reg[51][22]  ( .D(n10826), .SI(\mem2[51][21] ), .SE(test_se), 
        .CLK(n2018), .Q(\mem2[51][22] ), .QN(n31330) );
  SDFFX1 \mem2_reg[51][21]  ( .D(n10825), .SI(\mem2[51][20] ), .SE(test_se), 
        .CLK(n2018), .Q(\mem2[51][21] ), .QN(n31331) );
  SDFFX1 \mem2_reg[51][20]  ( .D(n10824), .SI(\mem2[51][19] ), .SE(test_se), 
        .CLK(n2018), .Q(\mem2[51][20] ), .QN(n31332) );
  SDFFX1 \mem2_reg[51][19]  ( .D(n10823), .SI(\mem2[51][18] ), .SE(test_se), 
        .CLK(n2018), .Q(\mem2[51][19] ), .QN(n31333) );
  SDFFX1 \mem2_reg[51][18]  ( .D(n10822), .SI(\mem2[51][17] ), .SE(test_se), 
        .CLK(n2018), .Q(\mem2[51][18] ), .QN(n31334) );
  SDFFX1 \mem2_reg[51][17]  ( .D(n10821), .SI(\mem2[51][16] ), .SE(test_se), 
        .CLK(n2019), .Q(\mem2[51][17] ), .QN(n31335) );
  SDFFX1 \mem2_reg[51][16]  ( .D(n10820), .SI(\mem2[50][23] ), .SE(test_se), 
        .CLK(n2019), .Q(\mem2[51][16] ), .QN(n31336) );
  SDFFX1 \mem2_reg[50][23]  ( .D(n10819), .SI(\mem2[50][22] ), .SE(test_se), 
        .CLK(n2019), .Q(\mem2[50][23] ), .QN(n31337) );
  SDFFX1 \mem2_reg[50][22]  ( .D(n10818), .SI(\mem2[50][21] ), .SE(test_se), 
        .CLK(n2019), .Q(\mem2[50][22] ), .QN(n31338) );
  SDFFX1 \mem2_reg[50][21]  ( .D(n10817), .SI(\mem2[50][20] ), .SE(test_se), 
        .CLK(n2019), .Q(\mem2[50][21] ), .QN(n31339) );
  SDFFX1 \mem2_reg[50][20]  ( .D(n10816), .SI(\mem2[50][19] ), .SE(test_se), 
        .CLK(n2019), .Q(\mem2[50][20] ), .QN(n31340) );
  SDFFX1 \mem2_reg[50][19]  ( .D(n10815), .SI(\mem2[50][18] ), .SE(test_se), 
        .CLK(n2019), .Q(\mem2[50][19] ), .QN(n31341) );
  SDFFX1 \mem2_reg[50][18]  ( .D(n10814), .SI(\mem2[50][17] ), .SE(test_se), 
        .CLK(n2019), .Q(\mem2[50][18] ), .QN(n31342) );
  SDFFX1 \mem2_reg[50][17]  ( .D(n10813), .SI(\mem2[50][16] ), .SE(test_se), 
        .CLK(n2019), .Q(\mem2[50][17] ), .QN(n31343) );
  SDFFX1 \mem2_reg[50][16]  ( .D(n10812), .SI(\mem2[49][23] ), .SE(test_se), 
        .CLK(n2019), .Q(\mem2[50][16] ), .QN(n31344) );
  SDFFX1 \mem2_reg[49][23]  ( .D(n10811), .SI(\mem2[49][22] ), .SE(test_se), 
        .CLK(n2019), .Q(\mem2[49][23] ), .QN(n31345) );
  SDFFX1 \mem2_reg[49][22]  ( .D(n10810), .SI(\mem2[49][21] ), .SE(test_se), 
        .CLK(n2019), .Q(\mem2[49][22] ), .QN(n31346) );
  SDFFX1 \mem2_reg[49][21]  ( .D(n10809), .SI(\mem2[49][20] ), .SE(test_se), 
        .CLK(n2020), .Q(\mem2[49][21] ), .QN(n31347) );
  SDFFX1 \mem2_reg[49][20]  ( .D(n10808), .SI(\mem2[49][19] ), .SE(test_se), 
        .CLK(n2020), .Q(\mem2[49][20] ), .QN(n31348) );
  SDFFX1 \mem2_reg[49][19]  ( .D(n10807), .SI(\mem2[49][18] ), .SE(test_se), 
        .CLK(n2020), .Q(\mem2[49][19] ), .QN(n31349) );
  SDFFX1 \mem2_reg[49][18]  ( .D(n10806), .SI(\mem2[49][17] ), .SE(test_se), 
        .CLK(n2020), .Q(\mem2[49][18] ), .QN(n31350) );
  SDFFX1 \mem2_reg[49][17]  ( .D(n10805), .SI(\mem2[49][16] ), .SE(test_se), 
        .CLK(n2020), .Q(\mem2[49][17] ), .QN(n31351) );
  SDFFX1 \mem2_reg[49][16]  ( .D(n10804), .SI(\mem2[48][23] ), .SE(test_se), 
        .CLK(n2020), .Q(\mem2[49][16] ), .QN(n31352) );
  SDFFX1 \mem2_reg[48][23]  ( .D(n10803), .SI(\mem2[48][22] ), .SE(test_se), 
        .CLK(n2020), .Q(\mem2[48][23] ), .QN(n31353) );
  SDFFX1 \mem2_reg[48][22]  ( .D(n10802), .SI(\mem2[48][21] ), .SE(test_se), 
        .CLK(n2020), .Q(\mem2[48][22] ), .QN(n31354) );
  SDFFX1 \mem2_reg[48][21]  ( .D(n10801), .SI(\mem2[48][20] ), .SE(test_se), 
        .CLK(n2020), .Q(\mem2[48][21] ), .QN(n31355) );
  SDFFX1 \mem2_reg[48][20]  ( .D(n10800), .SI(\mem2[48][19] ), .SE(test_se), 
        .CLK(n2020), .Q(\mem2[48][20] ), .QN(n31356) );
  SDFFX1 \mem2_reg[48][19]  ( .D(n10799), .SI(\mem2[48][18] ), .SE(test_se), 
        .CLK(n2020), .Q(\mem2[48][19] ), .QN(n31357) );
  SDFFX1 \mem2_reg[48][18]  ( .D(n10798), .SI(\mem2[48][17] ), .SE(test_se), 
        .CLK(n2020), .Q(\mem2[48][18] ), .QN(n31358) );
  SDFFX1 \mem2_reg[48][17]  ( .D(n10797), .SI(\mem2[48][16] ), .SE(test_se), 
        .CLK(n2021), .Q(\mem2[48][17] ), .QN(n31359) );
  SDFFX1 \mem2_reg[48][16]  ( .D(n10796), .SI(\mem2[47][23] ), .SE(test_se), 
        .CLK(n2021), .Q(\mem2[48][16] ), .QN(n31360) );
  SDFFX1 \mem2_reg[47][23]  ( .D(n10795), .SI(\mem2[47][22] ), .SE(test_se), 
        .CLK(n2021), .Q(\mem2[47][23] ), .QN(n31361) );
  SDFFX1 \mem2_reg[47][22]  ( .D(n10794), .SI(\mem2[47][21] ), .SE(test_se), 
        .CLK(n2021), .Q(\mem2[47][22] ), .QN(n31362) );
  SDFFX1 \mem2_reg[47][21]  ( .D(n10793), .SI(\mem2[47][20] ), .SE(test_se), 
        .CLK(n2021), .Q(\mem2[47][21] ), .QN(n31363) );
  SDFFX1 \mem2_reg[47][20]  ( .D(n10792), .SI(\mem2[47][19] ), .SE(test_se), 
        .CLK(n2021), .Q(\mem2[47][20] ), .QN(n31364) );
  SDFFX1 \mem2_reg[47][19]  ( .D(n10791), .SI(\mem2[47][18] ), .SE(test_se), 
        .CLK(n2021), .Q(\mem2[47][19] ), .QN(n31365) );
  SDFFX1 \mem2_reg[47][18]  ( .D(n10790), .SI(\mem2[47][17] ), .SE(test_se), 
        .CLK(n2021), .Q(\mem2[47][18] ), .QN(n31366) );
  SDFFX1 \mem2_reg[47][17]  ( .D(n10789), .SI(\mem2[47][16] ), .SE(test_se), 
        .CLK(n2021), .Q(\mem2[47][17] ), .QN(n31367) );
  SDFFX1 \mem2_reg[47][16]  ( .D(n10788), .SI(\mem2[46][23] ), .SE(test_se), 
        .CLK(n2021), .Q(\mem2[47][16] ), .QN(n31368) );
  SDFFX1 \mem2_reg[46][23]  ( .D(n10787), .SI(\mem2[46][22] ), .SE(test_se), 
        .CLK(n2021), .Q(\mem2[46][23] ), .QN(n31369) );
  SDFFX1 \mem2_reg[46][22]  ( .D(n10786), .SI(\mem2[46][21] ), .SE(test_se), 
        .CLK(n2021), .Q(\mem2[46][22] ), .QN(n31370) );
  SDFFX1 \mem2_reg[46][21]  ( .D(n10785), .SI(\mem2[46][20] ), .SE(test_se), 
        .CLK(n2022), .Q(\mem2[46][21] ), .QN(n31371) );
  SDFFX1 \mem2_reg[46][20]  ( .D(n10784), .SI(\mem2[46][19] ), .SE(test_se), 
        .CLK(n2022), .Q(\mem2[46][20] ), .QN(n31372) );
  SDFFX1 \mem2_reg[46][19]  ( .D(n10783), .SI(\mem2[46][18] ), .SE(test_se), 
        .CLK(n2022), .Q(\mem2[46][19] ), .QN(n31373) );
  SDFFX1 \mem2_reg[46][18]  ( .D(n10782), .SI(\mem2[46][17] ), .SE(test_se), 
        .CLK(n2022), .Q(\mem2[46][18] ), .QN(n31374) );
  SDFFX1 \mem2_reg[46][17]  ( .D(n10781), .SI(\mem2[46][16] ), .SE(test_se), 
        .CLK(n2022), .Q(\mem2[46][17] ), .QN(n31375) );
  SDFFX1 \mem2_reg[46][16]  ( .D(n10780), .SI(\mem2[45][23] ), .SE(test_se), 
        .CLK(n2022), .Q(\mem2[46][16] ), .QN(n31376) );
  SDFFX1 \mem2_reg[45][23]  ( .D(n10779), .SI(\mem2[45][22] ), .SE(test_se), 
        .CLK(n2022), .Q(\mem2[45][23] ), .QN(n31377) );
  SDFFX1 \mem2_reg[45][22]  ( .D(n10778), .SI(\mem2[45][21] ), .SE(test_se), 
        .CLK(n2022), .Q(\mem2[45][22] ), .QN(n31378) );
  SDFFX1 \mem2_reg[45][21]  ( .D(n10777), .SI(\mem2[45][20] ), .SE(test_se), 
        .CLK(n2022), .Q(\mem2[45][21] ), .QN(n31379) );
  SDFFX1 \mem2_reg[45][20]  ( .D(n10776), .SI(\mem2[45][19] ), .SE(test_se), 
        .CLK(n2022), .Q(\mem2[45][20] ), .QN(n31380) );
  SDFFX1 \mem2_reg[45][19]  ( .D(n10775), .SI(\mem2[45][18] ), .SE(test_se), 
        .CLK(n2022), .Q(\mem2[45][19] ), .QN(n31381) );
  SDFFX1 \mem2_reg[45][18]  ( .D(n10774), .SI(\mem2[45][17] ), .SE(test_se), 
        .CLK(n2022), .Q(\mem2[45][18] ), .QN(n31382) );
  SDFFX1 \mem2_reg[45][17]  ( .D(n10773), .SI(\mem2[45][16] ), .SE(test_se), 
        .CLK(n2023), .Q(\mem2[45][17] ), .QN(n31383) );
  SDFFX1 \mem2_reg[45][16]  ( .D(n10772), .SI(\mem2[44][23] ), .SE(test_se), 
        .CLK(n2023), .Q(\mem2[45][16] ), .QN(n31384) );
  SDFFX1 \mem2_reg[44][23]  ( .D(n10771), .SI(\mem2[44][22] ), .SE(test_se), 
        .CLK(n2023), .Q(\mem2[44][23] ), .QN(n31385) );
  SDFFX1 \mem2_reg[44][22]  ( .D(n10770), .SI(\mem2[44][21] ), .SE(test_se), 
        .CLK(n2023), .Q(\mem2[44][22] ), .QN(n31386) );
  SDFFX1 \mem2_reg[44][21]  ( .D(n10769), .SI(\mem2[44][20] ), .SE(test_se), 
        .CLK(n2023), .Q(\mem2[44][21] ), .QN(n31387) );
  SDFFX1 \mem2_reg[44][20]  ( .D(n10768), .SI(\mem2[44][19] ), .SE(test_se), 
        .CLK(n2023), .Q(\mem2[44][20] ), .QN(n31388) );
  SDFFX1 \mem2_reg[44][19]  ( .D(n10767), .SI(\mem2[44][18] ), .SE(test_se), 
        .CLK(n2023), .Q(\mem2[44][19] ), .QN(n31389) );
  SDFFX1 \mem2_reg[44][18]  ( .D(n10766), .SI(\mem2[44][17] ), .SE(test_se), 
        .CLK(n2023), .Q(\mem2[44][18] ), .QN(n31390) );
  SDFFX1 \mem2_reg[44][17]  ( .D(n10765), .SI(\mem2[44][16] ), .SE(test_se), 
        .CLK(n2023), .Q(\mem2[44][17] ), .QN(n31391) );
  SDFFX1 \mem2_reg[44][16]  ( .D(n10764), .SI(\mem2[43][23] ), .SE(test_se), 
        .CLK(n2023), .Q(\mem2[44][16] ), .QN(n31392) );
  SDFFX1 \mem2_reg[43][23]  ( .D(n10763), .SI(\mem2[43][22] ), .SE(test_se), 
        .CLK(n2023), .Q(\mem2[43][23] ), .QN(n31393) );
  SDFFX1 \mem2_reg[43][22]  ( .D(n10762), .SI(\mem2[43][21] ), .SE(test_se), 
        .CLK(n2023), .Q(\mem2[43][22] ), .QN(n31394) );
  SDFFX1 \mem2_reg[43][21]  ( .D(n10761), .SI(\mem2[43][20] ), .SE(test_se), 
        .CLK(n2024), .Q(\mem2[43][21] ), .QN(n31395) );
  SDFFX1 \mem2_reg[43][20]  ( .D(n10760), .SI(\mem2[43][19] ), .SE(test_se), 
        .CLK(n2024), .Q(\mem2[43][20] ), .QN(n31396) );
  SDFFX1 \mem2_reg[43][19]  ( .D(n10759), .SI(\mem2[43][18] ), .SE(test_se), 
        .CLK(n2024), .Q(\mem2[43][19] ), .QN(n31397) );
  SDFFX1 \mem2_reg[43][18]  ( .D(n10758), .SI(\mem2[43][17] ), .SE(test_se), 
        .CLK(n2024), .Q(\mem2[43][18] ), .QN(n31398) );
  SDFFX1 \mem2_reg[43][17]  ( .D(n10757), .SI(\mem2[43][16] ), .SE(test_se), 
        .CLK(n2024), .Q(\mem2[43][17] ), .QN(n31399) );
  SDFFX1 \mem2_reg[43][16]  ( .D(n10756), .SI(\mem2[42][23] ), .SE(test_se), 
        .CLK(n2024), .Q(\mem2[43][16] ), .QN(n31400) );
  SDFFX1 \mem2_reg[42][23]  ( .D(n10755), .SI(\mem2[42][22] ), .SE(test_se), 
        .CLK(n2024), .Q(\mem2[42][23] ), .QN(n31401) );
  SDFFX1 \mem2_reg[42][22]  ( .D(n10754), .SI(\mem2[42][21] ), .SE(test_se), 
        .CLK(n2024), .Q(\mem2[42][22] ), .QN(n31402) );
  SDFFX1 \mem2_reg[42][21]  ( .D(n10753), .SI(\mem2[42][20] ), .SE(test_se), 
        .CLK(n2024), .Q(\mem2[42][21] ), .QN(n31403) );
  SDFFX1 \mem2_reg[42][20]  ( .D(n10752), .SI(\mem2[42][19] ), .SE(test_se), 
        .CLK(n2024), .Q(\mem2[42][20] ), .QN(n31404) );
  SDFFX1 \mem2_reg[42][19]  ( .D(n10751), .SI(\mem2[42][18] ), .SE(test_se), 
        .CLK(n2024), .Q(\mem2[42][19] ), .QN(n31405) );
  SDFFX1 \mem2_reg[42][18]  ( .D(n10750), .SI(\mem2[42][17] ), .SE(test_se), 
        .CLK(n2024), .Q(\mem2[42][18] ), .QN(n31406) );
  SDFFX1 \mem2_reg[42][17]  ( .D(n10749), .SI(\mem2[42][16] ), .SE(test_se), 
        .CLK(n2025), .Q(\mem2[42][17] ), .QN(n31407) );
  SDFFX1 \mem2_reg[42][16]  ( .D(n10748), .SI(\mem2[41][23] ), .SE(test_se), 
        .CLK(n2025), .Q(\mem2[42][16] ), .QN(n31408) );
  SDFFX1 \mem2_reg[41][23]  ( .D(n10747), .SI(\mem2[41][22] ), .SE(test_se), 
        .CLK(n2025), .Q(\mem2[41][23] ), .QN(n31409) );
  SDFFX1 \mem2_reg[41][22]  ( .D(n10746), .SI(\mem2[41][21] ), .SE(test_se), 
        .CLK(n2025), .Q(\mem2[41][22] ), .QN(n31410) );
  SDFFX1 \mem2_reg[41][21]  ( .D(n10745), .SI(\mem2[41][20] ), .SE(test_se), 
        .CLK(n2025), .Q(\mem2[41][21] ), .QN(n31411) );
  SDFFX1 \mem2_reg[41][20]  ( .D(n10744), .SI(\mem2[41][19] ), .SE(test_se), 
        .CLK(n2025), .Q(\mem2[41][20] ), .QN(n31412) );
  SDFFX1 \mem2_reg[41][19]  ( .D(n10743), .SI(\mem2[41][18] ), .SE(test_se), 
        .CLK(n2025), .Q(\mem2[41][19] ), .QN(n31413) );
  SDFFX1 \mem2_reg[41][18]  ( .D(n10742), .SI(\mem2[41][17] ), .SE(test_se), 
        .CLK(n2025), .Q(\mem2[41][18] ), .QN(n31414) );
  SDFFX1 \mem2_reg[41][17]  ( .D(n10741), .SI(\mem2[41][16] ), .SE(test_se), 
        .CLK(n2025), .Q(\mem2[41][17] ), .QN(n31415) );
  SDFFX1 \mem2_reg[41][16]  ( .D(n10740), .SI(\mem2[40][23] ), .SE(test_se), 
        .CLK(n2025), .Q(\mem2[41][16] ), .QN(n31416) );
  SDFFX1 \mem2_reg[40][23]  ( .D(n10739), .SI(\mem2[40][22] ), .SE(test_se), 
        .CLK(n2025), .Q(\mem2[40][23] ), .QN(n31417) );
  SDFFX1 \mem2_reg[40][22]  ( .D(n10738), .SI(\mem2[40][21] ), .SE(test_se), 
        .CLK(n2025), .Q(\mem2[40][22] ), .QN(n31418) );
  SDFFX1 \mem2_reg[40][21]  ( .D(n10737), .SI(\mem2[40][20] ), .SE(test_se), 
        .CLK(n2026), .Q(\mem2[40][21] ), .QN(n31419) );
  SDFFX1 \mem2_reg[40][20]  ( .D(n10736), .SI(\mem2[40][19] ), .SE(test_se), 
        .CLK(n2026), .Q(\mem2[40][20] ), .QN(n31420) );
  SDFFX1 \mem2_reg[40][19]  ( .D(n10735), .SI(\mem2[40][18] ), .SE(test_se), 
        .CLK(n2026), .Q(\mem2[40][19] ), .QN(n31421) );
  SDFFX1 \mem2_reg[40][18]  ( .D(n10734), .SI(\mem2[40][17] ), .SE(test_se), 
        .CLK(n2026), .Q(\mem2[40][18] ), .QN(n31422) );
  SDFFX1 \mem2_reg[40][17]  ( .D(n10733), .SI(\mem2[40][16] ), .SE(test_se), 
        .CLK(n2026), .Q(\mem2[40][17] ), .QN(n31423) );
  SDFFX1 \mem2_reg[40][16]  ( .D(n10732), .SI(\mem2[39][23] ), .SE(test_se), 
        .CLK(n2026), .Q(\mem2[40][16] ), .QN(n31424) );
  SDFFX1 \mem2_reg[39][23]  ( .D(n10731), .SI(\mem2[39][22] ), .SE(test_se), 
        .CLK(n2026), .Q(\mem2[39][23] ), .QN(n31425) );
  SDFFX1 \mem2_reg[39][22]  ( .D(n10730), .SI(\mem2[39][21] ), .SE(test_se), 
        .CLK(n2026), .Q(\mem2[39][22] ), .QN(n31426) );
  SDFFX1 \mem2_reg[39][21]  ( .D(n10729), .SI(\mem2[39][20] ), .SE(test_se), 
        .CLK(n2026), .Q(\mem2[39][21] ), .QN(n31427) );
  SDFFX1 \mem2_reg[39][20]  ( .D(n10728), .SI(\mem2[39][19] ), .SE(test_se), 
        .CLK(n2026), .Q(\mem2[39][20] ), .QN(n31428) );
  SDFFX1 \mem2_reg[39][19]  ( .D(n10727), .SI(\mem2[39][18] ), .SE(test_se), 
        .CLK(n2026), .Q(\mem2[39][19] ), .QN(n31429) );
  SDFFX1 \mem2_reg[39][18]  ( .D(n10726), .SI(\mem2[39][17] ), .SE(test_se), 
        .CLK(n2026), .Q(\mem2[39][18] ), .QN(n31430) );
  SDFFX1 \mem2_reg[39][17]  ( .D(n10725), .SI(\mem2[39][16] ), .SE(test_se), 
        .CLK(n2027), .Q(\mem2[39][17] ), .QN(n31431) );
  SDFFX1 \mem2_reg[39][16]  ( .D(n10724), .SI(\mem2[38][23] ), .SE(test_se), 
        .CLK(n2027), .Q(\mem2[39][16] ), .QN(n31432) );
  SDFFX1 \mem2_reg[38][23]  ( .D(n10723), .SI(\mem2[38][22] ), .SE(test_se), 
        .CLK(n2027), .Q(\mem2[38][23] ), .QN(n31433) );
  SDFFX1 \mem2_reg[38][22]  ( .D(n10722), .SI(\mem2[38][21] ), .SE(test_se), 
        .CLK(n2027), .Q(\mem2[38][22] ), .QN(n31434) );
  SDFFX1 \mem2_reg[38][21]  ( .D(n10721), .SI(\mem2[38][20] ), .SE(test_se), 
        .CLK(n2027), .Q(\mem2[38][21] ), .QN(n31435) );
  SDFFX1 \mem2_reg[38][20]  ( .D(n10720), .SI(\mem2[38][19] ), .SE(test_se), 
        .CLK(n2027), .Q(\mem2[38][20] ), .QN(n31436) );
  SDFFX1 \mem2_reg[38][19]  ( .D(n10719), .SI(\mem2[38][18] ), .SE(test_se), 
        .CLK(n2027), .Q(\mem2[38][19] ), .QN(n31437) );
  SDFFX1 \mem2_reg[38][18]  ( .D(n10718), .SI(\mem2[38][17] ), .SE(test_se), 
        .CLK(n2027), .Q(\mem2[38][18] ), .QN(n31438) );
  SDFFX1 \mem2_reg[38][17]  ( .D(n10717), .SI(\mem2[38][16] ), .SE(test_se), 
        .CLK(n2027), .Q(\mem2[38][17] ), .QN(n31439) );
  SDFFX1 \mem2_reg[38][16]  ( .D(n10716), .SI(\mem2[37][23] ), .SE(test_se), 
        .CLK(n2027), .Q(\mem2[38][16] ), .QN(n31440) );
  SDFFX1 \mem2_reg[37][23]  ( .D(n10715), .SI(\mem2[37][22] ), .SE(test_se), 
        .CLK(n2027), .Q(\mem2[37][23] ), .QN(n31441) );
  SDFFX1 \mem2_reg[37][22]  ( .D(n10714), .SI(\mem2[37][21] ), .SE(test_se), 
        .CLK(n2027), .Q(\mem2[37][22] ), .QN(n31442) );
  SDFFX1 \mem2_reg[37][21]  ( .D(n10713), .SI(\mem2[37][20] ), .SE(test_se), 
        .CLK(n2028), .Q(\mem2[37][21] ), .QN(n31443) );
  SDFFX1 \mem2_reg[37][20]  ( .D(n10712), .SI(\mem2[37][19] ), .SE(test_se), 
        .CLK(n2028), .Q(\mem2[37][20] ), .QN(n31444) );
  SDFFX1 \mem2_reg[37][19]  ( .D(n10711), .SI(\mem2[37][18] ), .SE(test_se), 
        .CLK(n2028), .Q(\mem2[37][19] ), .QN(n31445) );
  SDFFX1 \mem2_reg[37][18]  ( .D(n10710), .SI(\mem2[37][17] ), .SE(test_se), 
        .CLK(n2028), .Q(\mem2[37][18] ), .QN(n31446) );
  SDFFX1 \mem2_reg[37][17]  ( .D(n10709), .SI(\mem2[37][16] ), .SE(test_se), 
        .CLK(n2028), .Q(\mem2[37][17] ), .QN(n31447) );
  SDFFX1 \mem2_reg[37][16]  ( .D(n10708), .SI(\mem2[36][23] ), .SE(test_se), 
        .CLK(n2028), .Q(\mem2[37][16] ), .QN(n31448) );
  SDFFX1 \mem2_reg[36][23]  ( .D(n10707), .SI(\mem2[36][22] ), .SE(test_se), 
        .CLK(n2028), .Q(\mem2[36][23] ), .QN(n31449) );
  SDFFX1 \mem2_reg[36][22]  ( .D(n10706), .SI(\mem2[36][21] ), .SE(test_se), 
        .CLK(n2028), .Q(\mem2[36][22] ), .QN(n31450) );
  SDFFX1 \mem2_reg[36][21]  ( .D(n10705), .SI(\mem2[36][20] ), .SE(test_se), 
        .CLK(n2028), .Q(\mem2[36][21] ), .QN(n31451) );
  SDFFX1 \mem2_reg[36][20]  ( .D(n10704), .SI(\mem2[36][19] ), .SE(test_se), 
        .CLK(n2028), .Q(\mem2[36][20] ), .QN(n31452) );
  SDFFX1 \mem2_reg[36][19]  ( .D(n10703), .SI(\mem2[36][18] ), .SE(test_se), 
        .CLK(n2028), .Q(\mem2[36][19] ), .QN(n31453) );
  SDFFX1 \mem2_reg[36][18]  ( .D(n10702), .SI(\mem2[36][17] ), .SE(test_se), 
        .CLK(n2028), .Q(\mem2[36][18] ), .QN(n31454) );
  SDFFX1 \mem2_reg[36][17]  ( .D(n10701), .SI(\mem2[36][16] ), .SE(test_se), 
        .CLK(n2029), .Q(\mem2[36][17] ), .QN(n31455) );
  SDFFX1 \mem2_reg[36][16]  ( .D(n10700), .SI(\mem2[35][23] ), .SE(test_se), 
        .CLK(n2029), .Q(\mem2[36][16] ), .QN(n31456) );
  SDFFX1 \mem2_reg[35][23]  ( .D(n10699), .SI(\mem2[35][22] ), .SE(test_se), 
        .CLK(n2029), .Q(\mem2[35][23] ), .QN(n31457) );
  SDFFX1 \mem2_reg[35][22]  ( .D(n10698), .SI(\mem2[35][21] ), .SE(test_se), 
        .CLK(n2029), .Q(\mem2[35][22] ), .QN(n31458) );
  SDFFX1 \mem2_reg[35][21]  ( .D(n10697), .SI(\mem2[35][20] ), .SE(test_se), 
        .CLK(n2029), .Q(\mem2[35][21] ), .QN(n31459) );
  SDFFX1 \mem2_reg[35][20]  ( .D(n10696), .SI(\mem2[35][19] ), .SE(test_se), 
        .CLK(n2029), .Q(\mem2[35][20] ), .QN(n31460) );
  SDFFX1 \mem2_reg[35][19]  ( .D(n10695), .SI(\mem2[35][18] ), .SE(test_se), 
        .CLK(n2029), .Q(\mem2[35][19] ), .QN(n31461) );
  SDFFX1 \mem2_reg[35][18]  ( .D(n10694), .SI(\mem2[35][17] ), .SE(test_se), 
        .CLK(n2029), .Q(\mem2[35][18] ), .QN(n31462) );
  SDFFX1 \mem2_reg[35][17]  ( .D(n10693), .SI(\mem2[35][16] ), .SE(test_se), 
        .CLK(n2029), .Q(\mem2[35][17] ), .QN(n31463) );
  SDFFX1 \mem2_reg[35][16]  ( .D(n10692), .SI(\mem2[34][23] ), .SE(test_se), 
        .CLK(n2029), .Q(\mem2[35][16] ), .QN(n31464) );
  SDFFX1 \mem2_reg[34][23]  ( .D(n10691), .SI(\mem2[34][22] ), .SE(test_se), 
        .CLK(n2029), .Q(\mem2[34][23] ), .QN(n31465) );
  SDFFX1 \mem2_reg[34][22]  ( .D(n10690), .SI(\mem2[34][21] ), .SE(test_se), 
        .CLK(n2029), .Q(\mem2[34][22] ), .QN(n31466) );
  SDFFX1 \mem2_reg[34][21]  ( .D(n10689), .SI(\mem2[34][20] ), .SE(test_se), 
        .CLK(n2030), .Q(\mem2[34][21] ), .QN(n31467) );
  SDFFX1 \mem2_reg[34][20]  ( .D(n10688), .SI(\mem2[34][19] ), .SE(test_se), 
        .CLK(n2030), .Q(\mem2[34][20] ), .QN(n31468) );
  SDFFX1 \mem2_reg[34][19]  ( .D(n10687), .SI(\mem2[34][18] ), .SE(test_se), 
        .CLK(n2030), .Q(\mem2[34][19] ), .QN(n31469) );
  SDFFX1 \mem2_reg[34][18]  ( .D(n10686), .SI(\mem2[34][17] ), .SE(test_se), 
        .CLK(n2030), .Q(\mem2[34][18] ), .QN(n31470) );
  SDFFX1 \mem2_reg[34][17]  ( .D(n10685), .SI(\mem2[34][16] ), .SE(test_se), 
        .CLK(n2030), .Q(\mem2[34][17] ), .QN(n31471) );
  SDFFX1 \mem2_reg[34][16]  ( .D(n10684), .SI(\mem2[33][23] ), .SE(test_se), 
        .CLK(n2030), .Q(\mem2[34][16] ), .QN(n31472) );
  SDFFX1 \mem2_reg[33][23]  ( .D(n10683), .SI(\mem2[33][22] ), .SE(test_se), 
        .CLK(n2030), .Q(\mem2[33][23] ), .QN(n31473) );
  SDFFX1 \mem2_reg[33][22]  ( .D(n10682), .SI(\mem2[33][21] ), .SE(test_se), 
        .CLK(n2030), .Q(\mem2[33][22] ), .QN(n31474) );
  SDFFX1 \mem2_reg[33][21]  ( .D(n10681), .SI(\mem2[33][20] ), .SE(test_se), 
        .CLK(n2030), .Q(\mem2[33][21] ), .QN(n31475) );
  SDFFX1 \mem2_reg[33][20]  ( .D(n10680), .SI(\mem2[33][19] ), .SE(test_se), 
        .CLK(n2030), .Q(\mem2[33][20] ), .QN(n31476) );
  SDFFX1 \mem2_reg[33][19]  ( .D(n10679), .SI(\mem2[33][18] ), .SE(test_se), 
        .CLK(n2030), .Q(\mem2[33][19] ), .QN(n31477) );
  SDFFX1 \mem2_reg[33][18]  ( .D(n10678), .SI(\mem2[33][17] ), .SE(test_se), 
        .CLK(n2030), .Q(\mem2[33][18] ), .QN(n31478) );
  SDFFX1 \mem2_reg[33][17]  ( .D(n10677), .SI(\mem2[33][16] ), .SE(test_se), 
        .CLK(n2031), .Q(\mem2[33][17] ), .QN(n31479) );
  SDFFX1 \mem2_reg[33][16]  ( .D(n10676), .SI(\mem2[32][23] ), .SE(test_se), 
        .CLK(n2031), .Q(\mem2[33][16] ), .QN(n31480) );
  SDFFX1 \mem2_reg[32][23]  ( .D(n10675), .SI(\mem2[32][22] ), .SE(test_se), 
        .CLK(n2031), .Q(\mem2[32][23] ), .QN(n31481) );
  SDFFX1 \mem2_reg[32][22]  ( .D(n10674), .SI(\mem2[32][21] ), .SE(test_se), 
        .CLK(n2031), .Q(\mem2[32][22] ), .QN(n31482) );
  SDFFX1 \mem2_reg[32][21]  ( .D(n10673), .SI(\mem2[32][20] ), .SE(test_se), 
        .CLK(n2031), .Q(\mem2[32][21] ), .QN(n31483) );
  SDFFX1 \mem2_reg[32][20]  ( .D(n10672), .SI(\mem2[32][19] ), .SE(test_se), 
        .CLK(n2031), .Q(\mem2[32][20] ), .QN(n31484) );
  SDFFX1 \mem2_reg[32][19]  ( .D(n10671), .SI(\mem2[32][18] ), .SE(test_se), 
        .CLK(n2031), .Q(\mem2[32][19] ), .QN(n31485) );
  SDFFX1 \mem2_reg[32][18]  ( .D(n10670), .SI(\mem2[32][17] ), .SE(test_se), 
        .CLK(n2031), .Q(\mem2[32][18] ), .QN(n31486) );
  SDFFX1 \mem2_reg[32][17]  ( .D(n10669), .SI(\mem2[32][16] ), .SE(test_se), 
        .CLK(n2031), .Q(\mem2[32][17] ), .QN(n31487) );
  SDFFX1 \mem2_reg[32][16]  ( .D(n10668), .SI(\mem2[31][23] ), .SE(test_se), 
        .CLK(n2031), .Q(\mem2[32][16] ), .QN(n31488) );
  SDFFX1 \mem2_reg[31][23]  ( .D(n10667), .SI(\mem2[31][22] ), .SE(test_se), 
        .CLK(n2031), .Q(\mem2[31][23] ), .QN(n31489) );
  SDFFX1 \mem2_reg[31][22]  ( .D(n10666), .SI(\mem2[31][21] ), .SE(test_se), 
        .CLK(n2031), .Q(\mem2[31][22] ), .QN(n31490) );
  SDFFX1 \mem2_reg[31][21]  ( .D(n10665), .SI(\mem2[31][20] ), .SE(test_se), 
        .CLK(n2032), .Q(\mem2[31][21] ), .QN(n31491) );
  SDFFX1 \mem2_reg[31][20]  ( .D(n10664), .SI(\mem2[31][19] ), .SE(test_se), 
        .CLK(n2032), .Q(\mem2[31][20] ), .QN(n31492) );
  SDFFX1 \mem2_reg[31][19]  ( .D(n10663), .SI(\mem2[31][18] ), .SE(test_se), 
        .CLK(n2032), .Q(\mem2[31][19] ), .QN(n31493) );
  SDFFX1 \mem2_reg[31][18]  ( .D(n10662), .SI(\mem2[31][17] ), .SE(test_se), 
        .CLK(n2032), .Q(\mem2[31][18] ), .QN(n31494) );
  SDFFX1 \mem2_reg[31][17]  ( .D(n10661), .SI(\mem2[31][16] ), .SE(test_se), 
        .CLK(n2032), .Q(\mem2[31][17] ), .QN(n31495) );
  SDFFX1 \mem2_reg[31][16]  ( .D(n10660), .SI(\mem2[30][23] ), .SE(test_se), 
        .CLK(n2032), .Q(\mem2[31][16] ), .QN(n31496) );
  SDFFX1 \mem2_reg[30][23]  ( .D(n10659), .SI(\mem2[30][22] ), .SE(test_se), 
        .CLK(n2032), .Q(\mem2[30][23] ), .QN(n31497) );
  SDFFX1 \mem2_reg[30][22]  ( .D(n10658), .SI(\mem2[30][21] ), .SE(test_se), 
        .CLK(n2032), .Q(\mem2[30][22] ), .QN(n31498) );
  SDFFX1 \mem2_reg[30][21]  ( .D(n10657), .SI(\mem2[30][20] ), .SE(test_se), 
        .CLK(n2032), .Q(\mem2[30][21] ), .QN(n31499) );
  SDFFX1 \mem2_reg[30][20]  ( .D(n10656), .SI(\mem2[30][19] ), .SE(test_se), 
        .CLK(n2032), .Q(\mem2[30][20] ), .QN(n31500) );
  SDFFX1 \mem2_reg[30][19]  ( .D(n10655), .SI(\mem2[30][18] ), .SE(test_se), 
        .CLK(n2032), .Q(\mem2[30][19] ), .QN(n31501) );
  SDFFX1 \mem2_reg[30][18]  ( .D(n10654), .SI(\mem2[30][17] ), .SE(test_se), 
        .CLK(n2032), .Q(\mem2[30][18] ), .QN(n31502) );
  SDFFX1 \mem2_reg[30][17]  ( .D(n10653), .SI(\mem2[30][16] ), .SE(test_se), 
        .CLK(n2033), .Q(\mem2[30][17] ), .QN(n31503) );
  SDFFX1 \mem2_reg[30][16]  ( .D(n10652), .SI(\mem2[29][23] ), .SE(test_se), 
        .CLK(n2033), .Q(\mem2[30][16] ), .QN(n31504) );
  SDFFX1 \mem2_reg[29][23]  ( .D(n10651), .SI(\mem2[29][22] ), .SE(test_se), 
        .CLK(n2033), .Q(\mem2[29][23] ), .QN(n31505) );
  SDFFX1 \mem2_reg[29][22]  ( .D(n10650), .SI(\mem2[29][21] ), .SE(test_se), 
        .CLK(n2033), .Q(\mem2[29][22] ), .QN(n31506) );
  SDFFX1 \mem2_reg[29][21]  ( .D(n10649), .SI(\mem2[29][20] ), .SE(test_se), 
        .CLK(n2033), .Q(\mem2[29][21] ), .QN(n31507) );
  SDFFX1 \mem2_reg[29][20]  ( .D(n10648), .SI(\mem2[29][19] ), .SE(test_se), 
        .CLK(n2033), .Q(\mem2[29][20] ), .QN(n31508) );
  SDFFX1 \mem2_reg[29][19]  ( .D(n10647), .SI(\mem2[29][18] ), .SE(test_se), 
        .CLK(n2033), .Q(\mem2[29][19] ), .QN(n31509) );
  SDFFX1 \mem2_reg[29][18]  ( .D(n10646), .SI(\mem2[29][17] ), .SE(test_se), 
        .CLK(n2033), .Q(\mem2[29][18] ), .QN(n31510) );
  SDFFX1 \mem2_reg[29][17]  ( .D(n10645), .SI(\mem2[29][16] ), .SE(test_se), 
        .CLK(n2033), .Q(\mem2[29][17] ), .QN(n31511) );
  SDFFX1 \mem2_reg[29][16]  ( .D(n10644), .SI(\mem2[28][23] ), .SE(test_se), 
        .CLK(n2033), .Q(\mem2[29][16] ), .QN(n31512) );
  SDFFX1 \mem2_reg[28][23]  ( .D(n10643), .SI(\mem2[28][22] ), .SE(test_se), 
        .CLK(n2033), .Q(\mem2[28][23] ), .QN(n31513) );
  SDFFX1 \mem2_reg[28][22]  ( .D(n10642), .SI(\mem2[28][21] ), .SE(test_se), 
        .CLK(n2033), .Q(\mem2[28][22] ), .QN(n31514) );
  SDFFX1 \mem2_reg[28][21]  ( .D(n10641), .SI(\mem2[28][20] ), .SE(test_se), 
        .CLK(n2034), .Q(\mem2[28][21] ), .QN(n31515) );
  SDFFX1 \mem2_reg[28][20]  ( .D(n10640), .SI(\mem2[28][19] ), .SE(test_se), 
        .CLK(n2034), .Q(\mem2[28][20] ), .QN(n31516) );
  SDFFX1 \mem2_reg[28][19]  ( .D(n10639), .SI(\mem2[28][18] ), .SE(test_se), 
        .CLK(n2034), .Q(\mem2[28][19] ), .QN(n31517) );
  SDFFX1 \mem2_reg[28][18]  ( .D(n10638), .SI(\mem2[28][17] ), .SE(test_se), 
        .CLK(n2034), .Q(\mem2[28][18] ), .QN(n31518) );
  SDFFX1 \mem2_reg[28][17]  ( .D(n10637), .SI(\mem2[28][16] ), .SE(test_se), 
        .CLK(n2034), .Q(\mem2[28][17] ), .QN(n31519) );
  SDFFX1 \mem2_reg[28][16]  ( .D(n10636), .SI(\mem2[27][23] ), .SE(test_se), 
        .CLK(n2034), .Q(\mem2[28][16] ), .QN(n31520) );
  SDFFX1 \mem2_reg[27][23]  ( .D(n10635), .SI(\mem2[27][22] ), .SE(test_se), 
        .CLK(n2034), .Q(\mem2[27][23] ), .QN(n31521) );
  SDFFX1 \mem2_reg[27][22]  ( .D(n10634), .SI(\mem2[27][21] ), .SE(test_se), 
        .CLK(n2034), .Q(\mem2[27][22] ), .QN(n31522) );
  SDFFX1 \mem2_reg[27][21]  ( .D(n10633), .SI(\mem2[27][20] ), .SE(test_se), 
        .CLK(n2034), .Q(\mem2[27][21] ), .QN(n31523) );
  SDFFX1 \mem2_reg[27][20]  ( .D(n10632), .SI(\mem2[27][19] ), .SE(test_se), 
        .CLK(n2034), .Q(\mem2[27][20] ), .QN(n31524) );
  SDFFX1 \mem2_reg[27][19]  ( .D(n10631), .SI(\mem2[27][18] ), .SE(test_se), 
        .CLK(n2034), .Q(\mem2[27][19] ), .QN(n31525) );
  SDFFX1 \mem2_reg[27][18]  ( .D(n10630), .SI(\mem2[27][17] ), .SE(test_se), 
        .CLK(n2034), .Q(\mem2[27][18] ), .QN(n31526) );
  SDFFX1 \mem2_reg[27][17]  ( .D(n10629), .SI(\mem2[27][16] ), .SE(test_se), 
        .CLK(n2035), .Q(\mem2[27][17] ), .QN(n31527) );
  SDFFX1 \mem2_reg[27][16]  ( .D(n10628), .SI(\mem2[26][23] ), .SE(test_se), 
        .CLK(n2035), .Q(\mem2[27][16] ), .QN(n31528) );
  SDFFX1 \mem2_reg[26][23]  ( .D(n10627), .SI(\mem2[26][22] ), .SE(test_se), 
        .CLK(n2035), .Q(\mem2[26][23] ), .QN(n31529) );
  SDFFX1 \mem2_reg[26][22]  ( .D(n10626), .SI(\mem2[26][21] ), .SE(test_se), 
        .CLK(n2035), .Q(\mem2[26][22] ), .QN(n31530) );
  SDFFX1 \mem2_reg[26][21]  ( .D(n10625), .SI(\mem2[26][20] ), .SE(test_se), 
        .CLK(n2035), .Q(\mem2[26][21] ), .QN(n31531) );
  SDFFX1 \mem2_reg[26][20]  ( .D(n10624), .SI(\mem2[26][19] ), .SE(test_se), 
        .CLK(n2035), .Q(\mem2[26][20] ), .QN(n31532) );
  SDFFX1 \mem2_reg[26][19]  ( .D(n10623), .SI(\mem2[26][18] ), .SE(test_se), 
        .CLK(n2035), .Q(\mem2[26][19] ), .QN(n31533) );
  SDFFX1 \mem2_reg[26][18]  ( .D(n10622), .SI(\mem2[26][17] ), .SE(test_se), 
        .CLK(n2035), .Q(\mem2[26][18] ), .QN(n31534) );
  SDFFX1 \mem2_reg[26][17]  ( .D(n10621), .SI(\mem2[26][16] ), .SE(test_se), 
        .CLK(n2035), .Q(\mem2[26][17] ), .QN(n31535) );
  SDFFX1 \mem2_reg[26][16]  ( .D(n10620), .SI(\mem2[25][23] ), .SE(test_se), 
        .CLK(n2035), .Q(\mem2[26][16] ), .QN(n31536) );
  SDFFX1 \mem2_reg[25][23]  ( .D(n10619), .SI(\mem2[25][22] ), .SE(test_se), 
        .CLK(n2035), .Q(\mem2[25][23] ), .QN(n31537) );
  SDFFX1 \mem2_reg[25][22]  ( .D(n10618), .SI(\mem2[25][21] ), .SE(test_se), 
        .CLK(n2035), .Q(\mem2[25][22] ), .QN(n31538) );
  SDFFX1 \mem2_reg[25][21]  ( .D(n10617), .SI(\mem2[25][20] ), .SE(test_se), 
        .CLK(n2036), .Q(\mem2[25][21] ), .QN(n31539) );
  SDFFX1 \mem2_reg[25][20]  ( .D(n10616), .SI(\mem2[25][19] ), .SE(test_se), 
        .CLK(n2036), .Q(\mem2[25][20] ), .QN(n31540) );
  SDFFX1 \mem2_reg[25][19]  ( .D(n10615), .SI(\mem2[25][18] ), .SE(test_se), 
        .CLK(n2036), .Q(\mem2[25][19] ), .QN(n31541) );
  SDFFX1 \mem2_reg[25][18]  ( .D(n10614), .SI(\mem2[25][17] ), .SE(test_se), 
        .CLK(n2036), .Q(\mem2[25][18] ), .QN(n31542) );
  SDFFX1 \mem2_reg[25][17]  ( .D(n10613), .SI(\mem2[25][16] ), .SE(test_se), 
        .CLK(n2036), .Q(\mem2[25][17] ), .QN(n31543) );
  SDFFX1 \mem2_reg[25][16]  ( .D(n10612), .SI(\mem2[24][23] ), .SE(test_se), 
        .CLK(n2036), .Q(\mem2[25][16] ), .QN(n31544) );
  SDFFX1 \mem2_reg[24][23]  ( .D(n10611), .SI(\mem2[24][22] ), .SE(test_se), 
        .CLK(n2036), .Q(\mem2[24][23] ), .QN(n31545) );
  SDFFX1 \mem2_reg[24][22]  ( .D(n10610), .SI(\mem2[24][21] ), .SE(test_se), 
        .CLK(n2036), .Q(\mem2[24][22] ), .QN(n31546) );
  SDFFX1 \mem2_reg[24][21]  ( .D(n10609), .SI(\mem2[24][20] ), .SE(test_se), 
        .CLK(n2036), .Q(\mem2[24][21] ), .QN(n31547) );
  SDFFX1 \mem2_reg[24][20]  ( .D(n10608), .SI(\mem2[24][19] ), .SE(test_se), 
        .CLK(n2036), .Q(\mem2[24][20] ), .QN(n31548) );
  SDFFX1 \mem2_reg[24][19]  ( .D(n10607), .SI(\mem2[24][18] ), .SE(test_se), 
        .CLK(n2036), .Q(\mem2[24][19] ), .QN(n31549) );
  SDFFX1 \mem2_reg[24][18]  ( .D(n10606), .SI(\mem2[24][17] ), .SE(test_se), 
        .CLK(n2036), .Q(\mem2[24][18] ), .QN(n31550) );
  SDFFX1 \mem2_reg[24][17]  ( .D(n10605), .SI(\mem2[24][16] ), .SE(test_se), 
        .CLK(n2037), .Q(\mem2[24][17] ), .QN(n31551) );
  SDFFX1 \mem2_reg[24][16]  ( .D(n10604), .SI(\mem2[23][23] ), .SE(test_se), 
        .CLK(n2037), .Q(\mem2[24][16] ), .QN(n31552) );
  SDFFX1 \mem2_reg[23][23]  ( .D(n10603), .SI(\mem2[23][22] ), .SE(test_se), 
        .CLK(n2037), .Q(\mem2[23][23] ), .QN(n31553) );
  SDFFX1 \mem2_reg[23][22]  ( .D(n10602), .SI(\mem2[23][21] ), .SE(test_se), 
        .CLK(n2037), .Q(\mem2[23][22] ), .QN(n31554) );
  SDFFX1 \mem2_reg[23][21]  ( .D(n10601), .SI(\mem2[23][20] ), .SE(test_se), 
        .CLK(n2037), .Q(\mem2[23][21] ), .QN(n31555) );
  SDFFX1 \mem2_reg[23][20]  ( .D(n10600), .SI(\mem2[23][19] ), .SE(test_se), 
        .CLK(n2037), .Q(\mem2[23][20] ), .QN(n31556) );
  SDFFX1 \mem2_reg[23][19]  ( .D(n10599), .SI(\mem2[23][18] ), .SE(test_se), 
        .CLK(n2037), .Q(\mem2[23][19] ), .QN(n31557) );
  SDFFX1 \mem2_reg[23][18]  ( .D(n10598), .SI(\mem2[23][17] ), .SE(test_se), 
        .CLK(n2037), .Q(\mem2[23][18] ), .QN(n31558) );
  SDFFX1 \mem2_reg[23][17]  ( .D(n10597), .SI(\mem2[23][16] ), .SE(test_se), 
        .CLK(n2037), .Q(\mem2[23][17] ), .QN(n31559) );
  SDFFX1 \mem2_reg[23][16]  ( .D(n10596), .SI(\mem2[22][23] ), .SE(test_se), 
        .CLK(n2037), .Q(\mem2[23][16] ), .QN(n31560) );
  SDFFX1 \mem2_reg[22][23]  ( .D(n10595), .SI(\mem2[22][22] ), .SE(test_se), 
        .CLK(n2037), .Q(\mem2[22][23] ), .QN(n31561) );
  SDFFX1 \mem2_reg[22][22]  ( .D(n10594), .SI(\mem2[22][21] ), .SE(test_se), 
        .CLK(n2037), .Q(\mem2[22][22] ), .QN(n31562) );
  SDFFX1 \mem2_reg[22][21]  ( .D(n10593), .SI(\mem2[22][20] ), .SE(test_se), 
        .CLK(n2038), .Q(\mem2[22][21] ), .QN(n31563) );
  SDFFX1 \mem2_reg[22][20]  ( .D(n10592), .SI(\mem2[22][19] ), .SE(test_se), 
        .CLK(n2038), .Q(\mem2[22][20] ), .QN(n31564) );
  SDFFX1 \mem2_reg[22][19]  ( .D(n10591), .SI(\mem2[22][18] ), .SE(test_se), 
        .CLK(n2038), .Q(\mem2[22][19] ), .QN(n31565) );
  SDFFX1 \mem2_reg[22][18]  ( .D(n10590), .SI(\mem2[22][17] ), .SE(test_se), 
        .CLK(n2038), .Q(\mem2[22][18] ), .QN(n31566) );
  SDFFX1 \mem2_reg[22][17]  ( .D(n10589), .SI(\mem2[22][16] ), .SE(test_se), 
        .CLK(n2038), .Q(\mem2[22][17] ), .QN(n31567) );
  SDFFX1 \mem2_reg[22][16]  ( .D(n10588), .SI(\mem2[21][23] ), .SE(test_se), 
        .CLK(n2038), .Q(\mem2[22][16] ), .QN(n31568) );
  SDFFX1 \mem2_reg[21][23]  ( .D(n10587), .SI(\mem2[21][22] ), .SE(test_se), 
        .CLK(n2038), .Q(\mem2[21][23] ), .QN(n31569) );
  SDFFX1 \mem2_reg[21][22]  ( .D(n10586), .SI(\mem2[21][21] ), .SE(test_se), 
        .CLK(n2038), .Q(\mem2[21][22] ), .QN(n31570) );
  SDFFX1 \mem2_reg[21][21]  ( .D(n10585), .SI(\mem2[21][20] ), .SE(test_se), 
        .CLK(n2038), .Q(\mem2[21][21] ), .QN(n31571) );
  SDFFX1 \mem2_reg[21][20]  ( .D(n10584), .SI(\mem2[21][19] ), .SE(test_se), 
        .CLK(n2038), .Q(\mem2[21][20] ), .QN(n31572) );
  SDFFX1 \mem2_reg[21][19]  ( .D(n10583), .SI(\mem2[21][18] ), .SE(test_se), 
        .CLK(n2038), .Q(\mem2[21][19] ), .QN(n31573) );
  SDFFX1 \mem2_reg[21][18]  ( .D(n10582), .SI(\mem2[21][17] ), .SE(test_se), 
        .CLK(n2038), .Q(\mem2[21][18] ), .QN(n31574) );
  SDFFX1 \mem2_reg[21][17]  ( .D(n10581), .SI(\mem2[21][16] ), .SE(test_se), 
        .CLK(n2039), .Q(\mem2[21][17] ), .QN(n31575) );
  SDFFX1 \mem2_reg[21][16]  ( .D(n10580), .SI(\mem2[20][23] ), .SE(test_se), 
        .CLK(n2039), .Q(\mem2[21][16] ), .QN(n31576) );
  SDFFX1 \mem2_reg[20][23]  ( .D(n10579), .SI(\mem2[20][22] ), .SE(test_se), 
        .CLK(n2039), .Q(\mem2[20][23] ), .QN(n31577) );
  SDFFX1 \mem2_reg[20][22]  ( .D(n10578), .SI(\mem2[20][21] ), .SE(test_se), 
        .CLK(n2039), .Q(\mem2[20][22] ), .QN(n31578) );
  SDFFX1 \mem2_reg[20][21]  ( .D(n10577), .SI(\mem2[20][20] ), .SE(test_se), 
        .CLK(n2039), .Q(\mem2[20][21] ), .QN(n31579) );
  SDFFX1 \mem2_reg[20][20]  ( .D(n10576), .SI(\mem2[20][19] ), .SE(test_se), 
        .CLK(n2039), .Q(\mem2[20][20] ), .QN(n31580) );
  SDFFX1 \mem2_reg[20][19]  ( .D(n10575), .SI(\mem2[20][18] ), .SE(test_se), 
        .CLK(n2039), .Q(\mem2[20][19] ), .QN(n31581) );
  SDFFX1 \mem2_reg[20][18]  ( .D(n10574), .SI(\mem2[20][17] ), .SE(test_se), 
        .CLK(n2039), .Q(\mem2[20][18] ), .QN(n31582) );
  SDFFX1 \mem2_reg[20][17]  ( .D(n10573), .SI(\mem2[20][16] ), .SE(test_se), 
        .CLK(n2039), .Q(\mem2[20][17] ), .QN(n31583) );
  SDFFX1 \mem2_reg[20][16]  ( .D(n10572), .SI(\mem2[19][23] ), .SE(test_se), 
        .CLK(n2039), .Q(\mem2[20][16] ), .QN(n31584) );
  SDFFX1 \mem2_reg[19][23]  ( .D(n10571), .SI(\mem2[19][22] ), .SE(test_se), 
        .CLK(n2039), .Q(\mem2[19][23] ), .QN(n31585) );
  SDFFX1 \mem2_reg[19][22]  ( .D(n10570), .SI(\mem2[19][21] ), .SE(test_se), 
        .CLK(n2039), .Q(\mem2[19][22] ), .QN(n31586) );
  SDFFX1 \mem2_reg[19][21]  ( .D(n10569), .SI(\mem2[19][20] ), .SE(test_se), 
        .CLK(n2040), .Q(\mem2[19][21] ), .QN(n31587) );
  SDFFX1 \mem2_reg[19][20]  ( .D(n10568), .SI(\mem2[19][19] ), .SE(test_se), 
        .CLK(n2040), .Q(\mem2[19][20] ), .QN(n31588) );
  SDFFX1 \mem2_reg[19][19]  ( .D(n10567), .SI(\mem2[19][18] ), .SE(test_se), 
        .CLK(n2040), .Q(\mem2[19][19] ), .QN(n31589) );
  SDFFX1 \mem2_reg[19][18]  ( .D(n10566), .SI(\mem2[19][17] ), .SE(test_se), 
        .CLK(n2040), .Q(\mem2[19][18] ), .QN(n31590) );
  SDFFX1 \mem2_reg[19][17]  ( .D(n10565), .SI(\mem2[19][16] ), .SE(test_se), 
        .CLK(n2040), .Q(\mem2[19][17] ), .QN(n31591) );
  SDFFX1 \mem2_reg[19][16]  ( .D(n10564), .SI(\mem2[18][23] ), .SE(test_se), 
        .CLK(n2040), .Q(\mem2[19][16] ), .QN(n31592) );
  SDFFX1 \mem2_reg[18][23]  ( .D(n10563), .SI(\mem2[18][22] ), .SE(test_se), 
        .CLK(n2040), .Q(\mem2[18][23] ), .QN(n31593) );
  SDFFX1 \mem2_reg[18][22]  ( .D(n10562), .SI(\mem2[18][21] ), .SE(test_se), 
        .CLK(n2040), .Q(\mem2[18][22] ), .QN(n31594) );
  SDFFX1 \mem2_reg[18][21]  ( .D(n10561), .SI(\mem2[18][20] ), .SE(test_se), 
        .CLK(n2040), .Q(\mem2[18][21] ), .QN(n31595) );
  SDFFX1 \mem2_reg[18][20]  ( .D(n10560), .SI(\mem2[18][19] ), .SE(test_se), 
        .CLK(n2040), .Q(\mem2[18][20] ), .QN(n31596) );
  SDFFX1 \mem2_reg[18][19]  ( .D(n10559), .SI(\mem2[18][18] ), .SE(test_se), 
        .CLK(n2040), .Q(\mem2[18][19] ), .QN(n31597) );
  SDFFX1 \mem2_reg[18][18]  ( .D(n10558), .SI(\mem2[18][17] ), .SE(test_se), 
        .CLK(n2040), .Q(\mem2[18][18] ), .QN(n31598) );
  SDFFX1 \mem2_reg[18][17]  ( .D(n10557), .SI(\mem2[18][16] ), .SE(test_se), 
        .CLK(n2041), .Q(\mem2[18][17] ), .QN(n31599) );
  SDFFX1 \mem2_reg[18][16]  ( .D(n10556), .SI(\mem2[17][23] ), .SE(test_se), 
        .CLK(n2041), .Q(\mem2[18][16] ), .QN(n31600) );
  SDFFX1 \mem2_reg[17][23]  ( .D(n10555), .SI(\mem2[17][22] ), .SE(test_se), 
        .CLK(n2041), .Q(\mem2[17][23] ), .QN(n31601) );
  SDFFX1 \mem2_reg[17][22]  ( .D(n10554), .SI(\mem2[17][21] ), .SE(test_se), 
        .CLK(n2041), .Q(\mem2[17][22] ), .QN(n31602) );
  SDFFX1 \mem2_reg[17][21]  ( .D(n10553), .SI(\mem2[17][20] ), .SE(test_se), 
        .CLK(n2041), .Q(\mem2[17][21] ), .QN(n31603) );
  SDFFX1 \mem2_reg[17][20]  ( .D(n10552), .SI(\mem2[17][19] ), .SE(test_se), 
        .CLK(n2041), .Q(\mem2[17][20] ), .QN(n31604) );
  SDFFX1 \mem2_reg[17][19]  ( .D(n10551), .SI(\mem2[17][18] ), .SE(test_se), 
        .CLK(n2041), .Q(\mem2[17][19] ), .QN(n31605) );
  SDFFX1 \mem2_reg[17][18]  ( .D(n10550), .SI(\mem2[17][17] ), .SE(test_se), 
        .CLK(n2041), .Q(\mem2[17][18] ), .QN(n31606) );
  SDFFX1 \mem2_reg[17][17]  ( .D(n10549), .SI(\mem2[17][16] ), .SE(test_se), 
        .CLK(n2041), .Q(\mem2[17][17] ), .QN(n31607) );
  SDFFX1 \mem2_reg[17][16]  ( .D(n10548), .SI(\mem2[16][23] ), .SE(test_se), 
        .CLK(n2041), .Q(\mem2[17][16] ), .QN(n31608) );
  SDFFX1 \mem2_reg[16][23]  ( .D(n10547), .SI(\mem2[16][22] ), .SE(test_se), 
        .CLK(n2041), .Q(\mem2[16][23] ), .QN(n31609) );
  SDFFX1 \mem2_reg[16][22]  ( .D(n10546), .SI(\mem2[16][21] ), .SE(test_se), 
        .CLK(n2041), .Q(\mem2[16][22] ), .QN(n31610) );
  SDFFX1 \mem2_reg[16][21]  ( .D(n10545), .SI(\mem2[16][20] ), .SE(test_se), 
        .CLK(n2042), .Q(\mem2[16][21] ), .QN(n31611) );
  SDFFX1 \mem2_reg[16][20]  ( .D(n10544), .SI(\mem2[16][19] ), .SE(test_se), 
        .CLK(n2042), .Q(\mem2[16][20] ), .QN(n31612) );
  SDFFX1 \mem2_reg[16][19]  ( .D(n10543), .SI(\mem2[16][18] ), .SE(test_se), 
        .CLK(n2042), .Q(\mem2[16][19] ), .QN(n31613) );
  SDFFX1 \mem2_reg[16][18]  ( .D(n10542), .SI(\mem2[16][17] ), .SE(test_se), 
        .CLK(n2042), .Q(\mem2[16][18] ), .QN(n31614) );
  SDFFX1 \mem2_reg[16][17]  ( .D(n10541), .SI(\mem2[16][16] ), .SE(test_se), 
        .CLK(n2042), .Q(\mem2[16][17] ), .QN(n31615) );
  SDFFX1 \mem2_reg[16][16]  ( .D(n10540), .SI(\mem2[15][23] ), .SE(test_se), 
        .CLK(n2042), .Q(\mem2[16][16] ), .QN(n31616) );
  SDFFX1 \mem2_reg[15][23]  ( .D(n10539), .SI(\mem2[15][22] ), .SE(test_se), 
        .CLK(n2042), .Q(\mem2[15][23] ), .QN(n31617) );
  SDFFX1 \mem2_reg[15][22]  ( .D(n10538), .SI(\mem2[15][21] ), .SE(test_se), 
        .CLK(n2042), .Q(\mem2[15][22] ), .QN(n31618) );
  SDFFX1 \mem2_reg[15][21]  ( .D(n10537), .SI(\mem2[15][20] ), .SE(test_se), 
        .CLK(n2042), .Q(\mem2[15][21] ), .QN(n31619) );
  SDFFX1 \mem2_reg[15][20]  ( .D(n10536), .SI(\mem2[15][19] ), .SE(test_se), 
        .CLK(n2042), .Q(\mem2[15][20] ), .QN(n31620) );
  SDFFX1 \mem2_reg[15][19]  ( .D(n10535), .SI(\mem2[15][18] ), .SE(test_se), 
        .CLK(n2042), .Q(\mem2[15][19] ), .QN(n31621) );
  SDFFX1 \mem2_reg[15][18]  ( .D(n10534), .SI(\mem2[15][17] ), .SE(test_se), 
        .CLK(n2042), .Q(\mem2[15][18] ), .QN(n31622) );
  SDFFX1 \mem2_reg[15][17]  ( .D(n10533), .SI(\mem2[15][16] ), .SE(test_se), 
        .CLK(n2043), .Q(\mem2[15][17] ), .QN(n31623) );
  SDFFX1 \mem2_reg[15][16]  ( .D(n10532), .SI(\mem2[14][23] ), .SE(test_se), 
        .CLK(n2043), .Q(\mem2[15][16] ), .QN(n31624) );
  SDFFX1 \mem2_reg[14][23]  ( .D(n10531), .SI(\mem2[14][22] ), .SE(test_se), 
        .CLK(n2043), .Q(\mem2[14][23] ), .QN(n31625) );
  SDFFX1 \mem2_reg[14][22]  ( .D(n10530), .SI(\mem2[14][21] ), .SE(test_se), 
        .CLK(n2043), .Q(\mem2[14][22] ), .QN(n31626) );
  SDFFX1 \mem2_reg[14][21]  ( .D(n10529), .SI(\mem2[14][20] ), .SE(test_se), 
        .CLK(n2043), .Q(\mem2[14][21] ), .QN(n31627) );
  SDFFX1 \mem2_reg[14][20]  ( .D(n10528), .SI(\mem2[14][19] ), .SE(test_se), 
        .CLK(n2043), .Q(\mem2[14][20] ), .QN(n31628) );
  SDFFX1 \mem2_reg[14][19]  ( .D(n10527), .SI(\mem2[14][18] ), .SE(test_se), 
        .CLK(n2043), .Q(\mem2[14][19] ), .QN(n31629) );
  SDFFX1 \mem2_reg[14][18]  ( .D(n10526), .SI(\mem2[14][17] ), .SE(test_se), 
        .CLK(n2043), .Q(\mem2[14][18] ), .QN(n31630) );
  SDFFX1 \mem2_reg[14][17]  ( .D(n10525), .SI(\mem2[14][16] ), .SE(test_se), 
        .CLK(n2043), .Q(\mem2[14][17] ), .QN(n31631) );
  SDFFX1 \mem2_reg[14][16]  ( .D(n10524), .SI(\mem2[13][23] ), .SE(test_se), 
        .CLK(n2043), .Q(\mem2[14][16] ), .QN(n31632) );
  SDFFX1 \mem2_reg[13][23]  ( .D(n10523), .SI(\mem2[13][22] ), .SE(test_se), 
        .CLK(n2043), .Q(\mem2[13][23] ), .QN(n31633) );
  SDFFX1 \mem2_reg[13][22]  ( .D(n10522), .SI(\mem2[13][21] ), .SE(test_se), 
        .CLK(n2043), .Q(\mem2[13][22] ), .QN(n31634) );
  SDFFX1 \mem2_reg[13][21]  ( .D(n10521), .SI(\mem2[13][20] ), .SE(test_se), 
        .CLK(n2044), .Q(\mem2[13][21] ), .QN(n31635) );
  SDFFX1 \mem2_reg[13][20]  ( .D(n10520), .SI(\mem2[13][19] ), .SE(test_se), 
        .CLK(n2044), .Q(\mem2[13][20] ), .QN(n31636) );
  SDFFX1 \mem2_reg[13][19]  ( .D(n10519), .SI(\mem2[13][18] ), .SE(test_se), 
        .CLK(n2044), .Q(\mem2[13][19] ), .QN(n31637) );
  SDFFX1 \mem2_reg[13][18]  ( .D(n10518), .SI(\mem2[13][17] ), .SE(test_se), 
        .CLK(n2044), .Q(\mem2[13][18] ), .QN(n31638) );
  SDFFX1 \mem2_reg[13][17]  ( .D(n10517), .SI(\mem2[13][16] ), .SE(test_se), 
        .CLK(n2044), .Q(\mem2[13][17] ), .QN(n31639) );
  SDFFX1 \mem2_reg[13][16]  ( .D(n10516), .SI(\mem2[12][23] ), .SE(test_se), 
        .CLK(n2044), .Q(\mem2[13][16] ), .QN(n31640) );
  SDFFX1 \mem2_reg[12][23]  ( .D(n10515), .SI(\mem2[12][22] ), .SE(test_se), 
        .CLK(n2044), .Q(\mem2[12][23] ), .QN(n31641) );
  SDFFX1 \mem2_reg[12][22]  ( .D(n10514), .SI(\mem2[12][21] ), .SE(test_se), 
        .CLK(n2044), .Q(\mem2[12][22] ), .QN(n31642) );
  SDFFX1 \mem2_reg[12][21]  ( .D(n10513), .SI(\mem2[12][20] ), .SE(test_se), 
        .CLK(n2044), .Q(\mem2[12][21] ), .QN(n31643) );
  SDFFX1 \mem2_reg[12][20]  ( .D(n10512), .SI(\mem2[12][19] ), .SE(test_se), 
        .CLK(n2044), .Q(\mem2[12][20] ), .QN(n31644) );
  SDFFX1 \mem2_reg[12][19]  ( .D(n10511), .SI(\mem2[12][18] ), .SE(test_se), 
        .CLK(n2044), .Q(\mem2[12][19] ), .QN(n31645) );
  SDFFX1 \mem2_reg[12][18]  ( .D(n10510), .SI(\mem2[12][17] ), .SE(test_se), 
        .CLK(n2044), .Q(\mem2[12][18] ), .QN(n31646) );
  SDFFX1 \mem2_reg[12][17]  ( .D(n10509), .SI(\mem2[12][16] ), .SE(test_se), 
        .CLK(n2045), .Q(\mem2[12][17] ), .QN(n31647) );
  SDFFX1 \mem2_reg[12][16]  ( .D(n10508), .SI(\mem2[11][23] ), .SE(test_se), 
        .CLK(n2045), .Q(\mem2[12][16] ), .QN(n31648) );
  SDFFX1 \mem2_reg[11][23]  ( .D(n10507), .SI(\mem2[11][22] ), .SE(test_se), 
        .CLK(n2053), .Q(\mem2[11][23] ), .QN(n31649) );
  SDFFX1 \mem2_reg[11][22]  ( .D(n10506), .SI(\mem2[11][21] ), .SE(test_se), 
        .CLK(n2053), .Q(\mem2[11][22] ), .QN(n31650) );
  SDFFX1 \mem2_reg[11][21]  ( .D(n10505), .SI(\mem2[11][20] ), .SE(test_se), 
        .CLK(n2053), .Q(\mem2[11][21] ), .QN(n31651) );
  SDFFX1 \mem2_reg[11][20]  ( .D(n10504), .SI(\mem2[11][19] ), .SE(test_se), 
        .CLK(n2053), .Q(\mem2[11][20] ), .QN(n31652) );
  SDFFX1 \mem2_reg[11][19]  ( .D(n10503), .SI(\mem2[11][18] ), .SE(test_se), 
        .CLK(n2053), .Q(\mem2[11][19] ), .QN(n31653) );
  SDFFX1 \mem2_reg[11][18]  ( .D(n10502), .SI(\mem2[11][17] ), .SE(test_se), 
        .CLK(n2053), .Q(\mem2[11][18] ), .QN(n31654) );
  SDFFX1 \mem2_reg[11][17]  ( .D(n10501), .SI(\mem2[11][16] ), .SE(test_se), 
        .CLK(n2053), .Q(\mem2[11][17] ), .QN(n31655) );
  SDFFX1 \mem2_reg[11][16]  ( .D(n10500), .SI(\mem2[10][23] ), .SE(test_se), 
        .CLK(n2053), .Q(\mem2[11][16] ), .QN(n31656) );
  SDFFX1 \mem2_reg[10][23]  ( .D(n10499), .SI(\mem2[10][22] ), .SE(test_se), 
        .CLK(n2053), .Q(\mem2[10][23] ), .QN(n31657) );
  SDFFX1 \mem2_reg[10][22]  ( .D(n10498), .SI(\mem2[10][21] ), .SE(test_se), 
        .CLK(n2053), .Q(\mem2[10][22] ), .QN(n31658) );
  SDFFX1 \mem2_reg[10][21]  ( .D(n10497), .SI(\mem2[10][20] ), .SE(test_se), 
        .CLK(n2054), .Q(\mem2[10][21] ), .QN(n31659) );
  SDFFX1 \mem2_reg[10][20]  ( .D(n10496), .SI(\mem2[10][19] ), .SE(test_se), 
        .CLK(n2054), .Q(\mem2[10][20] ), .QN(n31660) );
  SDFFX1 \mem2_reg[10][19]  ( .D(n10495), .SI(\mem2[10][18] ), .SE(test_se), 
        .CLK(n2054), .Q(\mem2[10][19] ), .QN(n31661) );
  SDFFX1 \mem2_reg[10][18]  ( .D(n10494), .SI(\mem2[10][17] ), .SE(test_se), 
        .CLK(n2054), .Q(\mem2[10][18] ), .QN(n31662) );
  SDFFX1 \mem2_reg[10][17]  ( .D(n10493), .SI(\mem2[10][16] ), .SE(test_se), 
        .CLK(n2054), .Q(\mem2[10][17] ), .QN(n31663) );
  SDFFX1 \mem2_reg[10][16]  ( .D(n10492), .SI(\mem2[9][23] ), .SE(test_se), 
        .CLK(n2054), .Q(\mem2[10][16] ), .QN(n31664) );
  SDFFX1 \mem2_reg[9][23]  ( .D(n10491), .SI(\mem2[9][22] ), .SE(test_se), 
        .CLK(n2054), .Q(\mem2[9][23] ), .QN(n31665) );
  SDFFX1 \mem2_reg[9][22]  ( .D(n10490), .SI(\mem2[9][21] ), .SE(test_se), 
        .CLK(n2054), .Q(\mem2[9][22] ), .QN(n31666) );
  SDFFX1 \mem2_reg[9][21]  ( .D(n10489), .SI(\mem2[9][20] ), .SE(test_se), 
        .CLK(n2054), .Q(\mem2[9][21] ), .QN(n31667) );
  SDFFX1 \mem2_reg[9][20]  ( .D(n10488), .SI(\mem2[9][19] ), .SE(test_se), 
        .CLK(n2054), .Q(\mem2[9][20] ), .QN(n31668) );
  SDFFX1 \mem2_reg[9][19]  ( .D(n10487), .SI(\mem2[9][18] ), .SE(test_se), 
        .CLK(n2054), .Q(\mem2[9][19] ), .QN(n31669) );
  SDFFX1 \mem2_reg[9][18]  ( .D(n10486), .SI(\mem2[9][17] ), .SE(test_se), 
        .CLK(n2054), .Q(\mem2[9][18] ), .QN(n31670) );
  SDFFX1 \mem2_reg[9][17]  ( .D(n10485), .SI(\mem2[9][16] ), .SE(test_se), 
        .CLK(n2055), .Q(\mem2[9][17] ), .QN(n31671) );
  SDFFX1 \mem2_reg[9][16]  ( .D(n10484), .SI(\mem2[8][23] ), .SE(test_se), 
        .CLK(n2055), .Q(\mem2[9][16] ), .QN(n31672) );
  SDFFX1 \mem2_reg[8][23]  ( .D(n10483), .SI(\mem2[8][22] ), .SE(test_se), 
        .CLK(n2055), .Q(\mem2[8][23] ), .QN(n31673) );
  SDFFX1 \mem2_reg[8][22]  ( .D(n10482), .SI(\mem2[8][21] ), .SE(test_se), 
        .CLK(n2055), .Q(\mem2[8][22] ), .QN(n31674) );
  SDFFX1 \mem2_reg[8][21]  ( .D(n10481), .SI(\mem2[8][20] ), .SE(test_se), 
        .CLK(n2055), .Q(\mem2[8][21] ), .QN(n31675) );
  SDFFX1 \mem2_reg[8][20]  ( .D(n10480), .SI(\mem2[8][19] ), .SE(test_se), 
        .CLK(n2055), .Q(\mem2[8][20] ), .QN(n31676) );
  SDFFX1 \mem2_reg[8][19]  ( .D(n10479), .SI(\mem2[8][18] ), .SE(test_se), 
        .CLK(n2055), .Q(\mem2[8][19] ), .QN(n31677) );
  SDFFX1 \mem2_reg[8][18]  ( .D(n10478), .SI(\mem2[8][17] ), .SE(test_se), 
        .CLK(n2055), .Q(\mem2[8][18] ), .QN(n31678) );
  SDFFX1 \mem2_reg[8][17]  ( .D(n10477), .SI(\mem2[8][16] ), .SE(test_se), 
        .CLK(n2055), .Q(\mem2[8][17] ), .QN(n31679) );
  SDFFX1 \mem2_reg[8][16]  ( .D(n10476), .SI(\mem2[7][23] ), .SE(test_se), 
        .CLK(n2055), .Q(\mem2[8][16] ), .QN(n31680) );
  SDFFX1 \mem2_reg[7][23]  ( .D(n10475), .SI(\mem2[7][22] ), .SE(test_se), 
        .CLK(n2063), .Q(\mem2[7][23] ), .QN(n31681) );
  SDFFX1 \mem2_reg[7][22]  ( .D(n10474), .SI(\mem2[7][21] ), .SE(test_se), 
        .CLK(n2063), .Q(\mem2[7][22] ), .QN(n31682) );
  SDFFX1 \mem2_reg[7][21]  ( .D(n10473), .SI(\mem2[7][20] ), .SE(test_se), 
        .CLK(n2064), .Q(\mem2[7][21] ), .QN(n31683) );
  SDFFX1 \mem2_reg[7][20]  ( .D(n10472), .SI(\mem2[7][19] ), .SE(test_se), 
        .CLK(n2064), .Q(\mem2[7][20] ), .QN(n31684) );
  SDFFX1 \mem2_reg[7][19]  ( .D(n10471), .SI(\mem2[7][18] ), .SE(test_se), 
        .CLK(n2064), .Q(\mem2[7][19] ), .QN(n31685) );
  SDFFX1 \mem2_reg[7][18]  ( .D(n10470), .SI(\mem2[7][17] ), .SE(test_se), 
        .CLK(n2064), .Q(\mem2[7][18] ), .QN(n31686) );
  SDFFX1 \mem2_reg[7][17]  ( .D(n10469), .SI(\mem2[7][16] ), .SE(test_se), 
        .CLK(n2064), .Q(\mem2[7][17] ), .QN(n31687) );
  SDFFX1 \mem2_reg[7][16]  ( .D(n10468), .SI(\mem2[6][23] ), .SE(test_se), 
        .CLK(n2064), .Q(\mem2[7][16] ), .QN(n31688) );
  SDFFX1 \mem2_reg[6][23]  ( .D(n10467), .SI(\mem2[6][22] ), .SE(test_se), 
        .CLK(n2064), .Q(\mem2[6][23] ), .QN(n31689) );
  SDFFX1 \mem2_reg[6][22]  ( .D(n10466), .SI(\mem2[6][21] ), .SE(test_se), 
        .CLK(n2064), .Q(\mem2[6][22] ), .QN(n31690) );
  SDFFX1 \mem2_reg[6][21]  ( .D(n10465), .SI(\mem2[6][20] ), .SE(test_se), 
        .CLK(n2064), .Q(\mem2[6][21] ), .QN(n31691) );
  SDFFX1 \mem2_reg[6][20]  ( .D(n10464), .SI(\mem2[6][19] ), .SE(test_se), 
        .CLK(n2064), .Q(\mem2[6][20] ), .QN(n31692) );
  SDFFX1 \mem2_reg[6][19]  ( .D(n10463), .SI(\mem2[6][18] ), .SE(test_se), 
        .CLK(n2064), .Q(\mem2[6][19] ), .QN(n31693) );
  SDFFX1 \mem2_reg[6][18]  ( .D(n10462), .SI(\mem2[6][17] ), .SE(test_se), 
        .CLK(n2064), .Q(\mem2[6][18] ), .QN(n31694) );
  SDFFX1 \mem2_reg[6][17]  ( .D(n10461), .SI(\mem2[6][16] ), .SE(test_se), 
        .CLK(n2065), .Q(\mem2[6][17] ), .QN(n31695) );
  SDFFX1 \mem2_reg[6][16]  ( .D(n10460), .SI(\mem2[5][23] ), .SE(test_se), 
        .CLK(n2065), .Q(\mem2[6][16] ), .QN(n31696) );
  SDFFX1 \mem2_reg[5][23]  ( .D(n10459), .SI(\mem2[5][22] ), .SE(test_se), 
        .CLK(n2065), .Q(\mem2[5][23] ), .QN(n31697) );
  SDFFX1 \mem2_reg[5][22]  ( .D(n10458), .SI(\mem2[5][21] ), .SE(test_se), 
        .CLK(n2065), .Q(\mem2[5][22] ), .QN(n31698) );
  SDFFX1 \mem2_reg[5][21]  ( .D(n10457), .SI(\mem2[5][20] ), .SE(test_se), 
        .CLK(n2065), .Q(\mem2[5][21] ), .QN(n31699) );
  SDFFX1 \mem2_reg[5][20]  ( .D(n10456), .SI(\mem2[5][19] ), .SE(test_se), 
        .CLK(n2065), .Q(\mem2[5][20] ), .QN(n31700) );
  SDFFX1 \mem2_reg[5][19]  ( .D(n10455), .SI(\mem2[5][18] ), .SE(test_se), 
        .CLK(n2065), .Q(\mem2[5][19] ), .QN(n31701) );
  SDFFX1 \mem2_reg[5][18]  ( .D(n10454), .SI(\mem2[5][17] ), .SE(test_se), 
        .CLK(n2065), .Q(\mem2[5][18] ), .QN(n31702) );
  SDFFX1 \mem2_reg[5][17]  ( .D(n10453), .SI(\mem2[5][16] ), .SE(test_se), 
        .CLK(n2065), .Q(\mem2[5][17] ), .QN(n31703) );
  SDFFX1 \mem2_reg[5][16]  ( .D(n10452), .SI(\mem2[4][23] ), .SE(test_se), 
        .CLK(n2065), .Q(\mem2[5][16] ), .QN(n31704) );
  SDFFX1 \mem2_reg[4][23]  ( .D(n10451), .SI(\mem2[4][22] ), .SE(test_se), 
        .CLK(n2065), .Q(\mem2[4][23] ), .QN(n31705) );
  SDFFX1 \mem2_reg[4][22]  ( .D(n10450), .SI(\mem2[4][21] ), .SE(test_se), 
        .CLK(n2065), .Q(\mem2[4][22] ), .QN(n31706) );
  SDFFX1 \mem2_reg[4][21]  ( .D(n10449), .SI(\mem2[4][20] ), .SE(test_se), 
        .CLK(n2066), .Q(\mem2[4][21] ), .QN(n31707) );
  SDFFX1 \mem2_reg[4][20]  ( .D(n10448), .SI(\mem2[4][19] ), .SE(test_se), 
        .CLK(n2066), .Q(\mem2[4][20] ), .QN(n31708) );
  SDFFX1 \mem2_reg[4][19]  ( .D(n10447), .SI(\mem2[4][18] ), .SE(test_se), 
        .CLK(n2066), .Q(\mem2[4][19] ), .QN(n31709) );
  SDFFX1 \mem2_reg[4][18]  ( .D(n10446), .SI(test_si5), .SE(test_se), .CLK(
        n2066), .Q(\mem2[4][18] ), .QN(n31710) );
  SDFFX1 \mem2_reg[4][17]  ( .D(n10445), .SI(\mem2[4][16] ), .SE(test_se), 
        .CLK(n1407), .Q(\mem2[4][17] ), .QN(n31711) );
  SDFFX1 \mem2_reg[4][16]  ( .D(n10444), .SI(\mem2[3][23] ), .SE(test_se), 
        .CLK(n1407), .Q(\mem2[4][16] ), .QN(n31712) );
  SDFFX1 \mem2_reg[3][23]  ( .D(n10443), .SI(\mem2[3][22] ), .SE(test_se), 
        .CLK(n1407), .Q(\mem2[3][23] ), .QN(n31713) );
  SDFFX1 \mem2_reg[3][22]  ( .D(n10442), .SI(\mem2[3][21] ), .SE(test_se), 
        .CLK(n1407), .Q(\mem2[3][22] ), .QN(n31714) );
  SDFFX1 \mem2_reg[3][21]  ( .D(n10441), .SI(\mem2[3][20] ), .SE(test_se), 
        .CLK(n1408), .Q(\mem2[3][21] ), .QN(n31715) );
  SDFFX1 \mem2_reg[3][20]  ( .D(n10440), .SI(\mem2[3][19] ), .SE(test_se), 
        .CLK(n1408), .Q(\mem2[3][20] ), .QN(n31716) );
  SDFFX1 \mem2_reg[3][19]  ( .D(n10439), .SI(\mem2[3][18] ), .SE(test_se), 
        .CLK(n1408), .Q(\mem2[3][19] ), .QN(n31717) );
  SDFFX1 \mem2_reg[3][18]  ( .D(n10438), .SI(\mem2[3][17] ), .SE(test_se), 
        .CLK(n1408), .Q(\mem2[3][18] ), .QN(n31718) );
  SDFFX1 \mem2_reg[3][17]  ( .D(n10437), .SI(\mem2[3][16] ), .SE(test_se), 
        .CLK(n1408), .Q(\mem2[3][17] ), .QN(n31719) );
  SDFFX1 \mem2_reg[3][16]  ( .D(n10436), .SI(\mem2[2][23] ), .SE(test_se), 
        .CLK(n1408), .Q(\mem2[3][16] ), .QN(n31720) );
  SDFFX1 \mem2_reg[2][23]  ( .D(n10435), .SI(\mem2[2][22] ), .SE(test_se), 
        .CLK(n1408), .Q(\mem2[2][23] ), .QN(n31721) );
  SDFFX1 \mem2_reg[2][22]  ( .D(n10434), .SI(\mem2[2][21] ), .SE(test_se), 
        .CLK(n1408), .Q(\mem2[2][22] ), .QN(n31722) );
  SDFFX1 \mem2_reg[2][21]  ( .D(n10433), .SI(\mem2[2][20] ), .SE(test_se), 
        .CLK(n1408), .Q(\mem2[2][21] ), .QN(n31723) );
  SDFFX1 \mem2_reg[2][20]  ( .D(n10432), .SI(\mem2[2][19] ), .SE(test_se), 
        .CLK(n1408), .Q(\mem2[2][20] ), .QN(n31724) );
  SDFFX1 \mem2_reg[2][19]  ( .D(n10431), .SI(\mem2[2][18] ), .SE(test_se), 
        .CLK(n1408), .Q(\mem2[2][19] ), .QN(n31725) );
  SDFFX1 \mem2_reg[2][18]  ( .D(n10430), .SI(\mem2[2][17] ), .SE(test_se), 
        .CLK(n1408), .Q(\mem2[2][18] ), .QN(n31726) );
  SDFFX1 \mem2_reg[2][17]  ( .D(n10429), .SI(\mem2[2][16] ), .SE(test_se), 
        .CLK(n1409), .Q(\mem2[2][17] ), .QN(n31727) );
  SDFFX1 \mem2_reg[2][16]  ( .D(n10428), .SI(\mem2[1][23] ), .SE(test_se), 
        .CLK(n1409), .Q(\mem2[2][16] ), .QN(n31728) );
  SDFFX1 \mem2_reg[1][23]  ( .D(n10427), .SI(\mem2[1][22] ), .SE(test_se), 
        .CLK(n1409), .Q(\mem2[1][23] ), .QN(n31729) );
  SDFFX1 \mem2_reg[1][22]  ( .D(n10426), .SI(\mem2[1][21] ), .SE(test_se), 
        .CLK(n1409), .Q(\mem2[1][22] ), .QN(n31730) );
  SDFFX1 \mem2_reg[1][21]  ( .D(n10425), .SI(\mem2[1][20] ), .SE(test_se), 
        .CLK(n1409), .Q(\mem2[1][21] ), .QN(n31731) );
  SDFFX1 \mem2_reg[1][20]  ( .D(n10424), .SI(\mem2[1][19] ), .SE(test_se), 
        .CLK(n1409), .Q(\mem2[1][20] ), .QN(n31732) );
  SDFFX1 \mem2_reg[1][19]  ( .D(n10423), .SI(\mem2[1][18] ), .SE(test_se), 
        .CLK(n1409), .Q(\mem2[1][19] ), .QN(n31733) );
  SDFFX1 \mem2_reg[1][18]  ( .D(n10422), .SI(\mem2[1][17] ), .SE(test_se), 
        .CLK(n1409), .Q(\mem2[1][18] ), .QN(n31734) );
  SDFFX1 \mem2_reg[1][17]  ( .D(n10421), .SI(\mem2[1][16] ), .SE(test_se), 
        .CLK(n1409), .Q(\mem2[1][17] ), .QN(n31735) );
  SDFFX1 \mem2_reg[1][16]  ( .D(n10420), .SI(\mem2[0][23] ), .SE(test_se), 
        .CLK(n1409), .Q(\mem2[1][16] ), .QN(n31736) );
  SDFFX1 \mem2_reg[0][23]  ( .D(n10419), .SI(\mem2[0][22] ), .SE(test_se), 
        .CLK(n1409), .Q(\mem2[0][23] ), .QN(n31737) );
  SDFFX1 \mem2_reg[0][22]  ( .D(n10418), .SI(\mem2[0][21] ), .SE(test_se), 
        .CLK(n1409), .Q(\mem2[0][22] ), .QN(n31738) );
  SDFFX1 \mem2_reg[0][21]  ( .D(n10417), .SI(\mem2[0][20] ), .SE(test_se), 
        .CLK(n1410), .Q(\mem2[0][21] ), .QN(n31739) );
  SDFFX1 \mem2_reg[0][20]  ( .D(n10416), .SI(\mem2[0][19] ), .SE(test_se), 
        .CLK(n1410), .Q(\mem2[0][20] ), .QN(n31740) );
  SDFFX1 \mem2_reg[0][19]  ( .D(n10415), .SI(\mem2[0][18] ), .SE(test_se), 
        .CLK(n1410), .Q(\mem2[0][19] ), .QN(n31741) );
  SDFFX1 \mem2_reg[0][18]  ( .D(n10414), .SI(\mem2[0][17] ), .SE(test_se), 
        .CLK(n1410), .Q(\mem2[0][18] ), .QN(n31742) );
  SDFFX1 \mem2_reg[0][17]  ( .D(n10413), .SI(\mem2[0][16] ), .SE(test_se), 
        .CLK(n1410), .Q(\mem2[0][17] ), .QN(n31743) );
  SDFFX1 \mem2_reg[0][16]  ( .D(n10412), .SI(\mem1[255][15] ), .SE(test_se), 
        .CLK(n1410), .Q(\mem2[0][16] ), .QN(n31744) );
  BSLEX1 \do_tri[2]  ( .INOUT1(n2201), .ENB(n21510), .INOUT2(do[2]) );
  BSLEX1 \do_tri[3]  ( .INOUT1(n2200), .ENB(n21510), .INOUT2(do[3]) );
  BSLEX1 \do_tri[4]  ( .INOUT1(n2199), .ENB(n21510), .INOUT2(do[4]) );
  BSLEX1 \do_tri[5]  ( .INOUT1(n2198), .ENB(n21510), .INOUT2(do[5]) );
  BSLEX1 \do_tri[6]  ( .INOUT1(n2197), .ENB(n21510), .INOUT2(do[6]) );
  BSLEX1 \do_tri[7]  ( .INOUT1(n2196), .ENB(n21510), .INOUT2(do[7]) );
  BSLEX1 \do_tri[8]  ( .INOUT1(n2195), .ENB(n21510), .INOUT2(do[8]) );
  BSLEX1 \do_tri[9]  ( .INOUT1(n2193), .ENB(n21510), .INOUT2(do[9]) );
  BSLEX1 \do_tri[10]  ( .INOUT1(n2192), .ENB(n21510), .INOUT2(do[10]) );
  BSLEX1 \do_tri[11]  ( .INOUT1(n2191), .ENB(n21510), .INOUT2(do[11]) );
  BSLEX1 \do_tri[12]  ( .INOUT1(n2190), .ENB(n21510), .INOUT2(do[12]) );
  BSLEX1 \do_tri[0]  ( .INOUT1(n2203), .ENB(n21510), .INOUT2(do[0]) );
  BSLEX1 \do_tri[1]  ( .INOUT1(n2202), .ENB(n21510), .INOUT2(do[1]) );
  BSLEX1 \do_tri[15]  ( .INOUT1(n2187), .ENB(n21510), .INOUT2(do[15]) );
  BSLEX1 \do_tri[13]  ( .INOUT1(n2189), .ENB(n21510), .INOUT2(do[13]) );
  BSLEX1 \do_tri[14]  ( .INOUT1(n2188), .ENB(n21510), .INOUT2(do[14]) );
  BSLEX1 \do_tri[18]  ( .INOUT1(n2184), .ENB(n21510), .INOUT2(do[18]) );
  BSLEX1 \do_tri[17]  ( .INOUT1(n2185), .ENB(n21510), .INOUT2(do[17]) );
  BSLEX1 \do_tri[16]  ( .INOUT1(n2186), .ENB(n21510), .INOUT2(do[16]) );
  BSLEX1 \do_tri[19]  ( .INOUT1(n2183), .ENB(n21510), .INOUT2(do[19]) );
  BSLEX1 \do_tri[20]  ( .INOUT1(n2182), .ENB(n21510), .INOUT2(do[20]) );
  BSLEX1 \do_tri[31]  ( .INOUT1(n2171), .ENB(n21510), .INOUT2(do[31]) );
  BSLEX1 \do_tri[21]  ( .INOUT1(n2181), .ENB(n21510), .INOUT2(do[21]) );
  BSLEX1 \do_tri[23]  ( .INOUT1(n2179), .ENB(n21510), .INOUT2(do[23]) );
  BSLEX1 \do_tri[27]  ( .INOUT1(n2175), .ENB(n21510), .INOUT2(do[27]) );
  BSLEX1 \do_tri[30]  ( .INOUT1(n2172), .ENB(n21510), .INOUT2(do[30]) );
  BSLEX1 \do_tri[26]  ( .INOUT1(n2176), .ENB(n21510), .INOUT2(do[26]) );
  BSLEX1 \do_tri[25]  ( .INOUT1(n2177), .ENB(n21510), .INOUT2(do[25]) );
  BSLEX1 \do_tri[29]  ( .INOUT1(n2173), .ENB(n21510), .INOUT2(do[29]) );
  BSLEX1 \do_tri[28]  ( .INOUT1(n2174), .ENB(n21510), .INOUT2(do[28]) );
  BSLEX1 \do_tri[22]  ( .INOUT1(n2180), .ENB(n21510), .INOUT2(do[22]) );
  BSLEX1 \do_tri[24]  ( .INOUT1(n2178), .ENB(n21510), .INOUT2(do[24]) );
  NBUFFX2 U2 ( .INP(n2132), .Z(n1409) );
  NBUFFX2 U3 ( .INP(n2132), .Z(n1408) );
  NBUFFX2 U4 ( .INP(n2077), .Z(n2065) );
  NBUFFX2 U5 ( .INP(n2078), .Z(n2064) );
  NBUFFX2 U6 ( .INP(n2078), .Z(n2054) );
  NBUFFX2 U7 ( .INP(n2079), .Z(n2044) );
  NBUFFX2 U8 ( .INP(n2079), .Z(n2043) );
  NBUFFX2 U9 ( .INP(n2079), .Z(n2042) );
  NBUFFX2 U10 ( .INP(n2079), .Z(n2041) );
  NBUFFX2 U11 ( .INP(n2080), .Z(n2040) );
  NBUFFX2 U12 ( .INP(n2080), .Z(n2039) );
  NBUFFX2 U13 ( .INP(n2080), .Z(n2038) );
  NBUFFX2 U14 ( .INP(n2080), .Z(n2037) );
  NBUFFX2 U15 ( .INP(n2080), .Z(n2036) );
  NBUFFX2 U16 ( .INP(n2080), .Z(n2035) );
  NBUFFX2 U17 ( .INP(n2080), .Z(n2034) );
  NBUFFX2 U18 ( .INP(n2080), .Z(n2033) );
  NBUFFX2 U19 ( .INP(n2080), .Z(n2032) );
  NBUFFX2 U20 ( .INP(n2080), .Z(n2031) );
  NBUFFX2 U21 ( .INP(n2080), .Z(n2030) );
  NBUFFX2 U22 ( .INP(n2080), .Z(n2029) );
  NBUFFX2 U23 ( .INP(n2081), .Z(n2028) );
  NBUFFX2 U24 ( .INP(n2081), .Z(n2027) );
  NBUFFX2 U25 ( .INP(n2081), .Z(n2026) );
  NBUFFX2 U26 ( .INP(n2081), .Z(n2025) );
  NBUFFX2 U27 ( .INP(n2081), .Z(n2024) );
  NBUFFX2 U28 ( .INP(n2081), .Z(n2023) );
  NBUFFX2 U29 ( .INP(n2081), .Z(n2022) );
  NBUFFX2 U30 ( .INP(n2081), .Z(n2021) );
  NBUFFX2 U31 ( .INP(n2081), .Z(n2020) );
  NBUFFX2 U32 ( .INP(n2081), .Z(n2019) );
  NBUFFX2 U33 ( .INP(n2081), .Z(n2018) );
  NBUFFX2 U34 ( .INP(n2081), .Z(n2017) );
  NBUFFX2 U35 ( .INP(n2082), .Z(n2016) );
  NBUFFX2 U36 ( .INP(n2082), .Z(n2015) );
  NBUFFX2 U37 ( .INP(n2082), .Z(n2014) );
  NBUFFX2 U38 ( .INP(n2082), .Z(n2013) );
  NBUFFX2 U39 ( .INP(n2082), .Z(n2012) );
  NBUFFX2 U40 ( .INP(n2082), .Z(n2011) );
  NBUFFX2 U41 ( .INP(n2082), .Z(n2010) );
  NBUFFX2 U42 ( .INP(n2082), .Z(n2009) );
  NBUFFX2 U43 ( .INP(n2082), .Z(n2008) );
  NBUFFX2 U44 ( .INP(n2082), .Z(n2007) );
  NBUFFX2 U45 ( .INP(n2082), .Z(n2006) );
  NBUFFX2 U46 ( .INP(n2082), .Z(n2005) );
  NBUFFX2 U47 ( .INP(n2083), .Z(n2004) );
  NBUFFX2 U48 ( .INP(n2083), .Z(n2003) );
  NBUFFX2 U49 ( .INP(n2083), .Z(n2002) );
  NBUFFX2 U50 ( .INP(n2083), .Z(n2001) );
  NBUFFX2 U51 ( .INP(n2083), .Z(n2000) );
  NBUFFX2 U52 ( .INP(n2083), .Z(n1999) );
  NBUFFX2 U53 ( .INP(n2083), .Z(n1998) );
  NBUFFX2 U54 ( .INP(n2083), .Z(n1997) );
  NBUFFX2 U55 ( .INP(n2083), .Z(n1996) );
  NBUFFX2 U56 ( .INP(n2083), .Z(n1995) );
  NBUFFX2 U57 ( .INP(n2083), .Z(n1994) );
  NBUFFX2 U58 ( .INP(n2083), .Z(n1993) );
  NBUFFX2 U59 ( .INP(n2084), .Z(n1992) );
  NBUFFX2 U60 ( .INP(n2084), .Z(n1991) );
  NBUFFX2 U61 ( .INP(n2084), .Z(n1990) );
  NBUFFX2 U62 ( .INP(n2084), .Z(n1989) );
  NBUFFX2 U63 ( .INP(n2084), .Z(n1988) );
  NBUFFX2 U64 ( .INP(n2084), .Z(n1987) );
  NBUFFX2 U65 ( .INP(n2084), .Z(n1986) );
  NBUFFX2 U66 ( .INP(n2084), .Z(n1985) );
  NBUFFX2 U67 ( .INP(n2084), .Z(n1984) );
  NBUFFX2 U68 ( .INP(n2084), .Z(n1983) );
  NBUFFX2 U69 ( .INP(n2084), .Z(n1982) );
  NBUFFX2 U70 ( .INP(n2084), .Z(n1981) );
  NBUFFX2 U71 ( .INP(n2085), .Z(n1980) );
  NBUFFX2 U72 ( .INP(n2085), .Z(n1979) );
  NBUFFX2 U73 ( .INP(n2085), .Z(n1978) );
  NBUFFX2 U74 ( .INP(n2085), .Z(n1977) );
  NBUFFX2 U75 ( .INP(n2085), .Z(n1976) );
  NBUFFX2 U76 ( .INP(n2085), .Z(n1975) );
  NBUFFX2 U77 ( .INP(n2085), .Z(n1974) );
  NBUFFX2 U78 ( .INP(n2085), .Z(n1973) );
  NBUFFX2 U79 ( .INP(n2085), .Z(n1972) );
  NBUFFX2 U80 ( .INP(n2085), .Z(n1971) );
  NBUFFX2 U81 ( .INP(n2085), .Z(n1970) );
  NBUFFX2 U82 ( .INP(n2085), .Z(n1969) );
  NBUFFX2 U83 ( .INP(n2086), .Z(n1968) );
  NBUFFX2 U84 ( .INP(n2086), .Z(n1967) );
  NBUFFX2 U85 ( .INP(n2086), .Z(n1966) );
  NBUFFX2 U86 ( .INP(n2086), .Z(n1965) );
  NBUFFX2 U87 ( .INP(n2086), .Z(n1964) );
  NBUFFX2 U88 ( .INP(n2086), .Z(n1963) );
  NBUFFX2 U89 ( .INP(n2086), .Z(n1962) );
  NBUFFX2 U90 ( .INP(n2086), .Z(n1961) );
  NBUFFX2 U91 ( .INP(n2086), .Z(n1960) );
  NBUFFX2 U92 ( .INP(n2086), .Z(n1959) );
  NBUFFX2 U93 ( .INP(n2086), .Z(n1958) );
  NBUFFX2 U94 ( .INP(n2086), .Z(n1957) );
  NBUFFX2 U95 ( .INP(n2087), .Z(n1956) );
  NBUFFX2 U96 ( .INP(n2087), .Z(n1955) );
  NBUFFX2 U97 ( .INP(n2087), .Z(n1954) );
  NBUFFX2 U98 ( .INP(n2087), .Z(n1953) );
  NBUFFX2 U99 ( .INP(n2087), .Z(n1952) );
  NBUFFX2 U100 ( .INP(n2087), .Z(n1951) );
  NBUFFX2 U101 ( .INP(n2087), .Z(n1950) );
  NBUFFX2 U102 ( .INP(n2087), .Z(n1949) );
  NBUFFX2 U103 ( .INP(n2087), .Z(n1948) );
  NBUFFX2 U104 ( .INP(n2087), .Z(n1947) );
  NBUFFX2 U105 ( .INP(n2087), .Z(n1946) );
  NBUFFX2 U106 ( .INP(n2087), .Z(n1945) );
  NBUFFX2 U107 ( .INP(n2088), .Z(n1944) );
  NBUFFX2 U108 ( .INP(n2088), .Z(n1943) );
  NBUFFX2 U109 ( .INP(n2088), .Z(n1942) );
  NBUFFX2 U110 ( .INP(n2088), .Z(n1941) );
  NBUFFX2 U111 ( .INP(n2088), .Z(n1940) );
  NBUFFX2 U112 ( .INP(n2088), .Z(n1939) );
  NBUFFX2 U113 ( .INP(n2088), .Z(n1938) );
  NBUFFX2 U114 ( .INP(n2088), .Z(n1937) );
  NBUFFX2 U115 ( .INP(n2088), .Z(n1936) );
  NBUFFX2 U116 ( .INP(n2088), .Z(n1935) );
  NBUFFX2 U117 ( .INP(n2088), .Z(n1934) );
  NBUFFX2 U118 ( .INP(n2088), .Z(n1933) );
  NBUFFX2 U119 ( .INP(n2089), .Z(n1932) );
  NBUFFX2 U120 ( .INP(n2089), .Z(n1931) );
  NBUFFX2 U121 ( .INP(n2089), .Z(n1930) );
  NBUFFX2 U122 ( .INP(n2089), .Z(n1929) );
  NBUFFX2 U123 ( .INP(n2089), .Z(n1928) );
  NBUFFX2 U124 ( .INP(n2089), .Z(n1927) );
  NBUFFX2 U125 ( .INP(n2089), .Z(n1926) );
  NBUFFX2 U126 ( .INP(n2089), .Z(n1925) );
  NBUFFX2 U127 ( .INP(n2089), .Z(n1924) );
  NBUFFX2 U128 ( .INP(n2089), .Z(n1923) );
  NBUFFX2 U129 ( .INP(n2089), .Z(n1922) );
  NBUFFX2 U130 ( .INP(n2089), .Z(n1921) );
  NBUFFX2 U131 ( .INP(n2090), .Z(n1920) );
  NBUFFX2 U132 ( .INP(n2090), .Z(n1919) );
  NBUFFX2 U133 ( .INP(n2090), .Z(n1918) );
  NBUFFX2 U134 ( .INP(n2090), .Z(n1917) );
  NBUFFX2 U135 ( .INP(n2090), .Z(n1916) );
  NBUFFX2 U136 ( .INP(n2090), .Z(n1915) );
  NBUFFX2 U137 ( .INP(n2090), .Z(n1914) );
  NBUFFX2 U138 ( .INP(n2090), .Z(n1913) );
  NBUFFX2 U139 ( .INP(n2090), .Z(n1912) );
  NBUFFX2 U140 ( .INP(n2090), .Z(n1911) );
  NBUFFX2 U141 ( .INP(n2090), .Z(n1910) );
  NBUFFX2 U142 ( .INP(n2090), .Z(n1909) );
  NBUFFX2 U143 ( .INP(n2091), .Z(n1908) );
  NBUFFX2 U144 ( .INP(n2091), .Z(n1907) );
  NBUFFX2 U145 ( .INP(n2091), .Z(n1906) );
  NBUFFX2 U146 ( .INP(n2091), .Z(n1905) );
  NBUFFX2 U147 ( .INP(n2091), .Z(n1904) );
  NBUFFX2 U148 ( .INP(n2091), .Z(n1903) );
  NBUFFX2 U149 ( .INP(n2091), .Z(n1902) );
  NBUFFX2 U150 ( .INP(n2091), .Z(n1901) );
  NBUFFX2 U151 ( .INP(n2091), .Z(n1900) );
  NBUFFX2 U152 ( .INP(n2091), .Z(n1899) );
  NBUFFX2 U153 ( .INP(n2091), .Z(n1898) );
  NBUFFX2 U154 ( .INP(n2091), .Z(n1897) );
  NBUFFX2 U155 ( .INP(n2092), .Z(n1896) );
  NBUFFX2 U156 ( .INP(n2092), .Z(n1895) );
  NBUFFX2 U157 ( .INP(n2092), .Z(n1894) );
  NBUFFX2 U158 ( .INP(n2092), .Z(n1893) );
  NBUFFX2 U159 ( .INP(n2092), .Z(n1892) );
  NBUFFX2 U160 ( .INP(n2092), .Z(n1891) );
  NBUFFX2 U161 ( .INP(n2092), .Z(n1890) );
  NBUFFX2 U162 ( .INP(n2092), .Z(n1889) );
  NBUFFX2 U163 ( .INP(n2092), .Z(n1888) );
  NBUFFX2 U164 ( .INP(n2092), .Z(n1887) );
  NBUFFX2 U165 ( .INP(n2092), .Z(n1886) );
  NBUFFX2 U166 ( .INP(n2092), .Z(n1885) );
  NBUFFX2 U167 ( .INP(n2077), .Z(n2070) );
  NBUFFX2 U168 ( .INP(n2077), .Z(n2069) );
  NBUFFX2 U169 ( .INP(n2078), .Z(n2063) );
  NBUFFX2 U170 ( .INP(n2078), .Z(n2062) );
  NBUFFX2 U171 ( .INP(n2078), .Z(n2053) );
  NBUFFX2 U172 ( .INP(n2079), .Z(n2052) );
  NBUFFX2 U173 ( .INP(n2079), .Z(n2051) );
  NBUFFX2 U174 ( .INP(n2093), .Z(n1884) );
  NBUFFX2 U175 ( .INP(n2093), .Z(n1883) );
  NBUFFX2 U176 ( .INP(n2093), .Z(n1882) );
  NBUFFX2 U177 ( .INP(n2093), .Z(n1881) );
  NBUFFX2 U178 ( .INP(n2093), .Z(n1880) );
  NBUFFX2 U179 ( .INP(n2093), .Z(n1879) );
  NBUFFX2 U180 ( .INP(n2093), .Z(n1878) );
  NBUFFX2 U181 ( .INP(n2093), .Z(n1877) );
  NBUFFX2 U182 ( .INP(n2093), .Z(n1876) );
  NBUFFX2 U183 ( .INP(n2093), .Z(n1875) );
  NBUFFX2 U184 ( .INP(n2093), .Z(n1874) );
  NBUFFX2 U185 ( .INP(n2093), .Z(n1873) );
  NBUFFX2 U186 ( .INP(n2094), .Z(n1872) );
  NBUFFX2 U187 ( .INP(n2094), .Z(n1871) );
  NBUFFX2 U188 ( .INP(n2094), .Z(n1870) );
  NBUFFX2 U189 ( .INP(n2094), .Z(n1869) );
  NBUFFX2 U190 ( .INP(n2094), .Z(n1868) );
  NBUFFX2 U191 ( .INP(n2094), .Z(n1867) );
  NBUFFX2 U192 ( .INP(n2094), .Z(n1866) );
  NBUFFX2 U193 ( .INP(n2094), .Z(n1865) );
  NBUFFX2 U194 ( .INP(n2094), .Z(n1864) );
  NBUFFX2 U195 ( .INP(n2094), .Z(n1863) );
  NBUFFX2 U196 ( .INP(n2094), .Z(n1862) );
  NBUFFX2 U197 ( .INP(n2094), .Z(n1861) );
  NBUFFX2 U198 ( .INP(n2095), .Z(n1860) );
  NBUFFX2 U199 ( .INP(n2095), .Z(n1859) );
  NBUFFX2 U200 ( .INP(n2095), .Z(n1858) );
  NBUFFX2 U201 ( .INP(n2095), .Z(n1857) );
  NBUFFX2 U202 ( .INP(n2095), .Z(n1856) );
  NBUFFX2 U203 ( .INP(n2095), .Z(n1855) );
  NBUFFX2 U204 ( .INP(n2095), .Z(n1854) );
  NBUFFX2 U205 ( .INP(n2095), .Z(n1853) );
  NBUFFX2 U206 ( .INP(n2095), .Z(n1852) );
  NBUFFX2 U207 ( .INP(n2095), .Z(n1851) );
  NBUFFX2 U208 ( .INP(n2095), .Z(n1850) );
  NBUFFX2 U209 ( .INP(n2095), .Z(n1849) );
  NBUFFX2 U210 ( .INP(n2096), .Z(n1848) );
  NBUFFX2 U211 ( .INP(n2096), .Z(n1847) );
  NBUFFX2 U212 ( .INP(n2096), .Z(n1846) );
  NBUFFX2 U213 ( .INP(n2096), .Z(n1845) );
  NBUFFX2 U214 ( .INP(n2096), .Z(n1844) );
  NBUFFX2 U215 ( .INP(n2096), .Z(n1843) );
  NBUFFX2 U216 ( .INP(n2096), .Z(n1842) );
  NBUFFX2 U217 ( .INP(n2096), .Z(n1841) );
  NBUFFX2 U218 ( .INP(n2077), .Z(n2074) );
  NBUFFX2 U219 ( .INP(n2077), .Z(n2071) );
  NBUFFX2 U220 ( .INP(n2077), .Z(n2068) );
  NBUFFX2 U221 ( .INP(n2077), .Z(n2067) );
  NBUFFX2 U222 ( .INP(n2077), .Z(n2066) );
  NBUFFX2 U223 ( .INP(n2078), .Z(n2061) );
  NBUFFX2 U224 ( .INP(n2078), .Z(n2060) );
  NBUFFX2 U225 ( .INP(n2078), .Z(n2059) );
  NBUFFX2 U226 ( .INP(n2079), .Z(n2050) );
  NBUFFX2 U227 ( .INP(n2079), .Z(n2049) );
  NBUFFX2 U228 ( .INP(n2079), .Z(n2048) );
  NBUFFX2 U229 ( .INP(n2096), .Z(n1840) );
  NBUFFX2 U230 ( .INP(n2096), .Z(n1839) );
  NBUFFX2 U231 ( .INP(n2096), .Z(n1838) );
  NBUFFX2 U232 ( .INP(n2096), .Z(n1837) );
  NBUFFX2 U233 ( .INP(n2097), .Z(n1836) );
  NBUFFX2 U234 ( .INP(n2097), .Z(n1835) );
  NBUFFX2 U235 ( .INP(n2097), .Z(n1834) );
  NBUFFX2 U236 ( .INP(n2097), .Z(n1833) );
  NBUFFX2 U237 ( .INP(n2097), .Z(n1832) );
  NBUFFX2 U238 ( .INP(n2097), .Z(n1831) );
  NBUFFX2 U239 ( .INP(n2097), .Z(n1830) );
  NBUFFX2 U240 ( .INP(n2097), .Z(n1829) );
  NBUFFX2 U241 ( .INP(n2097), .Z(n1828) );
  NBUFFX2 U242 ( .INP(n2097), .Z(n1827) );
  NBUFFX2 U243 ( .INP(n2097), .Z(n1826) );
  NBUFFX2 U244 ( .INP(n2097), .Z(n1825) );
  NBUFFX2 U245 ( .INP(n2098), .Z(n1824) );
  NBUFFX2 U246 ( .INP(n2098), .Z(n1823) );
  NBUFFX2 U247 ( .INP(n2098), .Z(n1822) );
  NBUFFX2 U248 ( .INP(n2098), .Z(n1821) );
  NBUFFX2 U249 ( .INP(n2098), .Z(n1820) );
  NBUFFX2 U250 ( .INP(n2098), .Z(n1819) );
  NBUFFX2 U251 ( .INP(n2098), .Z(n1818) );
  NBUFFX2 U252 ( .INP(n2098), .Z(n1817) );
  NBUFFX2 U253 ( .INP(n2098), .Z(n1816) );
  NBUFFX2 U254 ( .INP(n2098), .Z(n1815) );
  NBUFFX2 U255 ( .INP(n2098), .Z(n1814) );
  NBUFFX2 U256 ( .INP(n2098), .Z(n1813) );
  NBUFFX2 U257 ( .INP(n2099), .Z(n1812) );
  NBUFFX2 U258 ( .INP(n2099), .Z(n1811) );
  NBUFFX2 U259 ( .INP(n2099), .Z(n1810) );
  NBUFFX2 U260 ( .INP(n2099), .Z(n1809) );
  NBUFFX2 U261 ( .INP(n2099), .Z(n1808) );
  NBUFFX2 U262 ( .INP(n2099), .Z(n1807) );
  NBUFFX2 U263 ( .INP(n2099), .Z(n1806) );
  NBUFFX2 U264 ( .INP(n2099), .Z(n1805) );
  NBUFFX2 U265 ( .INP(n2099), .Z(n1804) );
  NBUFFX2 U266 ( .INP(n2099), .Z(n1803) );
  NBUFFX2 U267 ( .INP(n2099), .Z(n1802) );
  NBUFFX2 U268 ( .INP(n2099), .Z(n1801) );
  NBUFFX2 U269 ( .INP(n2100), .Z(n1800) );
  NBUFFX2 U270 ( .INP(n2100), .Z(n1799) );
  NBUFFX2 U271 ( .INP(n2100), .Z(n1798) );
  NBUFFX2 U272 ( .INP(n2100), .Z(n1797) );
  NBUFFX2 U273 ( .INP(n2100), .Z(n1796) );
  NBUFFX2 U274 ( .INP(n2100), .Z(n1795) );
  NBUFFX2 U275 ( .INP(n2100), .Z(n1794) );
  NBUFFX2 U276 ( .INP(n2100), .Z(n1793) );
  NBUFFX2 U277 ( .INP(n2100), .Z(n1792) );
  NBUFFX2 U278 ( .INP(n2100), .Z(n1791) );
  NBUFFX2 U279 ( .INP(n2100), .Z(n1790) );
  NBUFFX2 U280 ( .INP(n2100), .Z(n1789) );
  NBUFFX2 U281 ( .INP(n2101), .Z(n1788) );
  NBUFFX2 U282 ( .INP(n2101), .Z(n1787) );
  NBUFFX2 U283 ( .INP(n2101), .Z(n1786) );
  NBUFFX2 U284 ( .INP(n2101), .Z(n1785) );
  NBUFFX2 U285 ( .INP(n2101), .Z(n1784) );
  NBUFFX2 U286 ( .INP(n2101), .Z(n1783) );
  NBUFFX2 U287 ( .INP(n2101), .Z(n1782) );
  NBUFFX2 U288 ( .INP(n2101), .Z(n1781) );
  NBUFFX2 U289 ( .INP(n2101), .Z(n1780) );
  NBUFFX2 U290 ( .INP(n2101), .Z(n1779) );
  NBUFFX2 U291 ( .INP(n2101), .Z(n1778) );
  NBUFFX2 U292 ( .INP(n2101), .Z(n1777) );
  NBUFFX2 U293 ( .INP(n2102), .Z(n1776) );
  NBUFFX2 U294 ( .INP(n2102), .Z(n1775) );
  NBUFFX2 U295 ( .INP(n2102), .Z(n1774) );
  NBUFFX2 U296 ( .INP(n2102), .Z(n1773) );
  NBUFFX2 U297 ( .INP(n2102), .Z(n1772) );
  NBUFFX2 U298 ( .INP(n2102), .Z(n1771) );
  NBUFFX2 U299 ( .INP(n2102), .Z(n1770) );
  NBUFFX2 U300 ( .INP(n2102), .Z(n1769) );
  NBUFFX2 U301 ( .INP(n2102), .Z(n1768) );
  NBUFFX2 U302 ( .INP(n2102), .Z(n1767) );
  NBUFFX2 U303 ( .INP(n2102), .Z(n1766) );
  NBUFFX2 U304 ( .INP(n2102), .Z(n1765) );
  NBUFFX2 U305 ( .INP(n2103), .Z(n1764) );
  NBUFFX2 U306 ( .INP(n2103), .Z(n1763) );
  NBUFFX2 U307 ( .INP(n2103), .Z(n1762) );
  NBUFFX2 U308 ( .INP(n2103), .Z(n1761) );
  NBUFFX2 U309 ( .INP(n2103), .Z(n1760) );
  NBUFFX2 U310 ( .INP(n2103), .Z(n1759) );
  NBUFFX2 U311 ( .INP(n2103), .Z(n1758) );
  NBUFFX2 U312 ( .INP(n2103), .Z(n1757) );
  NBUFFX2 U313 ( .INP(n2103), .Z(n1756) );
  NBUFFX2 U314 ( .INP(n2103), .Z(n1755) );
  NBUFFX2 U315 ( .INP(n2103), .Z(n1754) );
  NBUFFX2 U316 ( .INP(n2103), .Z(n1753) );
  NBUFFX2 U317 ( .INP(n2104), .Z(n1752) );
  NBUFFX2 U318 ( .INP(n2104), .Z(n1751) );
  NBUFFX2 U319 ( .INP(n2104), .Z(n1750) );
  NBUFFX2 U320 ( .INP(n2104), .Z(n1749) );
  NBUFFX2 U321 ( .INP(n2104), .Z(n1748) );
  NBUFFX2 U322 ( .INP(n2104), .Z(n1747) );
  NBUFFX2 U323 ( .INP(n2104), .Z(n1746) );
  NBUFFX2 U324 ( .INP(n2104), .Z(n1745) );
  NBUFFX2 U325 ( .INP(n2104), .Z(n1744) );
  NBUFFX2 U326 ( .INP(n2104), .Z(n1743) );
  NBUFFX2 U327 ( .INP(n2104), .Z(n1742) );
  NBUFFX2 U328 ( .INP(n2104), .Z(n1741) );
  NBUFFX2 U329 ( .INP(n2077), .Z(n2075) );
  NBUFFX2 U330 ( .INP(n2077), .Z(n2073) );
  NBUFFX2 U331 ( .INP(n2077), .Z(n2072) );
  NBUFFX2 U332 ( .INP(n2078), .Z(n2058) );
  NBUFFX2 U333 ( .INP(n2078), .Z(n2057) );
  NBUFFX2 U334 ( .INP(n2078), .Z(n2056) );
  NBUFFX2 U335 ( .INP(n2078), .Z(n2055) );
  NBUFFX2 U336 ( .INP(n2079), .Z(n2047) );
  NBUFFX2 U337 ( .INP(n2079), .Z(n2046) );
  NBUFFX2 U338 ( .INP(n2079), .Z(n2045) );
  NBUFFX2 U339 ( .INP(n2105), .Z(n1740) );
  NBUFFX2 U340 ( .INP(n2105), .Z(n1739) );
  NBUFFX2 U341 ( .INP(n2105), .Z(n1738) );
  NBUFFX2 U342 ( .INP(n2118), .Z(n1580) );
  NBUFFX2 U343 ( .INP(n2118), .Z(n1579) );
  NBUFFX2 U344 ( .INP(n2118), .Z(n1578) );
  NBUFFX2 U345 ( .INP(n2118), .Z(n1577) );
  NBUFFX2 U346 ( .INP(n2118), .Z(n1576) );
  NBUFFX2 U347 ( .INP(n2118), .Z(n1575) );
  NBUFFX2 U348 ( .INP(n2118), .Z(n1574) );
  NBUFFX2 U349 ( .INP(n2118), .Z(n1573) );
  NBUFFX2 U350 ( .INP(n2119), .Z(n1572) );
  NBUFFX2 U351 ( .INP(n2119), .Z(n1571) );
  NBUFFX2 U352 ( .INP(n2119), .Z(n1570) );
  NBUFFX2 U353 ( .INP(n2119), .Z(n1569) );
  NBUFFX2 U354 ( .INP(n2119), .Z(n1568) );
  NBUFFX2 U355 ( .INP(n2119), .Z(n1567) );
  NBUFFX2 U356 ( .INP(n2119), .Z(n1566) );
  NBUFFX2 U357 ( .INP(n2119), .Z(n1565) );
  NBUFFX2 U358 ( .INP(n2119), .Z(n1564) );
  NBUFFX2 U359 ( .INP(n2119), .Z(n1563) );
  NBUFFX2 U360 ( .INP(n2119), .Z(n1562) );
  NBUFFX2 U361 ( .INP(n2119), .Z(n1561) );
  NBUFFX2 U362 ( .INP(n2120), .Z(n1560) );
  NBUFFX2 U363 ( .INP(n2120), .Z(n1559) );
  NBUFFX2 U364 ( .INP(n2120), .Z(n1558) );
  NBUFFX2 U365 ( .INP(n2120), .Z(n1557) );
  NBUFFX2 U366 ( .INP(n2120), .Z(n1556) );
  NBUFFX2 U367 ( .INP(n2120), .Z(n1555) );
  NBUFFX2 U368 ( .INP(n2120), .Z(n1554) );
  NBUFFX2 U369 ( .INP(n2120), .Z(n1553) );
  NBUFFX2 U370 ( .INP(n2120), .Z(n1552) );
  NBUFFX2 U371 ( .INP(n2120), .Z(n1551) );
  NBUFFX2 U372 ( .INP(n2120), .Z(n1550) );
  NBUFFX2 U373 ( .INP(n2120), .Z(n1549) );
  NBUFFX2 U374 ( .INP(n2121), .Z(n1548) );
  NBUFFX2 U375 ( .INP(n2121), .Z(n1547) );
  NBUFFX2 U376 ( .INP(n2121), .Z(n1546) );
  NBUFFX2 U377 ( .INP(n2121), .Z(n1545) );
  NBUFFX2 U378 ( .INP(n2121), .Z(n1544) );
  NBUFFX2 U379 ( .INP(n2121), .Z(n1543) );
  NBUFFX2 U380 ( .INP(n2121), .Z(n1542) );
  NBUFFX2 U381 ( .INP(n2121), .Z(n1541) );
  NBUFFX2 U382 ( .INP(n2121), .Z(n1540) );
  NBUFFX2 U383 ( .INP(n2121), .Z(n1539) );
  NBUFFX2 U384 ( .INP(n2121), .Z(n1538) );
  NBUFFX2 U385 ( .INP(n2121), .Z(n1537) );
  NBUFFX2 U386 ( .INP(n2122), .Z(n1536) );
  NBUFFX2 U387 ( .INP(n2122), .Z(n1535) );
  NBUFFX2 U388 ( .INP(n2122), .Z(n1534) );
  NBUFFX2 U389 ( .INP(n2122), .Z(n1533) );
  NBUFFX2 U390 ( .INP(n2122), .Z(n1532) );
  NBUFFX2 U391 ( .INP(n2122), .Z(n1531) );
  NBUFFX2 U392 ( .INP(n2122), .Z(n1530) );
  NBUFFX2 U393 ( .INP(n2122), .Z(n1529) );
  NBUFFX2 U394 ( .INP(n2122), .Z(n1528) );
  NBUFFX2 U395 ( .INP(n2122), .Z(n1527) );
  NBUFFX2 U396 ( .INP(n2122), .Z(n1526) );
  NBUFFX2 U397 ( .INP(n2122), .Z(n1525) );
  NBUFFX2 U398 ( .INP(n2123), .Z(n1524) );
  NBUFFX2 U399 ( .INP(n2123), .Z(n1523) );
  NBUFFX2 U400 ( .INP(n2123), .Z(n1522) );
  NBUFFX2 U401 ( .INP(n2123), .Z(n1521) );
  NBUFFX2 U402 ( .INP(n2123), .Z(n1520) );
  NBUFFX2 U403 ( .INP(n2123), .Z(n1519) );
  NBUFFX2 U404 ( .INP(n2123), .Z(n1518) );
  NBUFFX2 U405 ( .INP(n2123), .Z(n1517) );
  NBUFFX2 U406 ( .INP(n2123), .Z(n1516) );
  NBUFFX2 U407 ( .INP(n2123), .Z(n1515) );
  NBUFFX2 U408 ( .INP(n2123), .Z(n1514) );
  NBUFFX2 U409 ( .INP(n2123), .Z(n1513) );
  NBUFFX2 U410 ( .INP(n2124), .Z(n1512) );
  NBUFFX2 U411 ( .INP(n2124), .Z(n1511) );
  NBUFFX2 U412 ( .INP(n2124), .Z(n1510) );
  NBUFFX2 U413 ( .INP(n2124), .Z(n1509) );
  NBUFFX2 U414 ( .INP(n2124), .Z(n1508) );
  NBUFFX2 U415 ( .INP(n2124), .Z(n1507) );
  NBUFFX2 U416 ( .INP(n2124), .Z(n1506) );
  NBUFFX2 U417 ( .INP(n2124), .Z(n1505) );
  NBUFFX2 U418 ( .INP(n2124), .Z(n1504) );
  NBUFFX2 U419 ( .INP(n2124), .Z(n1503) );
  NBUFFX2 U420 ( .INP(n2124), .Z(n1502) );
  NBUFFX2 U421 ( .INP(n2124), .Z(n1501) );
  NBUFFX2 U422 ( .INP(n2125), .Z(n1500) );
  NBUFFX2 U423 ( .INP(n2125), .Z(n1499) );
  NBUFFX2 U424 ( .INP(n2125), .Z(n1498) );
  NBUFFX2 U425 ( .INP(n2125), .Z(n1497) );
  NBUFFX2 U426 ( .INP(n2125), .Z(n1496) );
  NBUFFX2 U427 ( .INP(n2125), .Z(n1495) );
  NBUFFX2 U428 ( .INP(n2125), .Z(n1494) );
  NBUFFX2 U429 ( .INP(n2125), .Z(n1493) );
  NBUFFX2 U430 ( .INP(n2125), .Z(n1492) );
  NBUFFX2 U431 ( .INP(n2125), .Z(n1491) );
  NBUFFX2 U432 ( .INP(n2125), .Z(n1490) );
  NBUFFX2 U433 ( .INP(n2125), .Z(n1489) );
  NBUFFX2 U434 ( .INP(n2126), .Z(n1488) );
  NBUFFX2 U435 ( .INP(n2126), .Z(n1487) );
  NBUFFX2 U436 ( .INP(n2126), .Z(n1486) );
  NBUFFX2 U437 ( .INP(n2126), .Z(n1485) );
  NBUFFX2 U438 ( .INP(n2126), .Z(n1484) );
  NBUFFX2 U439 ( .INP(n2126), .Z(n1483) );
  NBUFFX2 U440 ( .INP(n2126), .Z(n1482) );
  NBUFFX2 U441 ( .INP(n2126), .Z(n1481) );
  NBUFFX2 U442 ( .INP(n2126), .Z(n1480) );
  NBUFFX2 U443 ( .INP(n2126), .Z(n1479) );
  NBUFFX2 U444 ( .INP(n2126), .Z(n1478) );
  NBUFFX2 U445 ( .INP(n2126), .Z(n1477) );
  NBUFFX2 U446 ( .INP(n2127), .Z(n1476) );
  NBUFFX2 U447 ( .INP(n2127), .Z(n1475) );
  NBUFFX2 U448 ( .INP(n2127), .Z(n1474) );
  NBUFFX2 U449 ( .INP(n2127), .Z(n1473) );
  NBUFFX2 U450 ( .INP(n2127), .Z(n1472) );
  NBUFFX2 U451 ( .INP(n2127), .Z(n1471) );
  NBUFFX2 U452 ( .INP(n2127), .Z(n1470) );
  NBUFFX2 U453 ( .INP(n2127), .Z(n1469) );
  NBUFFX2 U454 ( .INP(n2127), .Z(n1468) );
  NBUFFX2 U455 ( .INP(n2127), .Z(n1467) );
  NBUFFX2 U456 ( .INP(n2127), .Z(n1466) );
  NBUFFX2 U457 ( .INP(n2127), .Z(n1465) );
  NBUFFX2 U458 ( .INP(n2128), .Z(n1464) );
  NBUFFX2 U459 ( .INP(n2128), .Z(n1463) );
  NBUFFX2 U460 ( .INP(n2128), .Z(n1462) );
  NBUFFX2 U461 ( .INP(n2128), .Z(n1461) );
  NBUFFX2 U462 ( .INP(n2128), .Z(n1460) );
  NBUFFX2 U463 ( .INP(n2128), .Z(n1459) );
  NBUFFX2 U464 ( .INP(n2128), .Z(n1458) );
  NBUFFX2 U465 ( .INP(n2128), .Z(n1457) );
  NBUFFX2 U466 ( .INP(n2128), .Z(n1456) );
  NBUFFX2 U467 ( .INP(n2128), .Z(n1455) );
  NBUFFX2 U468 ( .INP(n2128), .Z(n1454) );
  NBUFFX2 U469 ( .INP(n2128), .Z(n1453) );
  NBUFFX2 U470 ( .INP(n2129), .Z(n1452) );
  NBUFFX2 U471 ( .INP(n2129), .Z(n1451) );
  NBUFFX2 U472 ( .INP(n2129), .Z(n1450) );
  NBUFFX2 U473 ( .INP(n2129), .Z(n1449) );
  NBUFFX2 U474 ( .INP(n2129), .Z(n1448) );
  NBUFFX2 U475 ( .INP(n2129), .Z(n1447) );
  NBUFFX2 U476 ( .INP(n2129), .Z(n1446) );
  NBUFFX2 U477 ( .INP(n2129), .Z(n1445) );
  NBUFFX2 U478 ( .INP(n2129), .Z(n1444) );
  NBUFFX2 U479 ( .INP(n2129), .Z(n1443) );
  NBUFFX2 U480 ( .INP(n2129), .Z(n1442) );
  NBUFFX2 U481 ( .INP(n2129), .Z(n1441) );
  NBUFFX2 U482 ( .INP(n2130), .Z(n1440) );
  NBUFFX2 U483 ( .INP(n2130), .Z(n1439) );
  NBUFFX2 U484 ( .INP(n2130), .Z(n1438) );
  NBUFFX2 U485 ( .INP(n2130), .Z(n1437) );
  NBUFFX2 U486 ( .INP(n2130), .Z(n1436) );
  NBUFFX2 U487 ( .INP(n2130), .Z(n1435) );
  NBUFFX2 U488 ( .INP(n2130), .Z(n1434) );
  NBUFFX2 U489 ( .INP(n2130), .Z(n1433) );
  NBUFFX2 U490 ( .INP(n2130), .Z(n1432) );
  NBUFFX2 U491 ( .INP(n2130), .Z(n1431) );
  NBUFFX2 U492 ( .INP(n2130), .Z(n1430) );
  NBUFFX2 U493 ( .INP(n2130), .Z(n1429) );
  NBUFFX2 U494 ( .INP(n2131), .Z(n1428) );
  NBUFFX2 U495 ( .INP(n2131), .Z(n1427) );
  NBUFFX2 U496 ( .INP(n2131), .Z(n1426) );
  NBUFFX2 U497 ( .INP(n2131), .Z(n1425) );
  NBUFFX2 U498 ( .INP(n2131), .Z(n1424) );
  NBUFFX2 U499 ( .INP(n2131), .Z(n1423) );
  NBUFFX2 U500 ( .INP(n2131), .Z(n1422) );
  NBUFFX2 U501 ( .INP(n2131), .Z(n1421) );
  NBUFFX2 U502 ( .INP(n2131), .Z(n1420) );
  NBUFFX2 U503 ( .INP(n2131), .Z(n1419) );
  NBUFFX2 U504 ( .INP(n2131), .Z(n1418) );
  NBUFFX2 U505 ( .INP(n2131), .Z(n1417) );
  NBUFFX2 U506 ( .INP(n2132), .Z(n1416) );
  NBUFFX2 U507 ( .INP(n2132), .Z(n1415) );
  NBUFFX2 U508 ( .INP(n2132), .Z(n1414) );
  NBUFFX2 U509 ( .INP(n2132), .Z(n1413) );
  NBUFFX2 U510 ( .INP(n2132), .Z(n1412) );
  NBUFFX2 U511 ( .INP(n2132), .Z(n1411) );
  NBUFFX2 U512 ( .INP(n2132), .Z(n1410) );
  NBUFFX2 U513 ( .INP(n2132), .Z(n1407) );
  NBUFFX2 U514 ( .INP(n2132), .Z(n1406) );
  NBUFFX2 U515 ( .INP(n2132), .Z(n1405) );
  NBUFFX2 U516 ( .INP(n2133), .Z(n1404) );
  NBUFFX2 U517 ( .INP(n2133), .Z(n1403) );
  NBUFFX2 U518 ( .INP(n2133), .Z(n1402) );
  NBUFFX2 U519 ( .INP(n2133), .Z(n1401) );
  NBUFFX2 U520 ( .INP(n2133), .Z(n1400) );
  NBUFFX2 U521 ( .INP(n2133), .Z(n1399) );
  NBUFFX2 U522 ( .INP(n2133), .Z(n1398) );
  NBUFFX2 U523 ( .INP(n2133), .Z(n1397) );
  NBUFFX2 U524 ( .INP(n2133), .Z(n1396) );
  NBUFFX2 U525 ( .INP(n2133), .Z(n1395) );
  NBUFFX2 U526 ( .INP(n2133), .Z(n1394) );
  NBUFFX2 U527 ( .INP(n2133), .Z(n1393) );
  NBUFFX2 U528 ( .INP(n2105), .Z(n1736) );
  NBUFFX2 U529 ( .INP(n2105), .Z(n1735) );
  NBUFFX2 U530 ( .INP(n2105), .Z(n1734) );
  NBUFFX2 U531 ( .INP(n2105), .Z(n1733) );
  NBUFFX2 U532 ( .INP(n2105), .Z(n1732) );
  NBUFFX2 U533 ( .INP(n2105), .Z(n1731) );
  NBUFFX2 U534 ( .INP(n2105), .Z(n1730) );
  NBUFFX2 U535 ( .INP(n2105), .Z(n1729) );
  NBUFFX2 U536 ( .INP(n2106), .Z(n1728) );
  NBUFFX2 U537 ( .INP(n2106), .Z(n1727) );
  NBUFFX2 U538 ( .INP(n2106), .Z(n1726) );
  NBUFFX2 U539 ( .INP(n2106), .Z(n1725) );
  NBUFFX2 U540 ( .INP(n2106), .Z(n1724) );
  NBUFFX2 U541 ( .INP(n2106), .Z(n1723) );
  NBUFFX2 U542 ( .INP(n2106), .Z(n1722) );
  NBUFFX2 U543 ( .INP(n2106), .Z(n1721) );
  NBUFFX2 U544 ( .INP(n2106), .Z(n1720) );
  NBUFFX2 U545 ( .INP(n2106), .Z(n1719) );
  NBUFFX2 U546 ( .INP(n2106), .Z(n1718) );
  NBUFFX2 U547 ( .INP(n2106), .Z(n1717) );
  NBUFFX2 U548 ( .INP(n2107), .Z(n1716) );
  NBUFFX2 U549 ( .INP(n2107), .Z(n1715) );
  NBUFFX2 U550 ( .INP(n2107), .Z(n1714) );
  NBUFFX2 U551 ( .INP(n2107), .Z(n1713) );
  NBUFFX2 U552 ( .INP(n2107), .Z(n1712) );
  NBUFFX2 U553 ( .INP(n2107), .Z(n1711) );
  NBUFFX2 U554 ( .INP(n2107), .Z(n1710) );
  NBUFFX2 U555 ( .INP(n2107), .Z(n1709) );
  NBUFFX2 U556 ( .INP(n2107), .Z(n1708) );
  NBUFFX2 U557 ( .INP(n2107), .Z(n1707) );
  NBUFFX2 U558 ( .INP(n2107), .Z(n1706) );
  NBUFFX2 U559 ( .INP(n2107), .Z(n1705) );
  NBUFFX2 U560 ( .INP(n2108), .Z(n1704) );
  NBUFFX2 U561 ( .INP(n2108), .Z(n1703) );
  NBUFFX2 U562 ( .INP(n2108), .Z(n1702) );
  NBUFFX2 U563 ( .INP(n2108), .Z(n1701) );
  NBUFFX2 U564 ( .INP(n2108), .Z(n1700) );
  NBUFFX2 U565 ( .INP(n2108), .Z(n1699) );
  NBUFFX2 U566 ( .INP(n2108), .Z(n1698) );
  NBUFFX2 U567 ( .INP(n2108), .Z(n1697) );
  NBUFFX2 U568 ( .INP(n2108), .Z(n1696) );
  NBUFFX2 U569 ( .INP(n2108), .Z(n1695) );
  NBUFFX2 U570 ( .INP(n2108), .Z(n1694) );
  NBUFFX2 U571 ( .INP(n2108), .Z(n1693) );
  NBUFFX2 U572 ( .INP(n2109), .Z(n1692) );
  NBUFFX2 U573 ( .INP(n2109), .Z(n1691) );
  NBUFFX2 U574 ( .INP(n2109), .Z(n1690) );
  NBUFFX2 U575 ( .INP(n2109), .Z(n1689) );
  NBUFFX2 U576 ( .INP(n2109), .Z(n1688) );
  NBUFFX2 U577 ( .INP(n2109), .Z(n1687) );
  NBUFFX2 U578 ( .INP(n2109), .Z(n1686) );
  NBUFFX2 U579 ( .INP(n2109), .Z(n1685) );
  NBUFFX2 U580 ( .INP(n2109), .Z(n1684) );
  NBUFFX2 U581 ( .INP(n2109), .Z(n1683) );
  NBUFFX2 U582 ( .INP(n2109), .Z(n1682) );
  NBUFFX2 U583 ( .INP(n2109), .Z(n1681) );
  NBUFFX2 U584 ( .INP(n2110), .Z(n1680) );
  NBUFFX2 U585 ( .INP(n2110), .Z(n1679) );
  NBUFFX2 U586 ( .INP(n2110), .Z(n1678) );
  NBUFFX2 U587 ( .INP(n2110), .Z(n1677) );
  NBUFFX2 U588 ( .INP(n2110), .Z(n1676) );
  NBUFFX2 U589 ( .INP(n2110), .Z(n1675) );
  NBUFFX2 U590 ( .INP(n2110), .Z(n1674) );
  NBUFFX2 U591 ( .INP(n2110), .Z(n1673) );
  NBUFFX2 U592 ( .INP(n2110), .Z(n1672) );
  NBUFFX2 U593 ( .INP(n2110), .Z(n1671) );
  NBUFFX2 U594 ( .INP(n2110), .Z(n1670) );
  NBUFFX2 U595 ( .INP(n2110), .Z(n1669) );
  NBUFFX2 U596 ( .INP(n2111), .Z(n1668) );
  NBUFFX2 U597 ( .INP(n2111), .Z(n1667) );
  NBUFFX2 U598 ( .INP(n2111), .Z(n1666) );
  NBUFFX2 U599 ( .INP(n2111), .Z(n1665) );
  NBUFFX2 U600 ( .INP(n2111), .Z(n1664) );
  NBUFFX2 U601 ( .INP(n2111), .Z(n1663) );
  NBUFFX2 U602 ( .INP(n2111), .Z(n1662) );
  NBUFFX2 U603 ( .INP(n2111), .Z(n1661) );
  NBUFFX2 U604 ( .INP(n2111), .Z(n1660) );
  NBUFFX2 U605 ( .INP(n2111), .Z(n1659) );
  NBUFFX2 U606 ( .INP(n2111), .Z(n1658) );
  NBUFFX2 U607 ( .INP(n2111), .Z(n1657) );
  NBUFFX2 U608 ( .INP(n2112), .Z(n1656) );
  NBUFFX2 U609 ( .INP(n2112), .Z(n1655) );
  NBUFFX2 U610 ( .INP(n2112), .Z(n1654) );
  NBUFFX2 U611 ( .INP(n2112), .Z(n1653) );
  NBUFFX2 U612 ( .INP(n2112), .Z(n1652) );
  NBUFFX2 U613 ( .INP(n2112), .Z(n1651) );
  NBUFFX2 U614 ( .INP(n2112), .Z(n1650) );
  NBUFFX2 U615 ( .INP(n2112), .Z(n1649) );
  NBUFFX2 U616 ( .INP(n2112), .Z(n1648) );
  NBUFFX2 U617 ( .INP(n2112), .Z(n1647) );
  NBUFFX2 U618 ( .INP(n2112), .Z(n1646) );
  NBUFFX2 U619 ( .INP(n2112), .Z(n1645) );
  NBUFFX2 U620 ( .INP(n2113), .Z(n1644) );
  NBUFFX2 U621 ( .INP(n2113), .Z(n1643) );
  NBUFFX2 U622 ( .INP(n2113), .Z(n1642) );
  NBUFFX2 U623 ( .INP(n2113), .Z(n1641) );
  NBUFFX2 U624 ( .INP(n2113), .Z(n1640) );
  NBUFFX2 U625 ( .INP(n2113), .Z(n1639) );
  NBUFFX2 U626 ( .INP(n2113), .Z(n1638) );
  NBUFFX2 U627 ( .INP(n2113), .Z(n1637) );
  NBUFFX2 U628 ( .INP(n2113), .Z(n1636) );
  NBUFFX2 U629 ( .INP(n2113), .Z(n1635) );
  NBUFFX2 U630 ( .INP(n2113), .Z(n1634) );
  NBUFFX2 U631 ( .INP(n2113), .Z(n1633) );
  NBUFFX2 U632 ( .INP(n2114), .Z(n1632) );
  NBUFFX2 U633 ( .INP(n2114), .Z(n1631) );
  NBUFFX2 U634 ( .INP(n2114), .Z(n1630) );
  NBUFFX2 U635 ( .INP(n2114), .Z(n1629) );
  NBUFFX2 U636 ( .INP(n2114), .Z(n1628) );
  NBUFFX2 U637 ( .INP(n2114), .Z(n1627) );
  NBUFFX2 U638 ( .INP(n2114), .Z(n1626) );
  NBUFFX2 U639 ( .INP(n2114), .Z(n1625) );
  NBUFFX2 U640 ( .INP(n2114), .Z(n1624) );
  NBUFFX2 U641 ( .INP(n2114), .Z(n1623) );
  NBUFFX2 U642 ( .INP(n2114), .Z(n1622) );
  NBUFFX2 U643 ( .INP(n2114), .Z(n1621) );
  NBUFFX2 U644 ( .INP(n2115), .Z(n1620) );
  NBUFFX2 U645 ( .INP(n2115), .Z(n1619) );
  NBUFFX2 U646 ( .INP(n2115), .Z(n1618) );
  NBUFFX2 U647 ( .INP(n2115), .Z(n1617) );
  NBUFFX2 U648 ( .INP(n2115), .Z(n1616) );
  NBUFFX2 U649 ( .INP(n2115), .Z(n1615) );
  NBUFFX2 U650 ( .INP(n2115), .Z(n1614) );
  NBUFFX2 U651 ( .INP(n2115), .Z(n1613) );
  NBUFFX2 U652 ( .INP(n2115), .Z(n1612) );
  NBUFFX2 U653 ( .INP(n2115), .Z(n1611) );
  NBUFFX2 U654 ( .INP(n2115), .Z(n1610) );
  NBUFFX2 U655 ( .INP(n2115), .Z(n1609) );
  NBUFFX2 U656 ( .INP(n2116), .Z(n1608) );
  NBUFFX2 U657 ( .INP(n2116), .Z(n1607) );
  NBUFFX2 U658 ( .INP(n2116), .Z(n1606) );
  NBUFFX2 U659 ( .INP(n2116), .Z(n1605) );
  NBUFFX2 U660 ( .INP(n2116), .Z(n1604) );
  NBUFFX2 U661 ( .INP(n2116), .Z(n1603) );
  NBUFFX2 U662 ( .INP(n2116), .Z(n1602) );
  NBUFFX2 U663 ( .INP(n2116), .Z(n1601) );
  NBUFFX2 U664 ( .INP(n2116), .Z(n1600) );
  NBUFFX2 U665 ( .INP(n2116), .Z(n1599) );
  NBUFFX2 U666 ( .INP(n2116), .Z(n1598) );
  NBUFFX2 U667 ( .INP(n2116), .Z(n1597) );
  NBUFFX2 U668 ( .INP(n2117), .Z(n1596) );
  NBUFFX2 U669 ( .INP(n2117), .Z(n1595) );
  NBUFFX2 U670 ( .INP(n2117), .Z(n1594) );
  NBUFFX2 U671 ( .INP(n2117), .Z(n1593) );
  NBUFFX2 U672 ( .INP(n2117), .Z(n1592) );
  NBUFFX2 U673 ( .INP(n2117), .Z(n1591) );
  NBUFFX2 U674 ( .INP(n2117), .Z(n1590) );
  NBUFFX2 U675 ( .INP(n2117), .Z(n1589) );
  NBUFFX2 U676 ( .INP(n2117), .Z(n1588) );
  NBUFFX2 U677 ( .INP(n2117), .Z(n1587) );
  NBUFFX2 U678 ( .INP(n2117), .Z(n1586) );
  NBUFFX2 U679 ( .INP(n2117), .Z(n1585) );
  NBUFFX2 U680 ( .INP(n2118), .Z(n1584) );
  NBUFFX2 U681 ( .INP(n2118), .Z(n1583) );
  NBUFFX2 U682 ( .INP(n2118), .Z(n1582) );
  NBUFFX2 U683 ( .INP(n2118), .Z(n1581) );
  NBUFFX2 U684 ( .INP(n2105), .Z(n1737) );
  NBUFFX2 U685 ( .INP(n2077), .Z(n2076) );
  DELLN1X2 U686 ( .INP(n2206), .Z(n141) );
  NBUFFX2 U687 ( .INP(n2206), .Z(n143) );
  NBUFFX2 U688 ( .INP(n2206), .Z(n144) );
  NBUFFX2 U689 ( .INP(n2206), .Z(n145) );
  NBUFFX2 U690 ( .INP(n2206), .Z(n147) );
  NBUFFX2 U691 ( .INP(n2206), .Z(n148) );
  NBUFFX2 U692 ( .INP(n2206), .Z(n149) );
  NBUFFX2 U693 ( .INP(n2206), .Z(n151) );
  NBUFFX2 U694 ( .INP(n2206), .Z(n152) );
  NBUFFX2 U695 ( .INP(n2206), .Z(n153) );
  NBUFFX2 U696 ( .INP(n2206), .Z(n155) );
  NBUFFX2 U697 ( .INP(n2206), .Z(n156) );
  NBUFFX2 U698 ( .INP(n2206), .Z(n157) );
  NBUFFX2 U699 ( .INP(n2206), .Z(n159) );
  NBUFFX2 U700 ( .INP(n2206), .Z(n160) );
  NBUFFX2 U701 ( .INP(n2206), .Z(n161) );
  NBUFFX2 U702 ( .INP(n2206), .Z(n163) );
  NBUFFX2 U703 ( .INP(n2206), .Z(n164) );
  NBUFFX2 U704 ( .INP(n2206), .Z(n165) );
  NBUFFX2 U705 ( .INP(n2206), .Z(n167) );
  NBUFFX2 U706 ( .INP(n2206), .Z(n168) );
  NBUFFX2 U707 ( .INP(n2206), .Z(n169) );
  NBUFFX2 U708 ( .INP(n2206), .Z(n171) );
  NBUFFX2 U709 ( .INP(n2206), .Z(n172) );
  NBUFFX2 U710 ( .INP(n2151), .Z(n2080) );
  NBUFFX2 U711 ( .INP(n2151), .Z(n2081) );
  NBUFFX2 U712 ( .INP(n2151), .Z(n2082) );
  NBUFFX2 U713 ( .INP(n2150), .Z(n2083) );
  NBUFFX2 U714 ( .INP(n2150), .Z(n2084) );
  NBUFFX2 U715 ( .INP(n2150), .Z(n2085) );
  NBUFFX2 U716 ( .INP(n2149), .Z(n2086) );
  NBUFFX2 U717 ( .INP(n2149), .Z(n2087) );
  NBUFFX2 U718 ( .INP(n2149), .Z(n2088) );
  NBUFFX2 U719 ( .INP(n2148), .Z(n2089) );
  NBUFFX2 U720 ( .INP(n2148), .Z(n2090) );
  NBUFFX2 U721 ( .INP(n2148), .Z(n2091) );
  NBUFFX2 U722 ( .INP(n2147), .Z(n2092) );
  NBUFFX2 U723 ( .INP(n2147), .Z(n2093) );
  NBUFFX2 U724 ( .INP(n2147), .Z(n2094) );
  NBUFFX2 U725 ( .INP(n2146), .Z(n2095) );
  NBUFFX2 U726 ( .INP(n2146), .Z(n2096) );
  NBUFFX2 U727 ( .INP(n2146), .Z(n2097) );
  NBUFFX2 U728 ( .INP(n2145), .Z(n2098) );
  NBUFFX2 U729 ( .INP(n2145), .Z(n2099) );
  NBUFFX2 U730 ( .INP(n2145), .Z(n2100) );
  NBUFFX2 U731 ( .INP(n2144), .Z(n2101) );
  NBUFFX2 U732 ( .INP(n2144), .Z(n2102) );
  NBUFFX2 U733 ( .INP(n2144), .Z(n2103) );
  NBUFFX2 U734 ( .INP(n2143), .Z(n2104) );
  NBUFFX2 U735 ( .INP(n2152), .Z(n2078) );
  NBUFFX2 U736 ( .INP(n2152), .Z(n2079) );
  NBUFFX2 U737 ( .INP(n2152), .Z(n2077) );
  NBUFFX2 U738 ( .INP(n2138), .Z(n2119) );
  NBUFFX2 U739 ( .INP(n2138), .Z(n2120) );
  NBUFFX2 U740 ( .INP(n2138), .Z(n2121) );
  NBUFFX2 U741 ( .INP(n2137), .Z(n2122) );
  NBUFFX2 U742 ( .INP(n2137), .Z(n2123) );
  NBUFFX2 U743 ( .INP(n2137), .Z(n2124) );
  NBUFFX2 U744 ( .INP(n2136), .Z(n2125) );
  NBUFFX2 U745 ( .INP(n2136), .Z(n2126) );
  NBUFFX2 U746 ( .INP(n2136), .Z(n2127) );
  NBUFFX2 U747 ( .INP(n2135), .Z(n2128) );
  NBUFFX2 U748 ( .INP(n2135), .Z(n2129) );
  NBUFFX2 U749 ( .INP(n2135), .Z(n2130) );
  NBUFFX2 U750 ( .INP(n2134), .Z(n2131) );
  NBUFFX2 U751 ( .INP(n2134), .Z(n2132) );
  NBUFFX2 U752 ( .INP(n2134), .Z(n2133) );
  NBUFFX2 U753 ( .INP(n2143), .Z(n2106) );
  NBUFFX2 U754 ( .INP(n2142), .Z(n2107) );
  NBUFFX2 U755 ( .INP(n2142), .Z(n2108) );
  NBUFFX2 U756 ( .INP(n2142), .Z(n2109) );
  NBUFFX2 U757 ( .INP(n2141), .Z(n2110) );
  NBUFFX2 U758 ( .INP(n2141), .Z(n2111) );
  NBUFFX2 U759 ( .INP(n2141), .Z(n2112) );
  NBUFFX2 U760 ( .INP(n2140), .Z(n2113) );
  NBUFFX2 U761 ( .INP(n2140), .Z(n2114) );
  NBUFFX2 U762 ( .INP(n2140), .Z(n2115) );
  NBUFFX2 U763 ( .INP(n2139), .Z(n2116) );
  NBUFFX2 U764 ( .INP(n2139), .Z(n2117) );
  NBUFFX2 U765 ( .INP(n2139), .Z(n2118) );
  NBUFFX2 U766 ( .INP(n2143), .Z(n2105) );
  DELLN1X2 U767 ( .INP(n2215), .Z(n442) );
  DELLN1X2 U768 ( .INP(n2205), .Z(n98) );
  DELLN1X2 U769 ( .INP(n2220), .Z(n614) );
  NBUFFX2 U770 ( .INP(n2215), .Z(n444) );
  NBUFFX2 U771 ( .INP(n2205), .Z(n100) );
  NBUFFX2 U772 ( .INP(n2220), .Z(n616) );
  NBUFFX2 U773 ( .INP(n2215), .Z(n445) );
  NBUFFX2 U774 ( .INP(n2205), .Z(n101) );
  NBUFFX2 U775 ( .INP(n2220), .Z(n617) );
  NBUFFX2 U776 ( .INP(n2215), .Z(n446) );
  NBUFFX2 U777 ( .INP(n2205), .Z(n102) );
  NBUFFX2 U778 ( .INP(n2220), .Z(n618) );
  NBUFFX2 U779 ( .INP(n2215), .Z(n448) );
  NBUFFX2 U780 ( .INP(n2205), .Z(n104) );
  NBUFFX2 U781 ( .INP(n2220), .Z(n620) );
  NBUFFX2 U782 ( .INP(n2215), .Z(n449) );
  NBUFFX2 U783 ( .INP(n2205), .Z(n105) );
  NBUFFX2 U784 ( .INP(n2220), .Z(n621) );
  DELLN1X2 U785 ( .INP(n2210), .Z(n278) );
  NBUFFX2 U786 ( .INP(n2215), .Z(n450) );
  NBUFFX2 U787 ( .INP(n2205), .Z(n106) );
  NBUFFX2 U788 ( .INP(n2220), .Z(n622) );
  NBUFFX2 U789 ( .INP(n2210), .Z(n279) );
  NBUFFX2 U790 ( .INP(n2210), .Z(n280) );
  NBUFFX2 U791 ( .INP(n2215), .Z(n452) );
  NBUFFX2 U792 ( .INP(n2205), .Z(n108) );
  NBUFFX2 U793 ( .INP(n2220), .Z(n624) );
  NBUFFX2 U794 ( .INP(n2210), .Z(n281) );
  NBUFFX2 U795 ( .INP(n2215), .Z(n453) );
  NBUFFX2 U796 ( .INP(n2205), .Z(n109) );
  NBUFFX2 U797 ( .INP(n2220), .Z(n625) );
  NBUFFX2 U798 ( .INP(n2210), .Z(n282) );
  NBUFFX2 U799 ( .INP(n2215), .Z(n454) );
  NBUFFX2 U800 ( .INP(n2205), .Z(n110) );
  NBUFFX2 U801 ( .INP(n2220), .Z(n626) );
  NBUFFX2 U802 ( .INP(n2210), .Z(n283) );
  NBUFFX2 U803 ( .INP(n2210), .Z(n284) );
  NBUFFX2 U804 ( .INP(n2215), .Z(n456) );
  NBUFFX2 U805 ( .INP(n2205), .Z(n112) );
  NBUFFX2 U806 ( .INP(n2220), .Z(n628) );
  NBUFFX2 U807 ( .INP(n2210), .Z(n285) );
  NBUFFX2 U808 ( .INP(n2215), .Z(n457) );
  NBUFFX2 U809 ( .INP(n2205), .Z(n113) );
  NBUFFX2 U810 ( .INP(n2220), .Z(n629) );
  NBUFFX2 U811 ( .INP(n2210), .Z(n286) );
  NBUFFX2 U812 ( .INP(n2215), .Z(n458) );
  NBUFFX2 U813 ( .INP(n2205), .Z(n114) );
  NBUFFX2 U814 ( .INP(n2220), .Z(n630) );
  NBUFFX2 U815 ( .INP(n2210), .Z(n287) );
  NBUFFX2 U816 ( .INP(n2210), .Z(n288) );
  NBUFFX2 U817 ( .INP(n2215), .Z(n460) );
  NBUFFX2 U818 ( .INP(n2205), .Z(n116) );
  NBUFFX2 U819 ( .INP(n2220), .Z(n632) );
  NBUFFX2 U820 ( .INP(n2210), .Z(n289) );
  NBUFFX2 U821 ( .INP(n2215), .Z(n461) );
  NBUFFX2 U822 ( .INP(n2205), .Z(n117) );
  NBUFFX2 U823 ( .INP(n2220), .Z(n633) );
  NBUFFX2 U824 ( .INP(n2210), .Z(n290) );
  NBUFFX2 U825 ( .INP(n2215), .Z(n462) );
  NBUFFX2 U826 ( .INP(n2205), .Z(n118) );
  NBUFFX2 U827 ( .INP(n2220), .Z(n634) );
  NBUFFX2 U828 ( .INP(n2210), .Z(n291) );
  NBUFFX2 U829 ( .INP(n2210), .Z(n292) );
  NBUFFX2 U830 ( .INP(n2215), .Z(n464) );
  NBUFFX2 U831 ( .INP(n2205), .Z(n120) );
  NBUFFX2 U832 ( .INP(n2220), .Z(n636) );
  NBUFFX2 U833 ( .INP(n2210), .Z(n293) );
  NBUFFX2 U834 ( .INP(n2215), .Z(n465) );
  NBUFFX2 U835 ( .INP(n2205), .Z(n121) );
  NBUFFX2 U836 ( .INP(n2220), .Z(n637) );
  NBUFFX2 U837 ( .INP(n2210), .Z(n294) );
  NBUFFX2 U838 ( .INP(n2215), .Z(n466) );
  NBUFFX2 U839 ( .INP(n2205), .Z(n122) );
  NBUFFX2 U840 ( .INP(n2220), .Z(n638) );
  NBUFFX2 U841 ( .INP(n2210), .Z(n295) );
  NBUFFX2 U842 ( .INP(n2210), .Z(n296) );
  NBUFFX2 U843 ( .INP(n2215), .Z(n468) );
  NBUFFX2 U844 ( .INP(n2205), .Z(n124) );
  NBUFFX2 U845 ( .INP(n2220), .Z(n640) );
  NBUFFX2 U846 ( .INP(n2210), .Z(n297) );
  NBUFFX2 U847 ( .INP(n2215), .Z(n469) );
  NBUFFX2 U848 ( .INP(n2205), .Z(n125) );
  NBUFFX2 U849 ( .INP(n2220), .Z(n641) );
  NBUFFX2 U850 ( .INP(n2210), .Z(n298) );
  NBUFFX2 U851 ( .INP(n2215), .Z(n470) );
  NBUFFX2 U852 ( .INP(n2205), .Z(n126) );
  NBUFFX2 U853 ( .INP(n2220), .Z(n642) );
  NBUFFX2 U854 ( .INP(n2210), .Z(n299) );
  NBUFFX2 U855 ( .INP(n2210), .Z(n300) );
  NBUFFX2 U856 ( .INP(n2215), .Z(n472) );
  NBUFFX2 U857 ( .INP(n2205), .Z(n128) );
  NBUFFX2 U858 ( .INP(n2220), .Z(n644) );
  DELLN1X2 U859 ( .INP(n2216), .Z(n485) );
  DELLN1X2 U860 ( .INP(n2221), .Z(n657) );
  NBUFFX2 U861 ( .INP(n2216), .Z(n487) );
  NBUFFX2 U862 ( .INP(n2221), .Z(n659) );
  NBUFFX2 U863 ( .INP(n2216), .Z(n488) );
  NBUFFX2 U864 ( .INP(n2221), .Z(n660) );
  NBUFFX2 U865 ( .INP(n2216), .Z(n489) );
  NBUFFX2 U866 ( .INP(n2221), .Z(n661) );
  NBUFFX2 U867 ( .INP(n2216), .Z(n491) );
  NBUFFX2 U868 ( .INP(n2221), .Z(n663) );
  NBUFFX2 U869 ( .INP(n2216), .Z(n492) );
  NBUFFX2 U870 ( .INP(n2221), .Z(n664) );
  DELLN1X2 U871 ( .INP(n2211), .Z(n321) );
  NBUFFX2 U872 ( .INP(n2216), .Z(n493) );
  NBUFFX2 U873 ( .INP(n2221), .Z(n665) );
  NBUFFX2 U874 ( .INP(n2211), .Z(n322) );
  NBUFFX2 U875 ( .INP(n2211), .Z(n323) );
  NBUFFX2 U876 ( .INP(n2216), .Z(n495) );
  NBUFFX2 U877 ( .INP(n2221), .Z(n667) );
  NBUFFX2 U878 ( .INP(n2211), .Z(n324) );
  NBUFFX2 U879 ( .INP(n2216), .Z(n496) );
  NBUFFX2 U880 ( .INP(n2221), .Z(n668) );
  NBUFFX2 U881 ( .INP(n2211), .Z(n325) );
  NBUFFX2 U882 ( .INP(n2216), .Z(n497) );
  NBUFFX2 U883 ( .INP(n2221), .Z(n669) );
  NBUFFX2 U884 ( .INP(n2211), .Z(n326) );
  NBUFFX2 U885 ( .INP(n2211), .Z(n327) );
  NBUFFX2 U886 ( .INP(n2216), .Z(n499) );
  NBUFFX2 U887 ( .INP(n2221), .Z(n671) );
  NBUFFX2 U888 ( .INP(n2211), .Z(n328) );
  NBUFFX2 U889 ( .INP(n2216), .Z(n500) );
  NBUFFX2 U890 ( .INP(n2221), .Z(n672) );
  NBUFFX2 U891 ( .INP(n2211), .Z(n329) );
  NBUFFX2 U892 ( .INP(n2216), .Z(n501) );
  NBUFFX2 U893 ( .INP(n2221), .Z(n673) );
  NBUFFX2 U894 ( .INP(n2211), .Z(n330) );
  NBUFFX2 U895 ( .INP(n2211), .Z(n331) );
  NBUFFX2 U896 ( .INP(n2216), .Z(n503) );
  NBUFFX2 U897 ( .INP(n2221), .Z(n675) );
  NBUFFX2 U898 ( .INP(n2211), .Z(n332) );
  NBUFFX2 U899 ( .INP(n2216), .Z(n504) );
  NBUFFX2 U900 ( .INP(n2221), .Z(n676) );
  NBUFFX2 U901 ( .INP(n2211), .Z(n333) );
  NBUFFX2 U902 ( .INP(n2216), .Z(n505) );
  NBUFFX2 U903 ( .INP(n2221), .Z(n677) );
  NBUFFX2 U904 ( .INP(n2211), .Z(n334) );
  NBUFFX2 U905 ( .INP(n2211), .Z(n335) );
  NBUFFX2 U906 ( .INP(n2216), .Z(n507) );
  NBUFFX2 U907 ( .INP(n2221), .Z(n679) );
  NBUFFX2 U908 ( .INP(n2211), .Z(n336) );
  NBUFFX2 U909 ( .INP(n2216), .Z(n508) );
  NBUFFX2 U910 ( .INP(n2221), .Z(n680) );
  NBUFFX2 U911 ( .INP(n2211), .Z(n337) );
  NBUFFX2 U912 ( .INP(n2216), .Z(n509) );
  NBUFFX2 U913 ( .INP(n2221), .Z(n681) );
  NBUFFX2 U914 ( .INP(n2211), .Z(n338) );
  NBUFFX2 U915 ( .INP(n2211), .Z(n339) );
  NBUFFX2 U916 ( .INP(n2216), .Z(n511) );
  NBUFFX2 U917 ( .INP(n2221), .Z(n683) );
  NBUFFX2 U918 ( .INP(n2211), .Z(n340) );
  NBUFFX2 U919 ( .INP(n2216), .Z(n512) );
  NBUFFX2 U920 ( .INP(n2221), .Z(n684) );
  NBUFFX2 U921 ( .INP(n2211), .Z(n341) );
  NBUFFX2 U922 ( .INP(n2216), .Z(n513) );
  NBUFFX2 U923 ( .INP(n2221), .Z(n685) );
  NBUFFX2 U924 ( .INP(n2211), .Z(n342) );
  NBUFFX2 U925 ( .INP(n2211), .Z(n343) );
  NBUFFX2 U926 ( .INP(n2216), .Z(n515) );
  NBUFFX2 U927 ( .INP(n2221), .Z(n687) );
  DELLN1X2 U928 ( .INP(n2208), .Z(n235) );
  NBUFFX2 U929 ( .INP(n2208), .Z(n236) );
  NBUFFX2 U930 ( .INP(n2208), .Z(n237) );
  NBUFFX2 U931 ( .INP(n2208), .Z(n238) );
  NBUFFX2 U932 ( .INP(n2208), .Z(n239) );
  NBUFFX2 U933 ( .INP(n2208), .Z(n240) );
  NBUFFX2 U934 ( .INP(n2208), .Z(n241) );
  NBUFFX2 U935 ( .INP(n2208), .Z(n242) );
  NBUFFX2 U936 ( .INP(n2208), .Z(n243) );
  NBUFFX2 U937 ( .INP(n2208), .Z(n244) );
  NBUFFX2 U938 ( .INP(n2208), .Z(n245) );
  NBUFFX2 U939 ( .INP(n2208), .Z(n246) );
  NBUFFX2 U940 ( .INP(n2208), .Z(n247) );
  NBUFFX2 U941 ( .INP(n2208), .Z(n248) );
  NBUFFX2 U942 ( .INP(n2208), .Z(n249) );
  NBUFFX2 U943 ( .INP(n2208), .Z(n250) );
  NBUFFX2 U944 ( .INP(n2208), .Z(n251) );
  NBUFFX2 U945 ( .INP(n2208), .Z(n252) );
  NBUFFX2 U946 ( .INP(n2208), .Z(n253) );
  NBUFFX2 U947 ( .INP(n2208), .Z(n254) );
  NBUFFX2 U948 ( .INP(n2208), .Z(n255) );
  NBUFFX2 U949 ( .INP(n2208), .Z(n256) );
  NBUFFX2 U950 ( .INP(n2208), .Z(n257) );
  DELLN1X2 U951 ( .INP(n2213), .Z(n407) );
  DELLN1X2 U952 ( .INP(n2194), .Z(n63) );
  DELLN1X2 U953 ( .INP(n2218), .Z(n579) );
  NBUFFX2 U954 ( .INP(n2213), .Z(n408) );
  NBUFFX2 U955 ( .INP(n2194), .Z(n64) );
  NBUFFX2 U956 ( .INP(n2218), .Z(n580) );
  NBUFFX2 U957 ( .INP(n2213), .Z(n409) );
  NBUFFX2 U958 ( .INP(n2194), .Z(n65) );
  NBUFFX2 U959 ( .INP(n2218), .Z(n581) );
  NBUFFX2 U960 ( .INP(n2213), .Z(n410) );
  NBUFFX2 U961 ( .INP(n2194), .Z(n66) );
  NBUFFX2 U962 ( .INP(n2218), .Z(n582) );
  NBUFFX2 U963 ( .INP(n2213), .Z(n411) );
  NBUFFX2 U964 ( .INP(n2194), .Z(n67) );
  NBUFFX2 U965 ( .INP(n2218), .Z(n583) );
  NBUFFX2 U966 ( .INP(n2213), .Z(n412) );
  NBUFFX2 U967 ( .INP(n2194), .Z(n68) );
  NBUFFX2 U968 ( .INP(n2218), .Z(n584) );
  NBUFFX2 U969 ( .INP(n2213), .Z(n413) );
  NBUFFX2 U970 ( .INP(n2194), .Z(n69) );
  NBUFFX2 U971 ( .INP(n2218), .Z(n585) );
  NBUFFX2 U972 ( .INP(n2213), .Z(n414) );
  NBUFFX2 U973 ( .INP(n2194), .Z(n70) );
  NBUFFX2 U974 ( .INP(n2218), .Z(n586) );
  NBUFFX2 U975 ( .INP(n2213), .Z(n415) );
  NBUFFX2 U976 ( .INP(n2194), .Z(n71) );
  NBUFFX2 U977 ( .INP(n2218), .Z(n587) );
  NBUFFX2 U978 ( .INP(n2213), .Z(n416) );
  NBUFFX2 U979 ( .INP(n2194), .Z(n72) );
  NBUFFX2 U980 ( .INP(n2218), .Z(n588) );
  NBUFFX2 U981 ( .INP(n2213), .Z(n417) );
  NBUFFX2 U982 ( .INP(n2194), .Z(n73) );
  NBUFFX2 U983 ( .INP(n2218), .Z(n589) );
  NBUFFX2 U984 ( .INP(n2213), .Z(n418) );
  NBUFFX2 U985 ( .INP(n2194), .Z(n74) );
  NBUFFX2 U986 ( .INP(n2218), .Z(n590) );
  NBUFFX2 U987 ( .INP(n2213), .Z(n419) );
  NBUFFX2 U988 ( .INP(n2194), .Z(n75) );
  NBUFFX2 U989 ( .INP(n2218), .Z(n591) );
  NBUFFX2 U990 ( .INP(n2213), .Z(n420) );
  NBUFFX2 U991 ( .INP(n2194), .Z(n76) );
  NBUFFX2 U992 ( .INP(n2218), .Z(n592) );
  NBUFFX2 U993 ( .INP(n2213), .Z(n421) );
  NBUFFX2 U994 ( .INP(n2194), .Z(n77) );
  NBUFFX2 U995 ( .INP(n2218), .Z(n593) );
  NBUFFX2 U996 ( .INP(n2213), .Z(n422) );
  NBUFFX2 U997 ( .INP(n2194), .Z(n78) );
  NBUFFX2 U998 ( .INP(n2218), .Z(n594) );
  NBUFFX2 U999 ( .INP(n2213), .Z(n423) );
  NBUFFX2 U1000 ( .INP(n2194), .Z(n79) );
  NBUFFX2 U1001 ( .INP(n2218), .Z(n595) );
  NBUFFX2 U1002 ( .INP(n2213), .Z(n424) );
  NBUFFX2 U1003 ( .INP(n2194), .Z(n80) );
  NBUFFX2 U1004 ( .INP(n2218), .Z(n596) );
  NBUFFX2 U1005 ( .INP(n2213), .Z(n425) );
  NBUFFX2 U1006 ( .INP(n2194), .Z(n81) );
  NBUFFX2 U1007 ( .INP(n2218), .Z(n597) );
  NBUFFX2 U1008 ( .INP(n2213), .Z(n426) );
  NBUFFX2 U1009 ( .INP(n2194), .Z(n82) );
  NBUFFX2 U1010 ( .INP(n2218), .Z(n598) );
  NBUFFX2 U1011 ( .INP(n2213), .Z(n427) );
  NBUFFX2 U1012 ( .INP(n2194), .Z(n83) );
  NBUFFX2 U1013 ( .INP(n2218), .Z(n599) );
  NBUFFX2 U1014 ( .INP(n2213), .Z(n428) );
  NBUFFX2 U1015 ( .INP(n2194), .Z(n84) );
  NBUFFX2 U1016 ( .INP(n2218), .Z(n600) );
  NBUFFX2 U1017 ( .INP(n2213), .Z(n429) );
  NBUFFX2 U1018 ( .INP(n2194), .Z(n85) );
  NBUFFX2 U1019 ( .INP(n2218), .Z(n601) );
  DELLN1X2 U1020 ( .INP(n2207), .Z(n192) );
  NBUFFX2 U1021 ( .INP(n2207), .Z(n193) );
  NBUFFX2 U1022 ( .INP(n2207), .Z(n194) );
  NBUFFX2 U1023 ( .INP(n2207), .Z(n195) );
  NBUFFX2 U1024 ( .INP(n2207), .Z(n196) );
  NBUFFX2 U1025 ( .INP(n2207), .Z(n197) );
  NBUFFX2 U1026 ( .INP(n2207), .Z(n198) );
  NBUFFX2 U1027 ( .INP(n2207), .Z(n199) );
  NBUFFX2 U1028 ( .INP(n2207), .Z(n200) );
  NBUFFX2 U1029 ( .INP(n2207), .Z(n201) );
  NBUFFX2 U1030 ( .INP(n2207), .Z(n202) );
  NBUFFX2 U1031 ( .INP(n2207), .Z(n203) );
  NBUFFX2 U1032 ( .INP(n2207), .Z(n204) );
  NBUFFX2 U1033 ( .INP(n2207), .Z(n205) );
  NBUFFX2 U1034 ( .INP(n2207), .Z(n206) );
  NBUFFX2 U1035 ( .INP(n2207), .Z(n207) );
  NBUFFX2 U1036 ( .INP(n2207), .Z(n208) );
  NBUFFX2 U1037 ( .INP(n2207), .Z(n209) );
  NBUFFX2 U1038 ( .INP(n2207), .Z(n210) );
  NBUFFX2 U1039 ( .INP(n2207), .Z(n211) );
  NBUFFX2 U1040 ( .INP(n2207), .Z(n212) );
  NBUFFX2 U1041 ( .INP(n2207), .Z(n213) );
  NBUFFX2 U1042 ( .INP(n2207), .Z(n214) );
  DELLN1X2 U1043 ( .INP(n2212), .Z(n364) );
  DELLN1X2 U1044 ( .INP(n2170), .Z(n20) );
  DELLN1X2 U1045 ( .INP(n2217), .Z(n536) );
  NBUFFX2 U1046 ( .INP(n2212), .Z(n365) );
  NBUFFX2 U1047 ( .INP(n2170), .Z(n21) );
  NBUFFX2 U1048 ( .INP(n2217), .Z(n537) );
  NBUFFX2 U1049 ( .INP(n2212), .Z(n366) );
  NBUFFX2 U1050 ( .INP(n2170), .Z(n22) );
  NBUFFX2 U1051 ( .INP(n2217), .Z(n538) );
  NBUFFX2 U1052 ( .INP(n2212), .Z(n367) );
  NBUFFX2 U1053 ( .INP(n2170), .Z(n23) );
  NBUFFX2 U1054 ( .INP(n2217), .Z(n539) );
  NBUFFX2 U1055 ( .INP(n2212), .Z(n368) );
  NBUFFX2 U1056 ( .INP(n2170), .Z(n24) );
  NBUFFX2 U1057 ( .INP(n2217), .Z(n540) );
  NBUFFX2 U1058 ( .INP(n2212), .Z(n369) );
  NBUFFX2 U1059 ( .INP(n2170), .Z(n25) );
  NBUFFX2 U1060 ( .INP(n2217), .Z(n541) );
  NBUFFX2 U1061 ( .INP(n2212), .Z(n370) );
  NBUFFX2 U1062 ( .INP(n2170), .Z(n26) );
  NBUFFX2 U1063 ( .INP(n2217), .Z(n542) );
  NBUFFX2 U1064 ( .INP(n2212), .Z(n371) );
  NBUFFX2 U1065 ( .INP(n2170), .Z(n27) );
  NBUFFX2 U1066 ( .INP(n2217), .Z(n543) );
  NBUFFX2 U1067 ( .INP(n2212), .Z(n372) );
  NBUFFX2 U1068 ( .INP(n2170), .Z(n28) );
  NBUFFX2 U1069 ( .INP(n2217), .Z(n544) );
  NBUFFX2 U1070 ( .INP(n2212), .Z(n373) );
  NBUFFX2 U1071 ( .INP(n2170), .Z(n29) );
  NBUFFX2 U1072 ( .INP(n2217), .Z(n545) );
  NBUFFX2 U1073 ( .INP(n2212), .Z(n374) );
  NBUFFX2 U1074 ( .INP(n2170), .Z(n30) );
  NBUFFX2 U1075 ( .INP(n2217), .Z(n546) );
  NBUFFX2 U1076 ( .INP(n2212), .Z(n375) );
  NBUFFX2 U1077 ( .INP(n2170), .Z(n31) );
  NBUFFX2 U1078 ( .INP(n2217), .Z(n547) );
  NBUFFX2 U1079 ( .INP(n2212), .Z(n376) );
  NBUFFX2 U1080 ( .INP(n2170), .Z(n32) );
  NBUFFX2 U1081 ( .INP(n2217), .Z(n548) );
  NBUFFX2 U1082 ( .INP(n2212), .Z(n377) );
  NBUFFX2 U1083 ( .INP(n2170), .Z(n33) );
  NBUFFX2 U1084 ( .INP(n2217), .Z(n549) );
  NBUFFX2 U1085 ( .INP(n2212), .Z(n378) );
  NBUFFX2 U1086 ( .INP(n2170), .Z(n34) );
  NBUFFX2 U1087 ( .INP(n2217), .Z(n550) );
  NBUFFX2 U1088 ( .INP(n2212), .Z(n379) );
  NBUFFX2 U1089 ( .INP(n2170), .Z(n35) );
  NBUFFX2 U1090 ( .INP(n2217), .Z(n551) );
  NBUFFX2 U1091 ( .INP(n2212), .Z(n380) );
  NBUFFX2 U1092 ( .INP(n2170), .Z(n36) );
  NBUFFX2 U1093 ( .INP(n2217), .Z(n552) );
  NBUFFX2 U1094 ( .INP(n2212), .Z(n381) );
  NBUFFX2 U1095 ( .INP(n2170), .Z(n37) );
  NBUFFX2 U1096 ( .INP(n2217), .Z(n553) );
  NBUFFX2 U1097 ( .INP(n2212), .Z(n382) );
  NBUFFX2 U1098 ( .INP(n2170), .Z(n38) );
  NBUFFX2 U1099 ( .INP(n2217), .Z(n554) );
  NBUFFX2 U1100 ( .INP(n2212), .Z(n383) );
  NBUFFX2 U1101 ( .INP(n2170), .Z(n39) );
  NBUFFX2 U1102 ( .INP(n2217), .Z(n555) );
  NBUFFX2 U1103 ( .INP(n2212), .Z(n384) );
  NBUFFX2 U1104 ( .INP(n2170), .Z(n40) );
  NBUFFX2 U1105 ( .INP(n2217), .Z(n556) );
  NBUFFX2 U1106 ( .INP(n2212), .Z(n385) );
  NBUFFX2 U1107 ( .INP(n2170), .Z(n41) );
  NBUFFX2 U1108 ( .INP(n2217), .Z(n557) );
  NBUFFX2 U1109 ( .INP(n2212), .Z(n386) );
  NBUFFX2 U1110 ( .INP(n2170), .Z(n42) );
  NBUFFX2 U1111 ( .INP(n2217), .Z(n558) );
  NBUFFX2 U1112 ( .INP(n2210), .Z(n301) );
  NBUFFX2 U1113 ( .INP(n2215), .Z(n473) );
  NBUFFX2 U1114 ( .INP(n2205), .Z(n129) );
  NBUFFX2 U1115 ( .INP(n2220), .Z(n645) );
  NBUFFX2 U1116 ( .INP(n2211), .Z(n344) );
  NBUFFX2 U1117 ( .INP(n2216), .Z(n516) );
  NBUFFX2 U1118 ( .INP(n2221), .Z(n688) );
  NBUFFX2 U1119 ( .INP(n2208), .Z(n258) );
  NBUFFX2 U1120 ( .INP(n2213), .Z(n430) );
  NBUFFX2 U1121 ( .INP(n2194), .Z(n86) );
  NBUFFX2 U1122 ( .INP(n2218), .Z(n602) );
  NBUFFX2 U1123 ( .INP(n2207), .Z(n215) );
  NBUFFX2 U1124 ( .INP(n2212), .Z(n387) );
  NBUFFX2 U1125 ( .INP(n2170), .Z(n43) );
  NBUFFX2 U1126 ( .INP(n2217), .Z(n559) );
  NBUFFX2 U1127 ( .INP(clk), .Z(n2151) );
  NBUFFX2 U1128 ( .INP(clk), .Z(n2150) );
  NBUFFX2 U1129 ( .INP(clk), .Z(n2149) );
  NBUFFX2 U1130 ( .INP(clk), .Z(n2148) );
  NBUFFX2 U1131 ( .INP(clk), .Z(n2147) );
  NBUFFX2 U1132 ( .INP(clk), .Z(n2146) );
  NBUFFX2 U1133 ( .INP(clk), .Z(n2145) );
  NBUFFX2 U1134 ( .INP(clk), .Z(n2144) );
  NBUFFX2 U1135 ( .INP(clk), .Z(n2152) );
  NBUFFX2 U1136 ( .INP(clk), .Z(n2138) );
  NBUFFX2 U1137 ( .INP(clk), .Z(n2137) );
  NBUFFX2 U1138 ( .INP(clk), .Z(n2136) );
  NBUFFX2 U1139 ( .INP(clk), .Z(n2135) );
  NBUFFX2 U1140 ( .INP(clk), .Z(n2134) );
  NBUFFX2 U1141 ( .INP(clk), .Z(n2142) );
  NBUFFX2 U1142 ( .INP(clk), .Z(n2141) );
  NBUFFX2 U1143 ( .INP(clk), .Z(n2140) );
  NBUFFX2 U1144 ( .INP(clk), .Z(n2139) );
  NBUFFX2 U1145 ( .INP(clk), .Z(n2143) );
  NBUFFX2 U1146 ( .INP(di[16]), .Z(n1061) );
  NBUFFX2 U1147 ( .INP(di[17]), .Z(n1083) );
  NBUFFX2 U1148 ( .INP(di[18]), .Z(n1105) );
  NBUFFX2 U1149 ( .INP(di[19]), .Z(n1127) );
  NBUFFX2 U1150 ( .INP(di[20]), .Z(n1149) );
  NBUFFX2 U1151 ( .INP(di[21]), .Z(n1171) );
  NBUFFX2 U1152 ( .INP(di[22]), .Z(n1193) );
  NBUFFX2 U1153 ( .INP(di[23]), .Z(n1215) );
  NBUFFX2 U1154 ( .INP(di[16]), .Z(n1060) );
  NBUFFX2 U1155 ( .INP(di[17]), .Z(n1082) );
  NBUFFX2 U1156 ( .INP(di[18]), .Z(n1104) );
  NBUFFX2 U1157 ( .INP(di[19]), .Z(n1126) );
  NBUFFX2 U1158 ( .INP(di[20]), .Z(n1148) );
  NBUFFX2 U1159 ( .INP(di[21]), .Z(n1170) );
  NBUFFX2 U1160 ( .INP(di[22]), .Z(n1192) );
  NBUFFX2 U1161 ( .INP(di[23]), .Z(n1214) );
  NBUFFX2 U1162 ( .INP(di[16]), .Z(n1059) );
  NBUFFX2 U1163 ( .INP(di[17]), .Z(n1081) );
  NBUFFX2 U1164 ( .INP(di[18]), .Z(n1103) );
  NBUFFX2 U1165 ( .INP(di[19]), .Z(n1125) );
  NBUFFX2 U1166 ( .INP(di[20]), .Z(n1147) );
  NBUFFX2 U1167 ( .INP(di[21]), .Z(n1169) );
  NBUFFX2 U1168 ( .INP(di[22]), .Z(n1191) );
  NBUFFX2 U1169 ( .INP(di[23]), .Z(n1213) );
  NBUFFX2 U1170 ( .INP(di[16]), .Z(n1058) );
  NBUFFX2 U1171 ( .INP(di[17]), .Z(n1080) );
  NBUFFX2 U1172 ( .INP(di[18]), .Z(n1102) );
  NBUFFX2 U1173 ( .INP(di[19]), .Z(n1124) );
  NBUFFX2 U1174 ( .INP(di[20]), .Z(n1146) );
  NBUFFX2 U1175 ( .INP(di[21]), .Z(n1168) );
  NBUFFX2 U1176 ( .INP(di[22]), .Z(n1190) );
  NBUFFX2 U1177 ( .INP(di[23]), .Z(n1212) );
  NBUFFX2 U1178 ( .INP(di[16]), .Z(n1057) );
  NBUFFX2 U1179 ( .INP(di[17]), .Z(n1079) );
  NBUFFX2 U1180 ( .INP(di[18]), .Z(n1101) );
  NBUFFX2 U1181 ( .INP(di[19]), .Z(n1123) );
  NBUFFX2 U1182 ( .INP(di[20]), .Z(n1145) );
  NBUFFX2 U1183 ( .INP(di[21]), .Z(n1167) );
  NBUFFX2 U1184 ( .INP(di[22]), .Z(n1189) );
  NBUFFX2 U1185 ( .INP(di[23]), .Z(n1211) );
  NBUFFX2 U1186 ( .INP(di[16]), .Z(n1056) );
  NBUFFX2 U1187 ( .INP(di[17]), .Z(n1078) );
  NBUFFX2 U1188 ( .INP(di[18]), .Z(n1100) );
  NBUFFX2 U1189 ( .INP(di[19]), .Z(n1122) );
  NBUFFX2 U1190 ( .INP(di[20]), .Z(n1144) );
  NBUFFX2 U1191 ( .INP(di[21]), .Z(n1166) );
  NBUFFX2 U1192 ( .INP(di[22]), .Z(n1188) );
  NBUFFX2 U1193 ( .INP(di[23]), .Z(n1210) );
  NBUFFX2 U1194 ( .INP(di[16]), .Z(n1055) );
  NBUFFX2 U1195 ( .INP(di[17]), .Z(n1077) );
  NBUFFX2 U1196 ( .INP(di[18]), .Z(n1099) );
  NBUFFX2 U1197 ( .INP(di[19]), .Z(n1121) );
  NBUFFX2 U1198 ( .INP(di[20]), .Z(n1143) );
  NBUFFX2 U1199 ( .INP(di[21]), .Z(n1165) );
  NBUFFX2 U1200 ( .INP(di[22]), .Z(n1187) );
  NBUFFX2 U1201 ( .INP(di[23]), .Z(n1209) );
  NBUFFX2 U1202 ( .INP(di[16]), .Z(n1054) );
  NBUFFX2 U1203 ( .INP(di[17]), .Z(n1076) );
  NBUFFX2 U1204 ( .INP(di[18]), .Z(n1098) );
  NBUFFX2 U1205 ( .INP(di[19]), .Z(n1120) );
  NBUFFX2 U1206 ( .INP(di[20]), .Z(n1142) );
  NBUFFX2 U1207 ( .INP(di[21]), .Z(n1164) );
  NBUFFX2 U1208 ( .INP(di[22]), .Z(n1186) );
  NBUFFX2 U1209 ( .INP(di[23]), .Z(n1208) );
  NBUFFX2 U1210 ( .INP(di[16]), .Z(n1053) );
  NBUFFX2 U1211 ( .INP(di[17]), .Z(n1075) );
  NBUFFX2 U1212 ( .INP(di[18]), .Z(n1097) );
  NBUFFX2 U1213 ( .INP(di[19]), .Z(n1119) );
  NBUFFX2 U1214 ( .INP(di[20]), .Z(n1141) );
  NBUFFX2 U1215 ( .INP(di[21]), .Z(n1163) );
  NBUFFX2 U1216 ( .INP(di[22]), .Z(n1185) );
  NBUFFX2 U1217 ( .INP(di[23]), .Z(n1207) );
  NBUFFX2 U1218 ( .INP(di[16]), .Z(n1052) );
  NBUFFX2 U1219 ( .INP(di[17]), .Z(n1074) );
  NBUFFX2 U1220 ( .INP(di[18]), .Z(n1096) );
  NBUFFX2 U1221 ( .INP(di[19]), .Z(n1118) );
  NBUFFX2 U1222 ( .INP(di[20]), .Z(n1140) );
  NBUFFX2 U1223 ( .INP(di[21]), .Z(n1162) );
  NBUFFX2 U1224 ( .INP(di[22]), .Z(n1184) );
  NBUFFX2 U1225 ( .INP(di[23]), .Z(n1206) );
  NBUFFX2 U1226 ( .INP(di[16]), .Z(n1051) );
  NBUFFX2 U1227 ( .INP(di[17]), .Z(n1073) );
  NBUFFX2 U1228 ( .INP(di[18]), .Z(n1095) );
  NBUFFX2 U1229 ( .INP(di[19]), .Z(n1117) );
  NBUFFX2 U1230 ( .INP(di[20]), .Z(n1139) );
  NBUFFX2 U1231 ( .INP(di[21]), .Z(n1161) );
  NBUFFX2 U1232 ( .INP(di[22]), .Z(n1183) );
  NBUFFX2 U1233 ( .INP(di[23]), .Z(n1205) );
  NBUFFX2 U1234 ( .INP(di[16]), .Z(n1050) );
  NBUFFX2 U1235 ( .INP(di[17]), .Z(n1072) );
  NBUFFX2 U1236 ( .INP(di[18]), .Z(n1094) );
  NBUFFX2 U1237 ( .INP(di[19]), .Z(n1116) );
  NBUFFX2 U1238 ( .INP(di[20]), .Z(n1138) );
  NBUFFX2 U1239 ( .INP(di[21]), .Z(n1160) );
  NBUFFX2 U1240 ( .INP(di[22]), .Z(n1182) );
  NBUFFX2 U1241 ( .INP(di[23]), .Z(n1204) );
  NBUFFX2 U1242 ( .INP(di[16]), .Z(n1049) );
  NBUFFX2 U1243 ( .INP(di[17]), .Z(n1071) );
  NBUFFX2 U1244 ( .INP(di[18]), .Z(n1093) );
  NBUFFX2 U1245 ( .INP(di[19]), .Z(n1115) );
  NBUFFX2 U1246 ( .INP(di[20]), .Z(n1137) );
  NBUFFX2 U1247 ( .INP(di[21]), .Z(n1159) );
  NBUFFX2 U1248 ( .INP(di[22]), .Z(n1181) );
  NBUFFX2 U1249 ( .INP(di[23]), .Z(n1203) );
  NBUFFX2 U1250 ( .INP(di[16]), .Z(n1048) );
  NBUFFX2 U1251 ( .INP(di[17]), .Z(n1070) );
  NBUFFX2 U1252 ( .INP(di[18]), .Z(n1092) );
  NBUFFX2 U1253 ( .INP(di[19]), .Z(n1114) );
  NBUFFX2 U1254 ( .INP(di[20]), .Z(n1136) );
  NBUFFX2 U1255 ( .INP(di[21]), .Z(n1158) );
  NBUFFX2 U1256 ( .INP(di[22]), .Z(n1180) );
  NBUFFX2 U1257 ( .INP(di[23]), .Z(n1202) );
  NBUFFX2 U1258 ( .INP(di[16]), .Z(n1047) );
  NBUFFX2 U1259 ( .INP(di[17]), .Z(n1069) );
  NBUFFX2 U1260 ( .INP(di[18]), .Z(n1091) );
  NBUFFX2 U1261 ( .INP(di[19]), .Z(n1113) );
  NBUFFX2 U1262 ( .INP(di[20]), .Z(n1135) );
  NBUFFX2 U1263 ( .INP(di[21]), .Z(n1157) );
  NBUFFX2 U1264 ( .INP(di[22]), .Z(n1179) );
  NBUFFX2 U1265 ( .INP(di[23]), .Z(n1201) );
  NBUFFX2 U1266 ( .INP(di[16]), .Z(n1046) );
  NBUFFX2 U1267 ( .INP(di[17]), .Z(n1068) );
  NBUFFX2 U1268 ( .INP(di[18]), .Z(n1090) );
  NBUFFX2 U1269 ( .INP(di[19]), .Z(n1112) );
  NBUFFX2 U1270 ( .INP(di[20]), .Z(n1134) );
  NBUFFX2 U1271 ( .INP(di[21]), .Z(n1156) );
  NBUFFX2 U1272 ( .INP(di[22]), .Z(n1178) );
  NBUFFX2 U1273 ( .INP(di[23]), .Z(n1200) );
  NBUFFX2 U1274 ( .INP(di[16]), .Z(n1045) );
  NBUFFX2 U1275 ( .INP(di[17]), .Z(n1067) );
  NBUFFX2 U1276 ( .INP(di[18]), .Z(n1089) );
  NBUFFX2 U1277 ( .INP(di[19]), .Z(n1111) );
  NBUFFX2 U1278 ( .INP(di[20]), .Z(n1133) );
  NBUFFX2 U1279 ( .INP(di[21]), .Z(n1155) );
  NBUFFX2 U1280 ( .INP(di[22]), .Z(n1177) );
  NBUFFX2 U1281 ( .INP(di[23]), .Z(n1199) );
  NBUFFX2 U1282 ( .INP(di[16]), .Z(n1044) );
  NBUFFX2 U1283 ( .INP(di[17]), .Z(n1066) );
  NBUFFX2 U1284 ( .INP(di[18]), .Z(n1088) );
  NBUFFX2 U1285 ( .INP(di[19]), .Z(n1110) );
  NBUFFX2 U1286 ( .INP(di[20]), .Z(n1132) );
  NBUFFX2 U1287 ( .INP(di[21]), .Z(n1154) );
  NBUFFX2 U1288 ( .INP(di[22]), .Z(n1176) );
  NBUFFX2 U1289 ( .INP(di[23]), .Z(n1198) );
  NBUFFX2 U1290 ( .INP(di[16]), .Z(n1043) );
  NBUFFX2 U1291 ( .INP(di[17]), .Z(n1065) );
  NBUFFX2 U1292 ( .INP(di[18]), .Z(n1087) );
  NBUFFX2 U1293 ( .INP(di[19]), .Z(n1109) );
  NBUFFX2 U1294 ( .INP(di[20]), .Z(n1131) );
  NBUFFX2 U1295 ( .INP(di[21]), .Z(n1153) );
  NBUFFX2 U1296 ( .INP(di[22]), .Z(n1175) );
  NBUFFX2 U1297 ( .INP(di[23]), .Z(n1197) );
  NBUFFX2 U1298 ( .INP(di[16]), .Z(n1042) );
  NBUFFX2 U1299 ( .INP(di[17]), .Z(n1064) );
  NBUFFX2 U1300 ( .INP(di[18]), .Z(n1086) );
  NBUFFX2 U1301 ( .INP(di[19]), .Z(n1108) );
  NBUFFX2 U1302 ( .INP(di[20]), .Z(n1130) );
  NBUFFX2 U1303 ( .INP(di[21]), .Z(n1152) );
  NBUFFX2 U1304 ( .INP(di[22]), .Z(n1174) );
  NBUFFX2 U1305 ( .INP(di[23]), .Z(n1196) );
  NBUFFX2 U1306 ( .INP(di[16]), .Z(n1041) );
  NBUFFX2 U1307 ( .INP(di[17]), .Z(n1063) );
  NBUFFX2 U1308 ( .INP(di[18]), .Z(n1085) );
  NBUFFX2 U1309 ( .INP(di[19]), .Z(n1107) );
  NBUFFX2 U1310 ( .INP(di[20]), .Z(n1129) );
  NBUFFX2 U1311 ( .INP(di[21]), .Z(n1151) );
  NBUFFX2 U1312 ( .INP(di[22]), .Z(n1173) );
  NBUFFX2 U1313 ( .INP(di[23]), .Z(n1195) );
  NBUFFX2 U1314 ( .INP(di[24]), .Z(n1237) );
  NBUFFX2 U1315 ( .INP(di[25]), .Z(n1259) );
  NBUFFX2 U1316 ( .INP(di[26]), .Z(n1281) );
  NBUFFX2 U1317 ( .INP(di[27]), .Z(n1303) );
  NBUFFX2 U1318 ( .INP(di[28]), .Z(n1325) );
  NBUFFX2 U1319 ( .INP(di[29]), .Z(n1347) );
  NBUFFX2 U1320 ( .INP(di[30]), .Z(n1369) );
  NBUFFX2 U1321 ( .INP(di[31]), .Z(n1391) );
  NBUFFX2 U1322 ( .INP(di[24]), .Z(n1236) );
  NBUFFX2 U1323 ( .INP(di[25]), .Z(n1258) );
  NBUFFX2 U1324 ( .INP(di[26]), .Z(n1280) );
  NBUFFX2 U1325 ( .INP(di[27]), .Z(n1302) );
  NBUFFX2 U1326 ( .INP(di[28]), .Z(n1324) );
  NBUFFX2 U1327 ( .INP(di[29]), .Z(n1346) );
  NBUFFX2 U1328 ( .INP(di[30]), .Z(n1368) );
  NBUFFX2 U1329 ( .INP(di[31]), .Z(n1390) );
  NBUFFX2 U1330 ( .INP(di[24]), .Z(n1235) );
  NBUFFX2 U1331 ( .INP(di[25]), .Z(n1257) );
  NBUFFX2 U1332 ( .INP(di[26]), .Z(n1279) );
  NBUFFX2 U1333 ( .INP(di[27]), .Z(n1301) );
  NBUFFX2 U1334 ( .INP(di[28]), .Z(n1323) );
  NBUFFX2 U1335 ( .INP(di[29]), .Z(n1345) );
  NBUFFX2 U1336 ( .INP(di[30]), .Z(n1367) );
  NBUFFX2 U1337 ( .INP(di[31]), .Z(n1389) );
  NBUFFX2 U1338 ( .INP(di[24]), .Z(n1234) );
  NBUFFX2 U1339 ( .INP(di[25]), .Z(n1256) );
  NBUFFX2 U1340 ( .INP(di[26]), .Z(n1278) );
  NBUFFX2 U1341 ( .INP(di[27]), .Z(n1300) );
  NBUFFX2 U1342 ( .INP(di[28]), .Z(n1322) );
  NBUFFX2 U1343 ( .INP(di[29]), .Z(n1344) );
  NBUFFX2 U1344 ( .INP(di[30]), .Z(n1366) );
  NBUFFX2 U1345 ( .INP(di[31]), .Z(n1388) );
  NBUFFX2 U1346 ( .INP(di[24]), .Z(n1233) );
  NBUFFX2 U1347 ( .INP(di[25]), .Z(n1255) );
  NBUFFX2 U1348 ( .INP(di[26]), .Z(n1277) );
  NBUFFX2 U1349 ( .INP(di[27]), .Z(n1299) );
  NBUFFX2 U1350 ( .INP(di[28]), .Z(n1321) );
  NBUFFX2 U1351 ( .INP(di[29]), .Z(n1343) );
  NBUFFX2 U1352 ( .INP(di[30]), .Z(n1365) );
  NBUFFX2 U1353 ( .INP(di[31]), .Z(n1387) );
  NBUFFX2 U1354 ( .INP(di[24]), .Z(n1232) );
  NBUFFX2 U1355 ( .INP(di[25]), .Z(n1254) );
  NBUFFX2 U1356 ( .INP(di[26]), .Z(n1276) );
  NBUFFX2 U1357 ( .INP(di[27]), .Z(n1298) );
  NBUFFX2 U1358 ( .INP(di[28]), .Z(n1320) );
  NBUFFX2 U1359 ( .INP(di[29]), .Z(n1342) );
  NBUFFX2 U1360 ( .INP(di[30]), .Z(n1364) );
  NBUFFX2 U1361 ( .INP(di[31]), .Z(n1386) );
  NBUFFX2 U1362 ( .INP(di[24]), .Z(n1231) );
  NBUFFX2 U1363 ( .INP(di[25]), .Z(n1253) );
  NBUFFX2 U1364 ( .INP(di[26]), .Z(n1275) );
  NBUFFX2 U1365 ( .INP(di[27]), .Z(n1297) );
  NBUFFX2 U1366 ( .INP(di[28]), .Z(n1319) );
  NBUFFX2 U1367 ( .INP(di[29]), .Z(n1341) );
  NBUFFX2 U1368 ( .INP(di[30]), .Z(n1363) );
  NBUFFX2 U1369 ( .INP(di[31]), .Z(n1385) );
  NBUFFX2 U1370 ( .INP(di[24]), .Z(n1230) );
  NBUFFX2 U1371 ( .INP(di[25]), .Z(n1252) );
  NBUFFX2 U1372 ( .INP(di[26]), .Z(n1274) );
  NBUFFX2 U1373 ( .INP(di[27]), .Z(n1296) );
  NBUFFX2 U1374 ( .INP(di[28]), .Z(n1318) );
  NBUFFX2 U1375 ( .INP(di[29]), .Z(n1340) );
  NBUFFX2 U1376 ( .INP(di[30]), .Z(n1362) );
  NBUFFX2 U1377 ( .INP(di[31]), .Z(n1384) );
  NBUFFX2 U1378 ( .INP(di[24]), .Z(n1229) );
  NBUFFX2 U1379 ( .INP(di[25]), .Z(n1251) );
  NBUFFX2 U1380 ( .INP(di[26]), .Z(n1273) );
  NBUFFX2 U1381 ( .INP(di[27]), .Z(n1295) );
  NBUFFX2 U1382 ( .INP(di[28]), .Z(n1317) );
  NBUFFX2 U1383 ( .INP(di[29]), .Z(n1339) );
  NBUFFX2 U1384 ( .INP(di[30]), .Z(n1361) );
  NBUFFX2 U1385 ( .INP(di[31]), .Z(n1383) );
  NBUFFX2 U1386 ( .INP(di[24]), .Z(n1228) );
  NBUFFX2 U1387 ( .INP(di[25]), .Z(n1250) );
  NBUFFX2 U1388 ( .INP(di[26]), .Z(n1272) );
  NBUFFX2 U1389 ( .INP(di[27]), .Z(n1294) );
  NBUFFX2 U1390 ( .INP(di[28]), .Z(n1316) );
  NBUFFX2 U1391 ( .INP(di[29]), .Z(n1338) );
  NBUFFX2 U1392 ( .INP(di[30]), .Z(n1360) );
  NBUFFX2 U1393 ( .INP(di[31]), .Z(n1382) );
  NBUFFX2 U1394 ( .INP(di[24]), .Z(n1227) );
  NBUFFX2 U1395 ( .INP(di[25]), .Z(n1249) );
  NBUFFX2 U1396 ( .INP(di[26]), .Z(n1271) );
  NBUFFX2 U1397 ( .INP(di[27]), .Z(n1293) );
  NBUFFX2 U1398 ( .INP(di[28]), .Z(n1315) );
  NBUFFX2 U1399 ( .INP(di[29]), .Z(n1337) );
  NBUFFX2 U1400 ( .INP(di[30]), .Z(n1359) );
  NBUFFX2 U1401 ( .INP(di[31]), .Z(n1381) );
  NBUFFX2 U1402 ( .INP(di[24]), .Z(n1226) );
  NBUFFX2 U1403 ( .INP(di[25]), .Z(n1248) );
  NBUFFX2 U1404 ( .INP(di[26]), .Z(n1270) );
  NBUFFX2 U1405 ( .INP(di[27]), .Z(n1292) );
  NBUFFX2 U1406 ( .INP(di[28]), .Z(n1314) );
  NBUFFX2 U1407 ( .INP(di[29]), .Z(n1336) );
  NBUFFX2 U1408 ( .INP(di[30]), .Z(n1358) );
  NBUFFX2 U1409 ( .INP(di[31]), .Z(n1380) );
  NBUFFX2 U1410 ( .INP(di[24]), .Z(n1225) );
  NBUFFX2 U1411 ( .INP(di[25]), .Z(n1247) );
  NBUFFX2 U1412 ( .INP(di[26]), .Z(n1269) );
  NBUFFX2 U1413 ( .INP(di[27]), .Z(n1291) );
  NBUFFX2 U1414 ( .INP(di[28]), .Z(n1313) );
  NBUFFX2 U1415 ( .INP(di[29]), .Z(n1335) );
  NBUFFX2 U1416 ( .INP(di[30]), .Z(n1357) );
  NBUFFX2 U1417 ( .INP(di[31]), .Z(n1379) );
  NBUFFX2 U1418 ( .INP(di[24]), .Z(n1224) );
  NBUFFX2 U1419 ( .INP(di[25]), .Z(n1246) );
  NBUFFX2 U1420 ( .INP(di[26]), .Z(n1268) );
  NBUFFX2 U1421 ( .INP(di[27]), .Z(n1290) );
  NBUFFX2 U1422 ( .INP(di[28]), .Z(n1312) );
  NBUFFX2 U1423 ( .INP(di[29]), .Z(n1334) );
  NBUFFX2 U1424 ( .INP(di[30]), .Z(n1356) );
  NBUFFX2 U1425 ( .INP(di[31]), .Z(n1378) );
  NBUFFX2 U1426 ( .INP(di[24]), .Z(n1223) );
  NBUFFX2 U1427 ( .INP(di[25]), .Z(n1245) );
  NBUFFX2 U1428 ( .INP(di[26]), .Z(n1267) );
  NBUFFX2 U1429 ( .INP(di[27]), .Z(n1289) );
  NBUFFX2 U1430 ( .INP(di[28]), .Z(n1311) );
  NBUFFX2 U1431 ( .INP(di[29]), .Z(n1333) );
  NBUFFX2 U1432 ( .INP(di[30]), .Z(n1355) );
  NBUFFX2 U1433 ( .INP(di[31]), .Z(n1377) );
  NBUFFX2 U1434 ( .INP(di[24]), .Z(n1222) );
  NBUFFX2 U1435 ( .INP(di[25]), .Z(n1244) );
  NBUFFX2 U1436 ( .INP(di[26]), .Z(n1266) );
  NBUFFX2 U1437 ( .INP(di[27]), .Z(n1288) );
  NBUFFX2 U1438 ( .INP(di[28]), .Z(n1310) );
  NBUFFX2 U1439 ( .INP(di[29]), .Z(n1332) );
  NBUFFX2 U1440 ( .INP(di[30]), .Z(n1354) );
  NBUFFX2 U1441 ( .INP(di[31]), .Z(n1376) );
  NBUFFX2 U1442 ( .INP(di[24]), .Z(n1221) );
  NBUFFX2 U1443 ( .INP(di[25]), .Z(n1243) );
  NBUFFX2 U1444 ( .INP(di[26]), .Z(n1265) );
  NBUFFX2 U1445 ( .INP(di[27]), .Z(n1287) );
  NBUFFX2 U1446 ( .INP(di[28]), .Z(n1309) );
  NBUFFX2 U1447 ( .INP(di[29]), .Z(n1331) );
  NBUFFX2 U1448 ( .INP(di[30]), .Z(n1353) );
  NBUFFX2 U1449 ( .INP(di[31]), .Z(n1375) );
  NBUFFX2 U1450 ( .INP(di[24]), .Z(n1220) );
  NBUFFX2 U1451 ( .INP(di[25]), .Z(n1242) );
  NBUFFX2 U1452 ( .INP(di[26]), .Z(n1264) );
  NBUFFX2 U1453 ( .INP(di[27]), .Z(n1286) );
  NBUFFX2 U1454 ( .INP(di[28]), .Z(n1308) );
  NBUFFX2 U1455 ( .INP(di[29]), .Z(n1330) );
  NBUFFX2 U1456 ( .INP(di[30]), .Z(n1352) );
  NBUFFX2 U1457 ( .INP(di[31]), .Z(n1374) );
  NBUFFX2 U1458 ( .INP(di[24]), .Z(n1219) );
  NBUFFX2 U1459 ( .INP(di[25]), .Z(n1241) );
  NBUFFX2 U1460 ( .INP(di[26]), .Z(n1263) );
  NBUFFX2 U1461 ( .INP(di[27]), .Z(n1285) );
  NBUFFX2 U1462 ( .INP(di[28]), .Z(n1307) );
  NBUFFX2 U1463 ( .INP(di[29]), .Z(n1329) );
  NBUFFX2 U1464 ( .INP(di[30]), .Z(n1351) );
  NBUFFX2 U1465 ( .INP(di[31]), .Z(n1373) );
  NBUFFX2 U1466 ( .INP(di[24]), .Z(n1218) );
  NBUFFX2 U1467 ( .INP(di[25]), .Z(n1240) );
  NBUFFX2 U1468 ( .INP(di[26]), .Z(n1262) );
  NBUFFX2 U1469 ( .INP(di[27]), .Z(n1284) );
  NBUFFX2 U1470 ( .INP(di[28]), .Z(n1306) );
  NBUFFX2 U1471 ( .INP(di[29]), .Z(n1328) );
  NBUFFX2 U1472 ( .INP(di[30]), .Z(n1350) );
  NBUFFX2 U1473 ( .INP(di[31]), .Z(n1372) );
  NBUFFX2 U1474 ( .INP(di[24]), .Z(n1217) );
  NBUFFX2 U1475 ( .INP(di[25]), .Z(n1239) );
  NBUFFX2 U1476 ( .INP(di[26]), .Z(n1261) );
  NBUFFX2 U1477 ( .INP(di[27]), .Z(n1283) );
  NBUFFX2 U1478 ( .INP(di[28]), .Z(n1305) );
  NBUFFX2 U1479 ( .INP(di[29]), .Z(n1327) );
  NBUFFX2 U1480 ( .INP(di[30]), .Z(n1349) );
  NBUFFX2 U1481 ( .INP(di[31]), .Z(n1371) );
  NBUFFX2 U1482 ( .INP(di[8]), .Z(n885) );
  NBUFFX2 U1483 ( .INP(di[9]), .Z(n907) );
  NBUFFX2 U1484 ( .INP(di[10]), .Z(n929) );
  NBUFFX2 U1485 ( .INP(di[11]), .Z(n951) );
  NBUFFX2 U1486 ( .INP(di[12]), .Z(n973) );
  NBUFFX2 U1487 ( .INP(di[13]), .Z(n995) );
  NBUFFX2 U1488 ( .INP(di[14]), .Z(n1017) );
  NBUFFX2 U1489 ( .INP(di[15]), .Z(n1039) );
  NBUFFX2 U1490 ( .INP(di[8]), .Z(n884) );
  NBUFFX2 U1491 ( .INP(di[9]), .Z(n906) );
  NBUFFX2 U1492 ( .INP(di[10]), .Z(n928) );
  NBUFFX2 U1493 ( .INP(di[11]), .Z(n950) );
  NBUFFX2 U1494 ( .INP(di[12]), .Z(n972) );
  NBUFFX2 U1495 ( .INP(di[13]), .Z(n994) );
  NBUFFX2 U1496 ( .INP(di[14]), .Z(n1016) );
  NBUFFX2 U1497 ( .INP(di[15]), .Z(n1038) );
  NBUFFX2 U1498 ( .INP(di[8]), .Z(n883) );
  NBUFFX2 U1499 ( .INP(di[9]), .Z(n905) );
  NBUFFX2 U1500 ( .INP(di[10]), .Z(n927) );
  NBUFFX2 U1501 ( .INP(di[11]), .Z(n949) );
  NBUFFX2 U1502 ( .INP(di[12]), .Z(n971) );
  NBUFFX2 U1503 ( .INP(di[13]), .Z(n993) );
  NBUFFX2 U1504 ( .INP(di[14]), .Z(n1015) );
  NBUFFX2 U1505 ( .INP(di[15]), .Z(n1037) );
  NBUFFX2 U1506 ( .INP(di[8]), .Z(n882) );
  NBUFFX2 U1507 ( .INP(di[9]), .Z(n904) );
  NBUFFX2 U1508 ( .INP(di[10]), .Z(n926) );
  NBUFFX2 U1509 ( .INP(di[11]), .Z(n948) );
  NBUFFX2 U1510 ( .INP(di[12]), .Z(n970) );
  NBUFFX2 U1511 ( .INP(di[13]), .Z(n992) );
  NBUFFX2 U1512 ( .INP(di[14]), .Z(n1014) );
  NBUFFX2 U1513 ( .INP(di[15]), .Z(n1036) );
  NBUFFX2 U1514 ( .INP(di[8]), .Z(n881) );
  NBUFFX2 U1515 ( .INP(di[9]), .Z(n903) );
  NBUFFX2 U1516 ( .INP(di[10]), .Z(n925) );
  NBUFFX2 U1517 ( .INP(di[11]), .Z(n947) );
  NBUFFX2 U1518 ( .INP(di[12]), .Z(n969) );
  NBUFFX2 U1519 ( .INP(di[13]), .Z(n991) );
  NBUFFX2 U1520 ( .INP(di[14]), .Z(n1013) );
  NBUFFX2 U1521 ( .INP(di[15]), .Z(n1035) );
  NBUFFX2 U1522 ( .INP(di[8]), .Z(n880) );
  NBUFFX2 U1523 ( .INP(di[9]), .Z(n902) );
  NBUFFX2 U1524 ( .INP(di[10]), .Z(n924) );
  NBUFFX2 U1525 ( .INP(di[11]), .Z(n946) );
  NBUFFX2 U1526 ( .INP(di[12]), .Z(n968) );
  NBUFFX2 U1527 ( .INP(di[13]), .Z(n990) );
  NBUFFX2 U1528 ( .INP(di[14]), .Z(n1012) );
  NBUFFX2 U1529 ( .INP(di[15]), .Z(n1034) );
  NBUFFX2 U1530 ( .INP(di[8]), .Z(n879) );
  NBUFFX2 U1531 ( .INP(di[9]), .Z(n901) );
  NBUFFX2 U1532 ( .INP(di[10]), .Z(n923) );
  NBUFFX2 U1533 ( .INP(di[11]), .Z(n945) );
  NBUFFX2 U1534 ( .INP(di[12]), .Z(n967) );
  NBUFFX2 U1535 ( .INP(di[13]), .Z(n989) );
  NBUFFX2 U1536 ( .INP(di[14]), .Z(n1011) );
  NBUFFX2 U1537 ( .INP(di[15]), .Z(n1033) );
  NBUFFX2 U1538 ( .INP(di[8]), .Z(n878) );
  NBUFFX2 U1539 ( .INP(di[9]), .Z(n900) );
  NBUFFX2 U1540 ( .INP(di[10]), .Z(n922) );
  NBUFFX2 U1541 ( .INP(di[11]), .Z(n944) );
  NBUFFX2 U1542 ( .INP(di[12]), .Z(n966) );
  NBUFFX2 U1543 ( .INP(di[13]), .Z(n988) );
  NBUFFX2 U1544 ( .INP(di[14]), .Z(n1010) );
  NBUFFX2 U1545 ( .INP(di[15]), .Z(n1032) );
  NBUFFX2 U1546 ( .INP(di[8]), .Z(n877) );
  NBUFFX2 U1547 ( .INP(di[9]), .Z(n899) );
  NBUFFX2 U1548 ( .INP(di[10]), .Z(n921) );
  NBUFFX2 U1549 ( .INP(di[11]), .Z(n943) );
  NBUFFX2 U1550 ( .INP(di[12]), .Z(n965) );
  NBUFFX2 U1551 ( .INP(di[13]), .Z(n987) );
  NBUFFX2 U1552 ( .INP(di[14]), .Z(n1009) );
  NBUFFX2 U1553 ( .INP(di[15]), .Z(n1031) );
  NBUFFX2 U1554 ( .INP(di[8]), .Z(n876) );
  NBUFFX2 U1555 ( .INP(di[9]), .Z(n898) );
  NBUFFX2 U1556 ( .INP(di[10]), .Z(n920) );
  NBUFFX2 U1557 ( .INP(di[11]), .Z(n942) );
  NBUFFX2 U1558 ( .INP(di[12]), .Z(n964) );
  NBUFFX2 U1559 ( .INP(di[13]), .Z(n986) );
  NBUFFX2 U1560 ( .INP(di[14]), .Z(n1008) );
  NBUFFX2 U1561 ( .INP(di[15]), .Z(n1030) );
  NBUFFX2 U1562 ( .INP(di[8]), .Z(n875) );
  NBUFFX2 U1563 ( .INP(di[9]), .Z(n897) );
  NBUFFX2 U1564 ( .INP(di[10]), .Z(n919) );
  NBUFFX2 U1565 ( .INP(di[11]), .Z(n941) );
  NBUFFX2 U1566 ( .INP(di[12]), .Z(n963) );
  NBUFFX2 U1567 ( .INP(di[13]), .Z(n985) );
  NBUFFX2 U1568 ( .INP(di[14]), .Z(n1007) );
  NBUFFX2 U1569 ( .INP(di[15]), .Z(n1029) );
  NBUFFX2 U1570 ( .INP(di[8]), .Z(n874) );
  NBUFFX2 U1571 ( .INP(di[9]), .Z(n896) );
  NBUFFX2 U1572 ( .INP(di[10]), .Z(n918) );
  NBUFFX2 U1573 ( .INP(di[11]), .Z(n940) );
  NBUFFX2 U1574 ( .INP(di[12]), .Z(n962) );
  NBUFFX2 U1575 ( .INP(di[13]), .Z(n984) );
  NBUFFX2 U1576 ( .INP(di[14]), .Z(n1006) );
  NBUFFX2 U1577 ( .INP(di[15]), .Z(n1028) );
  NBUFFX2 U1578 ( .INP(di[8]), .Z(n873) );
  NBUFFX2 U1579 ( .INP(di[9]), .Z(n895) );
  NBUFFX2 U1580 ( .INP(di[10]), .Z(n917) );
  NBUFFX2 U1581 ( .INP(di[11]), .Z(n939) );
  NBUFFX2 U1582 ( .INP(di[12]), .Z(n961) );
  NBUFFX2 U1583 ( .INP(di[13]), .Z(n983) );
  NBUFFX2 U1584 ( .INP(di[14]), .Z(n1005) );
  NBUFFX2 U1585 ( .INP(di[15]), .Z(n1027) );
  NBUFFX2 U1586 ( .INP(di[8]), .Z(n872) );
  NBUFFX2 U1587 ( .INP(di[9]), .Z(n894) );
  NBUFFX2 U1588 ( .INP(di[10]), .Z(n916) );
  NBUFFX2 U1589 ( .INP(di[11]), .Z(n938) );
  NBUFFX2 U1590 ( .INP(di[12]), .Z(n960) );
  NBUFFX2 U1591 ( .INP(di[13]), .Z(n982) );
  NBUFFX2 U1592 ( .INP(di[14]), .Z(n1004) );
  NBUFFX2 U1593 ( .INP(di[15]), .Z(n1026) );
  NBUFFX2 U1594 ( .INP(di[8]), .Z(n871) );
  NBUFFX2 U1595 ( .INP(di[9]), .Z(n893) );
  NBUFFX2 U1596 ( .INP(di[10]), .Z(n915) );
  NBUFFX2 U1597 ( .INP(di[11]), .Z(n937) );
  NBUFFX2 U1598 ( .INP(di[12]), .Z(n959) );
  NBUFFX2 U1599 ( .INP(di[13]), .Z(n981) );
  NBUFFX2 U1600 ( .INP(di[14]), .Z(n1003) );
  NBUFFX2 U1601 ( .INP(di[15]), .Z(n1025) );
  NBUFFX2 U1602 ( .INP(di[8]), .Z(n870) );
  NBUFFX2 U1603 ( .INP(di[9]), .Z(n892) );
  NBUFFX2 U1604 ( .INP(di[10]), .Z(n914) );
  NBUFFX2 U1605 ( .INP(di[11]), .Z(n936) );
  NBUFFX2 U1606 ( .INP(di[12]), .Z(n958) );
  NBUFFX2 U1607 ( .INP(di[13]), .Z(n980) );
  NBUFFX2 U1608 ( .INP(di[14]), .Z(n1002) );
  NBUFFX2 U1609 ( .INP(di[15]), .Z(n1024) );
  NBUFFX2 U1610 ( .INP(di[8]), .Z(n869) );
  NBUFFX2 U1611 ( .INP(di[9]), .Z(n891) );
  NBUFFX2 U1612 ( .INP(di[10]), .Z(n913) );
  NBUFFX2 U1613 ( .INP(di[11]), .Z(n935) );
  NBUFFX2 U1614 ( .INP(di[12]), .Z(n957) );
  NBUFFX2 U1615 ( .INP(di[13]), .Z(n979) );
  NBUFFX2 U1616 ( .INP(di[14]), .Z(n1001) );
  NBUFFX2 U1617 ( .INP(di[15]), .Z(n1023) );
  NBUFFX2 U1618 ( .INP(di[8]), .Z(n868) );
  NBUFFX2 U1619 ( .INP(di[9]), .Z(n890) );
  NBUFFX2 U1620 ( .INP(di[10]), .Z(n912) );
  NBUFFX2 U1621 ( .INP(di[11]), .Z(n934) );
  NBUFFX2 U1622 ( .INP(di[12]), .Z(n956) );
  NBUFFX2 U1623 ( .INP(di[13]), .Z(n978) );
  NBUFFX2 U1624 ( .INP(di[14]), .Z(n1000) );
  NBUFFX2 U1625 ( .INP(di[15]), .Z(n1022) );
  NBUFFX2 U1626 ( .INP(di[8]), .Z(n867) );
  NBUFFX2 U1627 ( .INP(di[9]), .Z(n889) );
  NBUFFX2 U1628 ( .INP(di[10]), .Z(n911) );
  NBUFFX2 U1629 ( .INP(di[11]), .Z(n933) );
  NBUFFX2 U1630 ( .INP(di[12]), .Z(n955) );
  NBUFFX2 U1631 ( .INP(di[13]), .Z(n977) );
  NBUFFX2 U1632 ( .INP(di[14]), .Z(n999) );
  NBUFFX2 U1633 ( .INP(di[15]), .Z(n1021) );
  NBUFFX2 U1634 ( .INP(di[8]), .Z(n866) );
  NBUFFX2 U1635 ( .INP(di[9]), .Z(n888) );
  NBUFFX2 U1636 ( .INP(di[10]), .Z(n910) );
  NBUFFX2 U1637 ( .INP(di[11]), .Z(n932) );
  NBUFFX2 U1638 ( .INP(di[12]), .Z(n954) );
  NBUFFX2 U1639 ( .INP(di[13]), .Z(n976) );
  NBUFFX2 U1640 ( .INP(di[14]), .Z(n998) );
  NBUFFX2 U1641 ( .INP(di[15]), .Z(n1020) );
  NBUFFX2 U1642 ( .INP(di[8]), .Z(n865) );
  NBUFFX2 U1643 ( .INP(di[9]), .Z(n887) );
  NBUFFX2 U1644 ( .INP(di[10]), .Z(n909) );
  NBUFFX2 U1645 ( .INP(di[11]), .Z(n931) );
  NBUFFX2 U1646 ( .INP(di[12]), .Z(n953) );
  NBUFFX2 U1647 ( .INP(di[13]), .Z(n975) );
  NBUFFX2 U1648 ( .INP(di[14]), .Z(n997) );
  NBUFFX2 U1649 ( .INP(di[15]), .Z(n1019) );
  NBUFFX2 U1650 ( .INP(di[0]), .Z(n709) );
  NBUFFX2 U1651 ( .INP(di[1]), .Z(n731) );
  NBUFFX2 U1652 ( .INP(di[2]), .Z(n753) );
  NBUFFX2 U1653 ( .INP(di[3]), .Z(n775) );
  NBUFFX2 U1654 ( .INP(di[4]), .Z(n797) );
  NBUFFX2 U1655 ( .INP(di[5]), .Z(n819) );
  NBUFFX2 U1656 ( .INP(di[6]), .Z(n841) );
  NBUFFX2 U1657 ( .INP(di[7]), .Z(n863) );
  NBUFFX2 U1658 ( .INP(di[0]), .Z(n708) );
  NBUFFX2 U1659 ( .INP(di[1]), .Z(n730) );
  NBUFFX2 U1660 ( .INP(di[2]), .Z(n752) );
  NBUFFX2 U1661 ( .INP(di[3]), .Z(n774) );
  NBUFFX2 U1662 ( .INP(di[4]), .Z(n796) );
  NBUFFX2 U1663 ( .INP(di[5]), .Z(n818) );
  NBUFFX2 U1664 ( .INP(di[6]), .Z(n840) );
  NBUFFX2 U1665 ( .INP(di[7]), .Z(n862) );
  NBUFFX2 U1666 ( .INP(di[0]), .Z(n707) );
  NBUFFX2 U1667 ( .INP(di[1]), .Z(n729) );
  NBUFFX2 U1668 ( .INP(di[2]), .Z(n751) );
  NBUFFX2 U1669 ( .INP(di[3]), .Z(n773) );
  NBUFFX2 U1670 ( .INP(di[4]), .Z(n795) );
  NBUFFX2 U1671 ( .INP(di[5]), .Z(n817) );
  NBUFFX2 U1672 ( .INP(di[6]), .Z(n839) );
  NBUFFX2 U1673 ( .INP(di[7]), .Z(n861) );
  NBUFFX2 U1674 ( .INP(di[0]), .Z(n706) );
  NBUFFX2 U1675 ( .INP(di[1]), .Z(n728) );
  NBUFFX2 U1676 ( .INP(di[2]), .Z(n750) );
  NBUFFX2 U1677 ( .INP(di[3]), .Z(n772) );
  NBUFFX2 U1678 ( .INP(di[4]), .Z(n794) );
  NBUFFX2 U1679 ( .INP(di[5]), .Z(n816) );
  NBUFFX2 U1680 ( .INP(di[6]), .Z(n838) );
  NBUFFX2 U1681 ( .INP(di[7]), .Z(n860) );
  NBUFFX2 U1682 ( .INP(di[0]), .Z(n705) );
  NBUFFX2 U1683 ( .INP(di[1]), .Z(n727) );
  NBUFFX2 U1684 ( .INP(di[2]), .Z(n749) );
  NBUFFX2 U1685 ( .INP(di[3]), .Z(n771) );
  NBUFFX2 U1686 ( .INP(di[4]), .Z(n793) );
  NBUFFX2 U1687 ( .INP(di[5]), .Z(n815) );
  NBUFFX2 U1688 ( .INP(di[6]), .Z(n837) );
  NBUFFX2 U1689 ( .INP(di[7]), .Z(n859) );
  NBUFFX2 U1690 ( .INP(di[0]), .Z(n704) );
  NBUFFX2 U1691 ( .INP(di[1]), .Z(n726) );
  NBUFFX2 U1692 ( .INP(di[2]), .Z(n748) );
  NBUFFX2 U1693 ( .INP(di[3]), .Z(n770) );
  NBUFFX2 U1694 ( .INP(di[4]), .Z(n792) );
  NBUFFX2 U1695 ( .INP(di[5]), .Z(n814) );
  NBUFFX2 U1696 ( .INP(di[6]), .Z(n836) );
  NBUFFX2 U1697 ( .INP(di[7]), .Z(n858) );
  NBUFFX2 U1698 ( .INP(di[0]), .Z(n703) );
  NBUFFX2 U1699 ( .INP(di[1]), .Z(n725) );
  NBUFFX2 U1700 ( .INP(di[2]), .Z(n747) );
  NBUFFX2 U1701 ( .INP(di[3]), .Z(n769) );
  NBUFFX2 U1702 ( .INP(di[4]), .Z(n791) );
  NBUFFX2 U1703 ( .INP(di[5]), .Z(n813) );
  NBUFFX2 U1704 ( .INP(di[6]), .Z(n835) );
  NBUFFX2 U1705 ( .INP(di[7]), .Z(n857) );
  NBUFFX2 U1706 ( .INP(di[0]), .Z(n702) );
  NBUFFX2 U1707 ( .INP(di[1]), .Z(n724) );
  NBUFFX2 U1708 ( .INP(di[2]), .Z(n746) );
  NBUFFX2 U1709 ( .INP(di[3]), .Z(n768) );
  NBUFFX2 U1710 ( .INP(di[4]), .Z(n790) );
  NBUFFX2 U1711 ( .INP(di[5]), .Z(n812) );
  NBUFFX2 U1712 ( .INP(di[6]), .Z(n834) );
  NBUFFX2 U1713 ( .INP(di[7]), .Z(n856) );
  NBUFFX2 U1714 ( .INP(di[0]), .Z(n701) );
  NBUFFX2 U1715 ( .INP(di[1]), .Z(n723) );
  NBUFFX2 U1716 ( .INP(di[2]), .Z(n745) );
  NBUFFX2 U1717 ( .INP(di[3]), .Z(n767) );
  NBUFFX2 U1718 ( .INP(di[4]), .Z(n789) );
  NBUFFX2 U1719 ( .INP(di[5]), .Z(n811) );
  NBUFFX2 U1720 ( .INP(di[6]), .Z(n833) );
  NBUFFX2 U1721 ( .INP(di[7]), .Z(n855) );
  NBUFFX2 U1722 ( .INP(di[0]), .Z(n700) );
  NBUFFX2 U1723 ( .INP(di[1]), .Z(n722) );
  NBUFFX2 U1724 ( .INP(di[2]), .Z(n744) );
  NBUFFX2 U1725 ( .INP(di[3]), .Z(n766) );
  NBUFFX2 U1726 ( .INP(di[4]), .Z(n788) );
  NBUFFX2 U1727 ( .INP(di[5]), .Z(n810) );
  NBUFFX2 U1728 ( .INP(di[6]), .Z(n832) );
  NBUFFX2 U1729 ( .INP(di[7]), .Z(n854) );
  NBUFFX2 U1730 ( .INP(di[0]), .Z(n699) );
  NBUFFX2 U1731 ( .INP(di[1]), .Z(n721) );
  NBUFFX2 U1732 ( .INP(di[2]), .Z(n743) );
  NBUFFX2 U1733 ( .INP(di[3]), .Z(n765) );
  NBUFFX2 U1734 ( .INP(di[4]), .Z(n787) );
  NBUFFX2 U1735 ( .INP(di[5]), .Z(n809) );
  NBUFFX2 U1736 ( .INP(di[6]), .Z(n831) );
  NBUFFX2 U1737 ( .INP(di[7]), .Z(n853) );
  NBUFFX2 U1738 ( .INP(di[0]), .Z(n698) );
  NBUFFX2 U1739 ( .INP(di[1]), .Z(n720) );
  NBUFFX2 U1740 ( .INP(di[2]), .Z(n742) );
  NBUFFX2 U1741 ( .INP(di[3]), .Z(n764) );
  NBUFFX2 U1742 ( .INP(di[4]), .Z(n786) );
  NBUFFX2 U1743 ( .INP(di[5]), .Z(n808) );
  NBUFFX2 U1744 ( .INP(di[6]), .Z(n830) );
  NBUFFX2 U1745 ( .INP(di[7]), .Z(n852) );
  NBUFFX2 U1746 ( .INP(di[0]), .Z(n697) );
  NBUFFX2 U1747 ( .INP(di[1]), .Z(n719) );
  NBUFFX2 U1748 ( .INP(di[2]), .Z(n741) );
  NBUFFX2 U1749 ( .INP(di[3]), .Z(n763) );
  NBUFFX2 U1750 ( .INP(di[4]), .Z(n785) );
  NBUFFX2 U1751 ( .INP(di[5]), .Z(n807) );
  NBUFFX2 U1752 ( .INP(di[6]), .Z(n829) );
  NBUFFX2 U1753 ( .INP(di[7]), .Z(n851) );
  NBUFFX2 U1754 ( .INP(di[0]), .Z(n696) );
  NBUFFX2 U1755 ( .INP(di[1]), .Z(n718) );
  NBUFFX2 U1756 ( .INP(di[2]), .Z(n740) );
  NBUFFX2 U1757 ( .INP(di[3]), .Z(n762) );
  NBUFFX2 U1758 ( .INP(di[4]), .Z(n784) );
  NBUFFX2 U1759 ( .INP(di[5]), .Z(n806) );
  NBUFFX2 U1760 ( .INP(di[6]), .Z(n828) );
  NBUFFX2 U1761 ( .INP(di[7]), .Z(n850) );
  NBUFFX2 U1762 ( .INP(di[0]), .Z(n695) );
  NBUFFX2 U1763 ( .INP(di[1]), .Z(n717) );
  NBUFFX2 U1764 ( .INP(di[2]), .Z(n739) );
  NBUFFX2 U1765 ( .INP(di[3]), .Z(n761) );
  NBUFFX2 U1766 ( .INP(di[4]), .Z(n783) );
  NBUFFX2 U1767 ( .INP(di[5]), .Z(n805) );
  NBUFFX2 U1768 ( .INP(di[6]), .Z(n827) );
  NBUFFX2 U1769 ( .INP(di[7]), .Z(n849) );
  NBUFFX2 U1770 ( .INP(di[0]), .Z(n694) );
  NBUFFX2 U1771 ( .INP(di[1]), .Z(n716) );
  NBUFFX2 U1772 ( .INP(di[2]), .Z(n738) );
  NBUFFX2 U1773 ( .INP(di[3]), .Z(n760) );
  NBUFFX2 U1774 ( .INP(di[4]), .Z(n782) );
  NBUFFX2 U1775 ( .INP(di[5]), .Z(n804) );
  NBUFFX2 U1776 ( .INP(di[6]), .Z(n826) );
  NBUFFX2 U1777 ( .INP(di[7]), .Z(n848) );
  NBUFFX2 U1778 ( .INP(di[0]), .Z(n693) );
  NBUFFX2 U1779 ( .INP(di[1]), .Z(n715) );
  NBUFFX2 U1780 ( .INP(di[2]), .Z(n737) );
  NBUFFX2 U1781 ( .INP(di[3]), .Z(n759) );
  NBUFFX2 U1782 ( .INP(di[4]), .Z(n781) );
  NBUFFX2 U1783 ( .INP(di[5]), .Z(n803) );
  NBUFFX2 U1784 ( .INP(di[6]), .Z(n825) );
  NBUFFX2 U1785 ( .INP(di[7]), .Z(n847) );
  NBUFFX2 U1786 ( .INP(di[0]), .Z(n692) );
  NBUFFX2 U1787 ( .INP(di[1]), .Z(n714) );
  NBUFFX2 U1788 ( .INP(di[2]), .Z(n736) );
  NBUFFX2 U1789 ( .INP(di[3]), .Z(n758) );
  NBUFFX2 U1790 ( .INP(di[4]), .Z(n780) );
  NBUFFX2 U1791 ( .INP(di[5]), .Z(n802) );
  NBUFFX2 U1792 ( .INP(di[6]), .Z(n824) );
  NBUFFX2 U1793 ( .INP(di[7]), .Z(n846) );
  NBUFFX2 U1794 ( .INP(di[0]), .Z(n691) );
  NBUFFX2 U1795 ( .INP(di[1]), .Z(n713) );
  NBUFFX2 U1796 ( .INP(di[2]), .Z(n735) );
  NBUFFX2 U1797 ( .INP(di[3]), .Z(n757) );
  NBUFFX2 U1798 ( .INP(di[4]), .Z(n779) );
  NBUFFX2 U1799 ( .INP(di[5]), .Z(n801) );
  NBUFFX2 U1800 ( .INP(di[6]), .Z(n823) );
  NBUFFX2 U1801 ( .INP(di[7]), .Z(n845) );
  NBUFFX2 U1802 ( .INP(di[0]), .Z(n690) );
  NBUFFX2 U1803 ( .INP(di[1]), .Z(n712) );
  NBUFFX2 U1804 ( .INP(di[2]), .Z(n734) );
  NBUFFX2 U1805 ( .INP(di[3]), .Z(n756) );
  NBUFFX2 U1806 ( .INP(di[4]), .Z(n778) );
  NBUFFX2 U1807 ( .INP(di[5]), .Z(n800) );
  NBUFFX2 U1808 ( .INP(di[6]), .Z(n822) );
  NBUFFX2 U1809 ( .INP(di[7]), .Z(n844) );
  NBUFFX2 U1810 ( .INP(di[0]), .Z(n689) );
  NBUFFX2 U1811 ( .INP(di[1]), .Z(n711) );
  NBUFFX2 U1812 ( .INP(di[2]), .Z(n733) );
  NBUFFX2 U1813 ( .INP(di[3]), .Z(n755) );
  NBUFFX2 U1814 ( .INP(di[4]), .Z(n777) );
  NBUFFX2 U1815 ( .INP(di[5]), .Z(n799) );
  NBUFFX2 U1816 ( .INP(di[6]), .Z(n821) );
  NBUFFX2 U1817 ( .INP(di[7]), .Z(n843) );
  NBUFFX2 U1818 ( .INP(di[16]), .Z(n1062) );
  NBUFFX2 U1819 ( .INP(di[17]), .Z(n1084) );
  NBUFFX2 U1820 ( .INP(di[18]), .Z(n1106) );
  NBUFFX2 U1821 ( .INP(di[19]), .Z(n1128) );
  NBUFFX2 U1822 ( .INP(di[20]), .Z(n1150) );
  NBUFFX2 U1823 ( .INP(di[21]), .Z(n1172) );
  NBUFFX2 U1824 ( .INP(di[22]), .Z(n1194) );
  NBUFFX2 U1825 ( .INP(di[23]), .Z(n1216) );
  NBUFFX2 U1826 ( .INP(di[24]), .Z(n1238) );
  NBUFFX2 U1827 ( .INP(di[25]), .Z(n1260) );
  NBUFFX2 U1828 ( .INP(di[26]), .Z(n1282) );
  NBUFFX2 U1829 ( .INP(di[27]), .Z(n1304) );
  NBUFFX2 U1830 ( .INP(di[28]), .Z(n1326) );
  NBUFFX2 U1831 ( .INP(di[29]), .Z(n1348) );
  NBUFFX2 U1832 ( .INP(di[30]), .Z(n1370) );
  NBUFFX2 U1833 ( .INP(di[31]), .Z(n1392) );
  NBUFFX2 U1834 ( .INP(di[8]), .Z(n886) );
  NBUFFX2 U1835 ( .INP(di[9]), .Z(n908) );
  NBUFFX2 U1836 ( .INP(di[10]), .Z(n930) );
  NBUFFX2 U1837 ( .INP(di[11]), .Z(n952) );
  NBUFFX2 U1838 ( .INP(di[12]), .Z(n974) );
  NBUFFX2 U1839 ( .INP(di[13]), .Z(n996) );
  NBUFFX2 U1840 ( .INP(di[14]), .Z(n1018) );
  NBUFFX2 U1841 ( .INP(di[15]), .Z(n1040) );
  NBUFFX2 U1842 ( .INP(di[0]), .Z(n710) );
  NBUFFX2 U1843 ( .INP(di[1]), .Z(n732) );
  NBUFFX2 U1844 ( .INP(di[2]), .Z(n754) );
  NBUFFX2 U1845 ( .INP(di[3]), .Z(n776) );
  NBUFFX2 U1846 ( .INP(di[4]), .Z(n798) );
  NBUFFX2 U1847 ( .INP(di[5]), .Z(n820) );
  NBUFFX2 U1848 ( .INP(di[6]), .Z(n842) );
  NBUFFX2 U1849 ( .INP(di[7]), .Z(n864) );
  DELLN2X2 U1850 ( .INP(n2170), .Z(n1) );
  DELLN2X2 U1851 ( .INP(n2170), .Z(n2) );
  DELLN2X2 U1852 ( .INP(n2170), .Z(n3) );
  DELLN2X2 U1853 ( .INP(n2170), .Z(n4) );
  DELLN2X2 U1854 ( .INP(n2170), .Z(n5) );
  DELLN2X2 U1855 ( .INP(n2170), .Z(n6) );
  DELLN2X2 U1856 ( .INP(n2170), .Z(n7) );
  DELLN2X2 U1857 ( .INP(n2170), .Z(n8) );
  DELLN2X2 U1858 ( .INP(n2170), .Z(n9) );
  DELLN2X2 U1859 ( .INP(n2170), .Z(n10) );
  DELLN2X2 U1860 ( .INP(n2170), .Z(n11) );
  DELLN2X2 U1861 ( .INP(n2170), .Z(n12) );
  DELLN2X2 U1862 ( .INP(n2170), .Z(n13) );
  DELLN2X2 U1863 ( .INP(n2170), .Z(n14) );
  DELLN2X2 U1864 ( .INP(n2170), .Z(n15) );
  DELLN2X2 U1865 ( .INP(n2170), .Z(n16) );
  DELLN2X2 U1866 ( .INP(n2170), .Z(n17) );
  DELLN2X2 U1867 ( .INP(n2170), .Z(n18) );
  DELLN2X2 U1868 ( .INP(n2170), .Z(n19) );
  DELLN2X2 U1869 ( .INP(n2194), .Z(n44) );
  DELLN2X2 U1870 ( .INP(n2194), .Z(n45) );
  DELLN2X2 U1871 ( .INP(n2194), .Z(n46) );
  DELLN2X2 U1872 ( .INP(n2194), .Z(n47) );
  DELLN2X2 U1873 ( .INP(n2194), .Z(n48) );
  DELLN2X2 U1874 ( .INP(n2194), .Z(n49) );
  DELLN2X2 U1875 ( .INP(n2194), .Z(n50) );
  DELLN2X2 U1876 ( .INP(n2194), .Z(n51) );
  DELLN2X2 U1877 ( .INP(n2194), .Z(n52) );
  DELLN2X2 U1878 ( .INP(n2194), .Z(n53) );
  DELLN2X2 U1879 ( .INP(n2194), .Z(n54) );
  DELLN2X2 U1880 ( .INP(n2194), .Z(n55) );
  DELLN2X2 U1881 ( .INP(n2194), .Z(n56) );
  DELLN2X2 U1882 ( .INP(n2194), .Z(n57) );
  DELLN2X2 U1883 ( .INP(n2194), .Z(n58) );
  DELLN2X2 U1884 ( .INP(n2194), .Z(n59) );
  DELLN2X2 U1885 ( .INP(n2194), .Z(n60) );
  DELLN2X2 U1886 ( .INP(n2194), .Z(n61) );
  DELLN2X2 U1887 ( .INP(n2194), .Z(n62) );
  DELLN2X2 U1888 ( .INP(n2205), .Z(n87) );
  DELLN2X2 U1889 ( .INP(n2205), .Z(n88) );
  DELLN2X2 U1890 ( .INP(n2205), .Z(n89) );
  DELLN2X2 U1891 ( .INP(n2205), .Z(n90) );
  DELLN2X2 U1892 ( .INP(n2205), .Z(n91) );
  DELLN2X2 U1893 ( .INP(n2205), .Z(n92) );
  DELLN2X2 U1894 ( .INP(n2205), .Z(n93) );
  DELLN2X2 U1895 ( .INP(n2205), .Z(n94) );
  DELLN2X2 U1896 ( .INP(n2205), .Z(n95) );
  DELLN2X2 U1897 ( .INP(n2205), .Z(n96) );
  DELLN2X2 U1898 ( .INP(n2205), .Z(n97) );
  DELLN2X2 U1899 ( .INP(n2205), .Z(n99) );
  DELLN2X2 U1900 ( .INP(n2205), .Z(n103) );
  DELLN2X2 U1901 ( .INP(n2205), .Z(n107) );
  DELLN2X2 U1902 ( .INP(n2205), .Z(n111) );
  DELLN2X2 U1903 ( .INP(n2205), .Z(n115) );
  DELLN2X2 U1904 ( .INP(n2205), .Z(n119) );
  DELLN2X2 U1905 ( .INP(n2205), .Z(n123) );
  DELLN2X2 U1906 ( .INP(n2205), .Z(n127) );
  DELLN2X2 U1907 ( .INP(n2206), .Z(n130) );
  DELLN2X2 U1908 ( .INP(n2206), .Z(n131) );
  DELLN2X2 U1909 ( .INP(n2206), .Z(n132) );
  DELLN2X2 U1910 ( .INP(n2206), .Z(n133) );
  DELLN2X2 U1911 ( .INP(n2206), .Z(n134) );
  DELLN2X2 U1912 ( .INP(n2206), .Z(n135) );
  DELLN2X2 U1913 ( .INP(n2206), .Z(n136) );
  DELLN2X2 U1914 ( .INP(n2206), .Z(n137) );
  DELLN2X2 U1915 ( .INP(n2206), .Z(n138) );
  DELLN2X2 U1916 ( .INP(n2206), .Z(n139) );
  DELLN2X2 U1917 ( .INP(n2206), .Z(n140) );
  DELLN2X2 U1918 ( .INP(n2206), .Z(n142) );
  DELLN2X2 U1919 ( .INP(n2206), .Z(n146) );
  DELLN2X2 U1920 ( .INP(n2206), .Z(n150) );
  DELLN2X2 U1921 ( .INP(n2206), .Z(n154) );
  DELLN2X2 U1922 ( .INP(n2206), .Z(n158) );
  DELLN2X2 U1923 ( .INP(n2206), .Z(n162) );
  DELLN2X2 U1924 ( .INP(n2206), .Z(n166) );
  DELLN2X2 U1925 ( .INP(n2206), .Z(n170) );
  DELLN2X2 U1926 ( .INP(n2207), .Z(n173) );
  DELLN2X2 U1927 ( .INP(n2207), .Z(n174) );
  DELLN2X2 U1928 ( .INP(n2207), .Z(n175) );
  DELLN2X2 U1929 ( .INP(n2207), .Z(n176) );
  DELLN2X2 U1930 ( .INP(n2207), .Z(n177) );
  DELLN2X2 U1931 ( .INP(n2207), .Z(n178) );
  DELLN2X2 U1932 ( .INP(n2207), .Z(n179) );
  DELLN2X2 U1933 ( .INP(n2207), .Z(n180) );
  DELLN2X2 U1934 ( .INP(n2207), .Z(n181) );
  DELLN2X2 U1935 ( .INP(n2207), .Z(n182) );
  DELLN2X2 U1936 ( .INP(n2207), .Z(n183) );
  DELLN2X2 U1937 ( .INP(n2207), .Z(n184) );
  DELLN2X2 U1938 ( .INP(n2207), .Z(n185) );
  DELLN2X2 U1939 ( .INP(n2207), .Z(n186) );
  DELLN2X2 U1940 ( .INP(n2207), .Z(n187) );
  DELLN2X2 U1941 ( .INP(n2207), .Z(n188) );
  DELLN2X2 U1942 ( .INP(n2207), .Z(n189) );
  DELLN2X2 U1943 ( .INP(n2207), .Z(n190) );
  DELLN2X2 U1944 ( .INP(n2207), .Z(n191) );
  DELLN2X2 U1945 ( .INP(n2208), .Z(n216) );
  DELLN2X2 U1946 ( .INP(n2208), .Z(n217) );
  DELLN2X2 U1947 ( .INP(n2208), .Z(n218) );
  DELLN2X2 U1948 ( .INP(n2208), .Z(n219) );
  DELLN2X2 U1949 ( .INP(n2208), .Z(n220) );
  DELLN2X2 U1950 ( .INP(n2208), .Z(n221) );
  DELLN2X2 U1951 ( .INP(n2208), .Z(n222) );
  DELLN2X2 U1952 ( .INP(n2208), .Z(n223) );
  DELLN2X2 U1953 ( .INP(n2208), .Z(n224) );
  DELLN2X2 U1954 ( .INP(n2208), .Z(n225) );
  DELLN2X2 U1955 ( .INP(n2208), .Z(n226) );
  DELLN2X2 U1956 ( .INP(n2208), .Z(n227) );
  DELLN2X2 U1957 ( .INP(n2208), .Z(n228) );
  DELLN2X2 U1958 ( .INP(n2208), .Z(n229) );
  DELLN2X2 U1959 ( .INP(n2208), .Z(n230) );
  DELLN2X2 U1960 ( .INP(n2208), .Z(n231) );
  DELLN2X2 U1961 ( .INP(n2208), .Z(n232) );
  DELLN2X2 U1962 ( .INP(n2208), .Z(n233) );
  DELLN2X2 U1963 ( .INP(n2208), .Z(n234) );
  DELLN2X2 U1964 ( .INP(n2210), .Z(n259) );
  DELLN2X2 U1965 ( .INP(n2210), .Z(n260) );
  DELLN2X2 U1966 ( .INP(n2210), .Z(n261) );
  DELLN2X2 U1967 ( .INP(n2210), .Z(n262) );
  DELLN2X2 U1968 ( .INP(n2210), .Z(n263) );
  DELLN2X2 U1969 ( .INP(n2210), .Z(n264) );
  DELLN2X2 U1970 ( .INP(n2210), .Z(n265) );
  DELLN2X2 U1971 ( .INP(n2210), .Z(n266) );
  DELLN2X2 U1972 ( .INP(n2210), .Z(n267) );
  DELLN2X2 U1973 ( .INP(n2210), .Z(n268) );
  DELLN2X2 U1974 ( .INP(n2210), .Z(n269) );
  DELLN2X2 U1975 ( .INP(n2210), .Z(n270) );
  DELLN2X2 U1976 ( .INP(n2210), .Z(n271) );
  DELLN2X2 U1977 ( .INP(n2210), .Z(n272) );
  DELLN2X2 U1978 ( .INP(n2210), .Z(n273) );
  DELLN2X2 U1979 ( .INP(n2210), .Z(n274) );
  DELLN2X2 U1980 ( .INP(n2210), .Z(n275) );
  DELLN2X2 U1981 ( .INP(n2210), .Z(n276) );
  DELLN2X2 U1982 ( .INP(n2210), .Z(n277) );
  DELLN2X2 U1983 ( .INP(n2211), .Z(n302) );
  DELLN2X2 U1984 ( .INP(n2211), .Z(n303) );
  DELLN2X2 U1985 ( .INP(n2211), .Z(n304) );
  DELLN2X2 U1986 ( .INP(n2211), .Z(n305) );
  DELLN2X2 U1987 ( .INP(n2211), .Z(n306) );
  DELLN2X2 U1988 ( .INP(n2211), .Z(n307) );
  DELLN2X2 U1989 ( .INP(n2211), .Z(n308) );
  DELLN2X2 U1990 ( .INP(n2211), .Z(n309) );
  DELLN2X2 U1991 ( .INP(n2211), .Z(n310) );
  DELLN2X2 U1992 ( .INP(n2211), .Z(n311) );
  DELLN2X2 U1993 ( .INP(n2211), .Z(n312) );
  DELLN2X2 U1994 ( .INP(n2211), .Z(n313) );
  DELLN2X2 U1995 ( .INP(n2211), .Z(n314) );
  DELLN2X2 U1996 ( .INP(n2211), .Z(n315) );
  DELLN2X2 U1997 ( .INP(n2211), .Z(n316) );
  DELLN2X2 U1998 ( .INP(n2211), .Z(n317) );
  DELLN2X2 U1999 ( .INP(n2211), .Z(n318) );
  DELLN2X2 U2000 ( .INP(n2211), .Z(n319) );
  DELLN2X2 U2001 ( .INP(n2211), .Z(n320) );
  DELLN2X2 U2002 ( .INP(n2212), .Z(n345) );
  DELLN2X2 U2003 ( .INP(n2212), .Z(n346) );
  DELLN2X2 U2004 ( .INP(n2212), .Z(n347) );
  DELLN2X2 U2005 ( .INP(n2212), .Z(n348) );
  DELLN2X2 U2006 ( .INP(n2212), .Z(n349) );
  DELLN2X2 U2007 ( .INP(n2212), .Z(n350) );
  DELLN2X2 U2008 ( .INP(n2212), .Z(n351) );
  DELLN2X2 U2009 ( .INP(n2212), .Z(n352) );
  DELLN2X2 U2010 ( .INP(n2212), .Z(n353) );
  DELLN2X2 U2011 ( .INP(n2212), .Z(n354) );
  DELLN2X2 U2012 ( .INP(n2212), .Z(n355) );
  DELLN2X2 U2013 ( .INP(n2212), .Z(n356) );
  DELLN2X2 U2014 ( .INP(n2212), .Z(n357) );
  DELLN2X2 U2015 ( .INP(n2212), .Z(n358) );
  DELLN2X2 U2016 ( .INP(n2212), .Z(n359) );
  DELLN2X2 U2017 ( .INP(n2212), .Z(n360) );
  DELLN2X2 U2018 ( .INP(n2212), .Z(n361) );
  DELLN2X2 U2019 ( .INP(n2212), .Z(n362) );
  DELLN2X2 U2020 ( .INP(n2212), .Z(n363) );
  DELLN2X2 U2021 ( .INP(n2213), .Z(n388) );
  DELLN2X2 U2022 ( .INP(n2213), .Z(n389) );
  DELLN2X2 U2023 ( .INP(n2213), .Z(n390) );
  DELLN2X2 U2024 ( .INP(n2213), .Z(n391) );
  DELLN2X2 U2025 ( .INP(n2213), .Z(n392) );
  DELLN2X2 U2026 ( .INP(n2213), .Z(n393) );
  DELLN2X2 U2027 ( .INP(n2213), .Z(n394) );
  DELLN2X2 U2028 ( .INP(n2213), .Z(n395) );
  DELLN2X2 U2029 ( .INP(n2213), .Z(n396) );
  DELLN2X2 U2030 ( .INP(n2213), .Z(n397) );
  DELLN2X2 U2031 ( .INP(n2213), .Z(n398) );
  DELLN2X2 U2032 ( .INP(n2213), .Z(n399) );
  DELLN2X2 U2033 ( .INP(n2213), .Z(n400) );
  DELLN2X2 U2034 ( .INP(n2213), .Z(n401) );
  DELLN2X2 U2035 ( .INP(n2213), .Z(n402) );
  DELLN2X2 U2036 ( .INP(n2213), .Z(n403) );
  DELLN2X2 U2037 ( .INP(n2213), .Z(n404) );
  DELLN2X2 U2038 ( .INP(n2213), .Z(n405) );
  DELLN2X2 U2039 ( .INP(n2213), .Z(n406) );
  DELLN2X2 U2040 ( .INP(n2215), .Z(n431) );
  DELLN2X2 U2041 ( .INP(n2215), .Z(n432) );
  DELLN2X2 U2042 ( .INP(n2215), .Z(n433) );
  DELLN2X2 U2043 ( .INP(n2215), .Z(n434) );
  DELLN2X2 U2044 ( .INP(n2215), .Z(n435) );
  DELLN2X2 U2045 ( .INP(n2215), .Z(n436) );
  DELLN2X2 U2046 ( .INP(n2215), .Z(n437) );
  DELLN2X2 U2047 ( .INP(n2215), .Z(n438) );
  DELLN2X2 U2048 ( .INP(n2215), .Z(n439) );
  DELLN2X2 U2049 ( .INP(n2215), .Z(n440) );
  DELLN2X2 U2050 ( .INP(n2215), .Z(n441) );
  DELLN2X2 U2051 ( .INP(n2215), .Z(n443) );
  DELLN2X2 U2052 ( .INP(n2215), .Z(n447) );
  DELLN2X2 U2053 ( .INP(n2215), .Z(n451) );
  DELLN2X2 U2054 ( .INP(n2215), .Z(n455) );
  DELLN2X2 U2055 ( .INP(n2215), .Z(n459) );
  DELLN2X2 U2056 ( .INP(n2215), .Z(n463) );
  DELLN2X2 U2057 ( .INP(n2215), .Z(n467) );
  DELLN2X2 U2058 ( .INP(n2215), .Z(n471) );
  DELLN2X2 U2059 ( .INP(n2216), .Z(n474) );
  DELLN2X2 U2060 ( .INP(n2216), .Z(n475) );
  DELLN2X2 U2061 ( .INP(n2216), .Z(n476) );
  DELLN2X2 U2062 ( .INP(n2216), .Z(n477) );
  DELLN2X2 U2063 ( .INP(n2216), .Z(n478) );
  DELLN2X2 U2064 ( .INP(n2216), .Z(n479) );
  DELLN2X2 U2065 ( .INP(n2216), .Z(n480) );
  DELLN2X2 U2066 ( .INP(n2216), .Z(n481) );
  DELLN2X2 U2067 ( .INP(n2216), .Z(n482) );
  DELLN2X2 U2068 ( .INP(n2216), .Z(n483) );
  DELLN2X2 U2069 ( .INP(n2216), .Z(n484) );
  DELLN2X2 U2070 ( .INP(n2216), .Z(n486) );
  DELLN2X2 U2071 ( .INP(n2216), .Z(n490) );
  DELLN2X2 U2072 ( .INP(n2216), .Z(n494) );
  DELLN2X2 U2073 ( .INP(n2216), .Z(n498) );
  DELLN2X2 U2074 ( .INP(n2216), .Z(n502) );
  DELLN2X2 U2075 ( .INP(n2216), .Z(n506) );
  DELLN2X2 U2076 ( .INP(n2216), .Z(n510) );
  DELLN2X2 U2077 ( .INP(n2216), .Z(n514) );
  DELLN2X2 U2078 ( .INP(n2217), .Z(n517) );
  DELLN2X2 U2079 ( .INP(n2217), .Z(n518) );
  DELLN2X2 U2080 ( .INP(n2217), .Z(n519) );
  DELLN2X2 U2081 ( .INP(n2217), .Z(n520) );
  DELLN2X2 U2082 ( .INP(n2217), .Z(n521) );
  DELLN2X2 U2083 ( .INP(n2217), .Z(n522) );
  DELLN2X2 U2084 ( .INP(n2217), .Z(n523) );
  DELLN2X2 U2085 ( .INP(n2217), .Z(n524) );
  DELLN2X2 U2086 ( .INP(n2217), .Z(n525) );
  DELLN2X2 U2087 ( .INP(n2217), .Z(n526) );
  DELLN2X2 U2088 ( .INP(n2217), .Z(n527) );
  DELLN2X2 U2089 ( .INP(n2217), .Z(n528) );
  DELLN2X2 U2090 ( .INP(n2217), .Z(n529) );
  DELLN2X2 U2091 ( .INP(n2217), .Z(n530) );
  DELLN2X2 U2092 ( .INP(n2217), .Z(n531) );
  DELLN2X2 U2093 ( .INP(n2217), .Z(n532) );
  DELLN2X2 U2094 ( .INP(n2217), .Z(n533) );
  DELLN2X2 U2095 ( .INP(n2217), .Z(n534) );
  DELLN2X2 U2096 ( .INP(n2217), .Z(n535) );
  DELLN2X2 U2097 ( .INP(n2218), .Z(n560) );
  DELLN2X2 U2098 ( .INP(n2218), .Z(n561) );
  DELLN2X2 U2099 ( .INP(n2218), .Z(n562) );
  DELLN2X2 U2100 ( .INP(n2218), .Z(n563) );
  DELLN2X2 U2101 ( .INP(n2218), .Z(n564) );
  DELLN2X2 U2102 ( .INP(n2218), .Z(n565) );
  DELLN2X2 U2103 ( .INP(n2218), .Z(n566) );
  DELLN2X2 U2104 ( .INP(n2218), .Z(n567) );
  DELLN2X2 U2105 ( .INP(n2218), .Z(n568) );
  DELLN2X2 U2106 ( .INP(n2218), .Z(n569) );
  DELLN2X2 U2107 ( .INP(n2218), .Z(n570) );
  DELLN2X2 U2108 ( .INP(n2218), .Z(n571) );
  DELLN2X2 U2109 ( .INP(n2218), .Z(n572) );
  DELLN2X2 U2110 ( .INP(n2218), .Z(n573) );
  DELLN2X2 U2111 ( .INP(n2218), .Z(n574) );
  DELLN2X2 U2112 ( .INP(n2218), .Z(n575) );
  DELLN2X2 U2113 ( .INP(n2218), .Z(n576) );
  DELLN2X2 U2114 ( .INP(n2218), .Z(n577) );
  DELLN2X2 U2115 ( .INP(n2218), .Z(n578) );
  DELLN2X2 U2116 ( .INP(n2220), .Z(n603) );
  DELLN2X2 U2117 ( .INP(n2220), .Z(n604) );
  DELLN2X2 U2118 ( .INP(n2220), .Z(n605) );
  DELLN2X2 U2119 ( .INP(n2220), .Z(n606) );
  DELLN2X2 U2120 ( .INP(n2220), .Z(n607) );
  DELLN2X2 U2121 ( .INP(n2220), .Z(n608) );
  DELLN2X2 U2122 ( .INP(n2220), .Z(n609) );
  DELLN2X2 U2123 ( .INP(n2220), .Z(n610) );
  DELLN2X2 U2124 ( .INP(n2220), .Z(n611) );
  DELLN2X2 U2125 ( .INP(n2220), .Z(n612) );
  DELLN2X2 U2126 ( .INP(n2220), .Z(n613) );
  DELLN2X2 U2127 ( .INP(n2220), .Z(n615) );
  DELLN2X2 U2128 ( .INP(n2220), .Z(n619) );
  DELLN2X2 U2129 ( .INP(n2220), .Z(n623) );
  DELLN2X2 U2130 ( .INP(n2220), .Z(n627) );
  DELLN2X2 U2131 ( .INP(n2220), .Z(n631) );
  DELLN2X2 U2132 ( .INP(n2220), .Z(n635) );
  DELLN2X2 U2133 ( .INP(n2220), .Z(n639) );
  DELLN2X2 U2134 ( .INP(n2220), .Z(n643) );
  DELLN2X2 U2135 ( .INP(n2221), .Z(n646) );
  DELLN2X2 U2136 ( .INP(n2221), .Z(n647) );
  DELLN2X2 U2137 ( .INP(n2221), .Z(n648) );
  DELLN2X2 U2138 ( .INP(n2221), .Z(n649) );
  DELLN2X2 U2139 ( .INP(n2221), .Z(n650) );
  DELLN2X2 U2140 ( .INP(n2221), .Z(n651) );
  DELLN2X2 U2141 ( .INP(n2221), .Z(n652) );
  DELLN2X2 U2142 ( .INP(n2221), .Z(n653) );
  DELLN2X2 U2143 ( .INP(n2221), .Z(n654) );
  DELLN2X2 U2144 ( .INP(n2221), .Z(n655) );
  DELLN2X2 U2145 ( .INP(n2221), .Z(n656) );
  DELLN2X2 U2146 ( .INP(n2221), .Z(n658) );
  DELLN2X2 U2147 ( .INP(n2221), .Z(n662) );
  DELLN2X2 U2148 ( .INP(n2221), .Z(n666) );
  DELLN2X2 U2149 ( .INP(n2221), .Z(n670) );
  DELLN2X2 U2150 ( .INP(n2221), .Z(n674) );
  DELLN2X2 U2151 ( .INP(n2221), .Z(n678) );
  DELLN2X2 U2152 ( .INP(n2221), .Z(n682) );
  DELLN2X2 U2153 ( .INP(n2221), .Z(n686) );
  OR4X1 U2154 ( .IN1(n2153), .IN2(n2154), .IN3(n2155), .IN4(n2156), .Q(n2203)
         );
  AO221X1 U2155 ( .IN1(n2157), .IN2(n2158), .IN3(n2159), .IN4(n2160), .IN5(
        n2161), .Q(n2156) );
  AO22X1 U2156 ( .IN1(n2162), .IN2(n2163), .IN3(n2164), .IN4(n2165), .Q(n2161)
         );
  NAND4X0 U2157 ( .IN1(n2166), .IN2(n2167), .IN3(n2168), .IN4(n2169), .QN(
        n2165) );
  OA221X1 U2158 ( .IN1(n24552), .IN2(n43), .IN3(n24560), .IN4(n86), .IN5(n2204), .Q(n2169) );
  OA22X1 U2159 ( .IN1(n24568), .IN2(n129), .IN3(n24576), .IN4(n172), .Q(n2204)
         );
  OA221X1 U2160 ( .IN1(n24520), .IN2(n215), .IN3(n24528), .IN4(n258), .IN5(
        n2209), .Q(n2168) );
  OA22X1 U2161 ( .IN1(n24536), .IN2(n301), .IN3(n24544), .IN4(n344), .Q(n2209)
         );
  OA221X1 U2162 ( .IN1(n24488), .IN2(n387), .IN3(n24496), .IN4(n430), .IN5(
        n2214), .Q(n2167) );
  OA22X1 U2163 ( .IN1(n24504), .IN2(n473), .IN3(n24512), .IN4(n516), .Q(n2214)
         );
  OA221X1 U2164 ( .IN1(n24456), .IN2(n559), .IN3(n24464), .IN4(n602), .IN5(
        n2219), .Q(n2166) );
  OA22X1 U2165 ( .IN1(n24472), .IN2(n645), .IN3(n24480), .IN4(n688), .Q(n2219)
         );
  NAND4X0 U2166 ( .IN1(n2222), .IN2(n2223), .IN3(n2224), .IN4(n2225), .QN(
        n2163) );
  OA221X1 U2167 ( .IN1(n24424), .IN2(n43), .IN3(n24432), .IN4(n86), .IN5(n2226), .Q(n2225) );
  OA22X1 U2168 ( .IN1(n24440), .IN2(n129), .IN3(n24448), .IN4(n172), .Q(n2226)
         );
  OA221X1 U2169 ( .IN1(n24392), .IN2(n215), .IN3(n24400), .IN4(n258), .IN5(
        n2227), .Q(n2224) );
  OA22X1 U2170 ( .IN1(n24408), .IN2(n301), .IN3(n24416), .IN4(n344), .Q(n2227)
         );
  OA221X1 U2171 ( .IN1(n24360), .IN2(n387), .IN3(n24368), .IN4(n430), .IN5(
        n2228), .Q(n2223) );
  OA22X1 U2172 ( .IN1(n24376), .IN2(n473), .IN3(n24384), .IN4(n516), .Q(n2228)
         );
  OA221X1 U2173 ( .IN1(n24328), .IN2(n559), .IN3(n24336), .IN4(n602), .IN5(
        n2229), .Q(n2222) );
  OA22X1 U2174 ( .IN1(n24344), .IN2(n645), .IN3(n24352), .IN4(n688), .Q(n2229)
         );
  NAND4X0 U2175 ( .IN1(n2230), .IN2(n2231), .IN3(n2232), .IN4(n2233), .QN(
        n2160) );
  OA221X1 U2176 ( .IN1(n24296), .IN2(n43), .IN3(n24304), .IN4(n86), .IN5(n2234), .Q(n2233) );
  OA22X1 U2177 ( .IN1(n24312), .IN2(n129), .IN3(n24320), .IN4(n172), .Q(n2234)
         );
  OA221X1 U2178 ( .IN1(n24264), .IN2(n215), .IN3(n24272), .IN4(n258), .IN5(
        n2235), .Q(n2232) );
  OA22X1 U2179 ( .IN1(n24280), .IN2(n301), .IN3(n24288), .IN4(n344), .Q(n2235)
         );
  OA221X1 U2180 ( .IN1(n24232), .IN2(n387), .IN3(n24240), .IN4(n430), .IN5(
        n2236), .Q(n2231) );
  OA22X1 U2181 ( .IN1(n24248), .IN2(n473), .IN3(n24256), .IN4(n516), .Q(n2236)
         );
  OA221X1 U2182 ( .IN1(n24200), .IN2(n559), .IN3(n24208), .IN4(n602), .IN5(
        n2237), .Q(n2230) );
  OA22X1 U2183 ( .IN1(n24216), .IN2(n645), .IN3(n24224), .IN4(n688), .Q(n2237)
         );
  NAND4X0 U2184 ( .IN1(n2238), .IN2(n2239), .IN3(n2240), .IN4(n2241), .QN(
        n2158) );
  OA221X1 U2185 ( .IN1(n24168), .IN2(n43), .IN3(n24176), .IN4(n86), .IN5(n2242), .Q(n2241) );
  OA22X1 U2186 ( .IN1(n24184), .IN2(n129), .IN3(n24192), .IN4(n172), .Q(n2242)
         );
  OA221X1 U2187 ( .IN1(n24136), .IN2(n215), .IN3(n24144), .IN4(n258), .IN5(
        n2243), .Q(n2240) );
  OA22X1 U2188 ( .IN1(n24152), .IN2(n301), .IN3(n24160), .IN4(n344), .Q(n2243)
         );
  OA221X1 U2189 ( .IN1(n24104), .IN2(n387), .IN3(n24112), .IN4(n430), .IN5(
        n2244), .Q(n2239) );
  OA22X1 U2190 ( .IN1(n24120), .IN2(n473), .IN3(n24128), .IN4(n516), .Q(n2244)
         );
  OA221X1 U2191 ( .IN1(n24072), .IN2(n559), .IN3(n24080), .IN4(n602), .IN5(
        n2245), .Q(n2238) );
  OA22X1 U2192 ( .IN1(n24088), .IN2(n645), .IN3(n24096), .IN4(n688), .Q(n2245)
         );
  AO221X1 U2193 ( .IN1(n2246), .IN2(n2247), .IN3(n2248), .IN4(n2249), .IN5(
        n2250), .Q(n2155) );
  AO22X1 U2194 ( .IN1(n2251), .IN2(n2252), .IN3(n2253), .IN4(n2254), .Q(n2250)
         );
  NAND4X0 U2195 ( .IN1(n2255), .IN2(n2256), .IN3(n2257), .IN4(n2258), .QN(
        n2254) );
  OA221X1 U2196 ( .IN1(n24040), .IN2(n43), .IN3(n24048), .IN4(n86), .IN5(n2259), .Q(n2258) );
  OA22X1 U2197 ( .IN1(n24056), .IN2(n129), .IN3(n24064), .IN4(n172), .Q(n2259)
         );
  OA221X1 U2198 ( .IN1(n24008), .IN2(n215), .IN3(n24016), .IN4(n258), .IN5(
        n2260), .Q(n2257) );
  OA22X1 U2199 ( .IN1(n24024), .IN2(n301), .IN3(n24032), .IN4(n344), .Q(n2260)
         );
  OA221X1 U2200 ( .IN1(n23976), .IN2(n387), .IN3(n23984), .IN4(n430), .IN5(
        n2261), .Q(n2256) );
  OA22X1 U2201 ( .IN1(n23992), .IN2(n473), .IN3(n24000), .IN4(n516), .Q(n2261)
         );
  OA221X1 U2202 ( .IN1(n23944), .IN2(n559), .IN3(n23952), .IN4(n602), .IN5(
        n2262), .Q(n2255) );
  OA22X1 U2203 ( .IN1(n23960), .IN2(n645), .IN3(n23968), .IN4(n688), .Q(n2262)
         );
  NAND4X0 U2204 ( .IN1(n2263), .IN2(n2264), .IN3(n2265), .IN4(n2266), .QN(
        n2252) );
  OA221X1 U2205 ( .IN1(n23912), .IN2(n43), .IN3(n23920), .IN4(n86), .IN5(n2267), .Q(n2266) );
  OA22X1 U2206 ( .IN1(n23928), .IN2(n129), .IN3(n23936), .IN4(n172), .Q(n2267)
         );
  OA221X1 U2207 ( .IN1(n23880), .IN2(n215), .IN3(n23888), .IN4(n258), .IN5(
        n2268), .Q(n2265) );
  OA22X1 U2208 ( .IN1(n23896), .IN2(n301), .IN3(n23904), .IN4(n344), .Q(n2268)
         );
  OA221X1 U2209 ( .IN1(n23848), .IN2(n387), .IN3(n23856), .IN4(n430), .IN5(
        n2269), .Q(n2264) );
  OA22X1 U2210 ( .IN1(n23864), .IN2(n473), .IN3(n23872), .IN4(n516), .Q(n2269)
         );
  OA221X1 U2211 ( .IN1(n23816), .IN2(n559), .IN3(n23824), .IN4(n602), .IN5(
        n2270), .Q(n2263) );
  OA22X1 U2212 ( .IN1(n23832), .IN2(n645), .IN3(n23840), .IN4(n688), .Q(n2270)
         );
  NAND4X0 U2213 ( .IN1(n2271), .IN2(n2272), .IN3(n2273), .IN4(n2274), .QN(
        n2249) );
  OA221X1 U2214 ( .IN1(n23784), .IN2(n43), .IN3(n23792), .IN4(n86), .IN5(n2275), .Q(n2274) );
  OA22X1 U2215 ( .IN1(n23800), .IN2(n129), .IN3(n23808), .IN4(n172), .Q(n2275)
         );
  OA221X1 U2216 ( .IN1(n23752), .IN2(n215), .IN3(n23760), .IN4(n258), .IN5(
        n2276), .Q(n2273) );
  OA22X1 U2217 ( .IN1(n23768), .IN2(n301), .IN3(n23776), .IN4(n344), .Q(n2276)
         );
  OA221X1 U2218 ( .IN1(n23720), .IN2(n387), .IN3(n23728), .IN4(n430), .IN5(
        n2277), .Q(n2272) );
  OA22X1 U2219 ( .IN1(n23736), .IN2(n473), .IN3(n23744), .IN4(n516), .Q(n2277)
         );
  OA221X1 U2220 ( .IN1(n23688), .IN2(n559), .IN3(n23696), .IN4(n602), .IN5(
        n2278), .Q(n2271) );
  OA22X1 U2221 ( .IN1(n23704), .IN2(n645), .IN3(n23712), .IN4(n688), .Q(n2278)
         );
  NAND4X0 U2222 ( .IN1(n2279), .IN2(n2280), .IN3(n2281), .IN4(n2282), .QN(
        n2247) );
  OA221X1 U2223 ( .IN1(n23656), .IN2(n43), .IN3(n23664), .IN4(n86), .IN5(n2283), .Q(n2282) );
  OA22X1 U2224 ( .IN1(n23672), .IN2(n129), .IN3(n23680), .IN4(n172), .Q(n2283)
         );
  OA221X1 U2225 ( .IN1(n23624), .IN2(n215), .IN3(n23632), .IN4(n258), .IN5(
        n2284), .Q(n2281) );
  OA22X1 U2226 ( .IN1(n23640), .IN2(n301), .IN3(n23648), .IN4(n344), .Q(n2284)
         );
  OA221X1 U2227 ( .IN1(n23592), .IN2(n387), .IN3(n23600), .IN4(n430), .IN5(
        n2285), .Q(n2280) );
  OA22X1 U2228 ( .IN1(n23608), .IN2(n473), .IN3(n23616), .IN4(n516), .Q(n2285)
         );
  OA221X1 U2229 ( .IN1(n23560), .IN2(n559), .IN3(n23568), .IN4(n602), .IN5(
        n2286), .Q(n2279) );
  OA22X1 U2230 ( .IN1(n23576), .IN2(n645), .IN3(n23584), .IN4(n688), .Q(n2286)
         );
  AO221X1 U2231 ( .IN1(n2287), .IN2(n2288), .IN3(n2289), .IN4(n2290), .IN5(
        n2291), .Q(n2154) );
  AO22X1 U2232 ( .IN1(n2292), .IN2(n2293), .IN3(n2294), .IN4(n2295), .Q(n2291)
         );
  NAND4X0 U2233 ( .IN1(n2296), .IN2(n2297), .IN3(n2298), .IN4(n2299), .QN(
        n2295) );
  OA221X1 U2234 ( .IN1(n25576), .IN2(n42), .IN3(n25584), .IN4(n85), .IN5(n2300), .Q(n2299) );
  OA22X1 U2235 ( .IN1(n25592), .IN2(n128), .IN3(n25600), .IN4(n171), .Q(n2300)
         );
  OA221X1 U2236 ( .IN1(n25544), .IN2(n214), .IN3(n25552), .IN4(n257), .IN5(
        n2301), .Q(n2298) );
  OA22X1 U2237 ( .IN1(n25560), .IN2(n300), .IN3(n25568), .IN4(n343), .Q(n2301)
         );
  OA221X1 U2238 ( .IN1(n25512), .IN2(n386), .IN3(n25520), .IN4(n429), .IN5(
        n2302), .Q(n2297) );
  OA22X1 U2239 ( .IN1(n25528), .IN2(n472), .IN3(n25536), .IN4(n515), .Q(n2302)
         );
  OA221X1 U2240 ( .IN1(n25480), .IN2(n558), .IN3(n25488), .IN4(n601), .IN5(
        n2303), .Q(n2296) );
  OA22X1 U2241 ( .IN1(n25496), .IN2(n644), .IN3(n25504), .IN4(n687), .Q(n2303)
         );
  NAND4X0 U2242 ( .IN1(n2304), .IN2(n2305), .IN3(n2306), .IN4(n2307), .QN(
        n2293) );
  OA221X1 U2243 ( .IN1(n25448), .IN2(n42), .IN3(n25456), .IN4(n85), .IN5(n2308), .Q(n2307) );
  OA22X1 U2244 ( .IN1(n25464), .IN2(n128), .IN3(n25472), .IN4(n171), .Q(n2308)
         );
  OA221X1 U2245 ( .IN1(n25416), .IN2(n214), .IN3(n25424), .IN4(n257), .IN5(
        n2309), .Q(n2306) );
  OA22X1 U2246 ( .IN1(n25432), .IN2(n300), .IN3(n25440), .IN4(n343), .Q(n2309)
         );
  OA221X1 U2247 ( .IN1(n25384), .IN2(n386), .IN3(n25392), .IN4(n429), .IN5(
        n2310), .Q(n2305) );
  OA22X1 U2248 ( .IN1(n25400), .IN2(n472), .IN3(n25408), .IN4(n515), .Q(n2310)
         );
  OA221X1 U2249 ( .IN1(n25352), .IN2(n558), .IN3(n25360), .IN4(n601), .IN5(
        n2311), .Q(n2304) );
  OA22X1 U2250 ( .IN1(n25368), .IN2(n644), .IN3(n25376), .IN4(n687), .Q(n2311)
         );
  NAND4X0 U2251 ( .IN1(n2312), .IN2(n2313), .IN3(n2314), .IN4(n2315), .QN(
        n2290) );
  OA221X1 U2252 ( .IN1(n25320), .IN2(n42), .IN3(n25328), .IN4(n85), .IN5(n2316), .Q(n2315) );
  OA22X1 U2253 ( .IN1(n25336), .IN2(n128), .IN3(n25344), .IN4(n171), .Q(n2316)
         );
  OA221X1 U2254 ( .IN1(n25288), .IN2(n214), .IN3(n25296), .IN4(n257), .IN5(
        n2317), .Q(n2314) );
  OA22X1 U2255 ( .IN1(n25304), .IN2(n300), .IN3(n25312), .IN4(n343), .Q(n2317)
         );
  OA221X1 U2256 ( .IN1(n25256), .IN2(n386), .IN3(n25264), .IN4(n429), .IN5(
        n2318), .Q(n2313) );
  OA22X1 U2257 ( .IN1(n25272), .IN2(n472), .IN3(n25280), .IN4(n515), .Q(n2318)
         );
  OA221X1 U2258 ( .IN1(n25224), .IN2(n558), .IN3(n25232), .IN4(n601), .IN5(
        n2319), .Q(n2312) );
  OA22X1 U2259 ( .IN1(n25240), .IN2(n644), .IN3(n25248), .IN4(n687), .Q(n2319)
         );
  NAND4X0 U2260 ( .IN1(n2320), .IN2(n2321), .IN3(n2322), .IN4(n2323), .QN(
        n2288) );
  OA221X1 U2261 ( .IN1(n25192), .IN2(n42), .IN3(n25200), .IN4(n85), .IN5(n2324), .Q(n2323) );
  OA22X1 U2262 ( .IN1(n25208), .IN2(n128), .IN3(n25216), .IN4(n171), .Q(n2324)
         );
  OA221X1 U2263 ( .IN1(n25160), .IN2(n214), .IN3(n25168), .IN4(n257), .IN5(
        n2325), .Q(n2322) );
  OA22X1 U2264 ( .IN1(n25176), .IN2(n300), .IN3(n25184), .IN4(n343), .Q(n2325)
         );
  OA221X1 U2265 ( .IN1(n25128), .IN2(n386), .IN3(n25136), .IN4(n429), .IN5(
        n2326), .Q(n2321) );
  OA22X1 U2266 ( .IN1(n25144), .IN2(n472), .IN3(n25152), .IN4(n515), .Q(n2326)
         );
  OA221X1 U2267 ( .IN1(n25096), .IN2(n558), .IN3(n25104), .IN4(n601), .IN5(
        n2327), .Q(n2320) );
  OA22X1 U2268 ( .IN1(n25112), .IN2(n644), .IN3(n25120), .IN4(n687), .Q(n2327)
         );
  AO221X1 U2269 ( .IN1(n2328), .IN2(n2329), .IN3(n2330), .IN4(n2331), .IN5(
        n2332), .Q(n2153) );
  AO22X1 U2270 ( .IN1(n2333), .IN2(n2334), .IN3(n2335), .IN4(n2336), .Q(n2332)
         );
  NAND4X0 U2271 ( .IN1(n2337), .IN2(n2338), .IN3(n2339), .IN4(n2340), .QN(
        n2336) );
  OA221X1 U2272 ( .IN1(n25064), .IN2(n42), .IN3(n25072), .IN4(n85), .IN5(n2341), .Q(n2340) );
  OA22X1 U2273 ( .IN1(n25080), .IN2(n128), .IN3(n25088), .IN4(n171), .Q(n2341)
         );
  OA221X1 U2274 ( .IN1(n25032), .IN2(n214), .IN3(n25040), .IN4(n257), .IN5(
        n2342), .Q(n2339) );
  OA22X1 U2275 ( .IN1(n25048), .IN2(n300), .IN3(n25056), .IN4(n343), .Q(n2342)
         );
  OA221X1 U2276 ( .IN1(n25000), .IN2(n386), .IN3(n25008), .IN4(n429), .IN5(
        n2343), .Q(n2338) );
  OA22X1 U2277 ( .IN1(n25016), .IN2(n472), .IN3(n25024), .IN4(n515), .Q(n2343)
         );
  OA221X1 U2278 ( .IN1(n24968), .IN2(n558), .IN3(n24976), .IN4(n601), .IN5(
        n2344), .Q(n2337) );
  OA22X1 U2279 ( .IN1(n24984), .IN2(n644), .IN3(n24992), .IN4(n687), .Q(n2344)
         );
  NAND4X0 U2280 ( .IN1(n2345), .IN2(n2346), .IN3(n2347), .IN4(n2348), .QN(
        n2334) );
  OA221X1 U2281 ( .IN1(n24936), .IN2(n42), .IN3(n24944), .IN4(n85), .IN5(n2349), .Q(n2348) );
  OA22X1 U2282 ( .IN1(n24952), .IN2(n128), .IN3(n24960), .IN4(n171), .Q(n2349)
         );
  OA221X1 U2283 ( .IN1(n24904), .IN2(n214), .IN3(n24912), .IN4(n257), .IN5(
        n2350), .Q(n2347) );
  OA22X1 U2284 ( .IN1(n24920), .IN2(n300), .IN3(n24928), .IN4(n343), .Q(n2350)
         );
  OA221X1 U2285 ( .IN1(n24872), .IN2(n386), .IN3(n24880), .IN4(n429), .IN5(
        n2351), .Q(n2346) );
  OA22X1 U2286 ( .IN1(n24888), .IN2(n472), .IN3(n24896), .IN4(n515), .Q(n2351)
         );
  OA221X1 U2287 ( .IN1(n24840), .IN2(n558), .IN3(n24848), .IN4(n601), .IN5(
        n2352), .Q(n2345) );
  OA22X1 U2288 ( .IN1(n24856), .IN2(n644), .IN3(n24864), .IN4(n687), .Q(n2352)
         );
  NAND4X0 U2289 ( .IN1(n2353), .IN2(n2354), .IN3(n2355), .IN4(n2356), .QN(
        n2331) );
  OA221X1 U2290 ( .IN1(n24808), .IN2(n42), .IN3(n24816), .IN4(n85), .IN5(n2357), .Q(n2356) );
  OA22X1 U2291 ( .IN1(n24824), .IN2(n128), .IN3(n24832), .IN4(n171), .Q(n2357)
         );
  OA221X1 U2292 ( .IN1(n24776), .IN2(n214), .IN3(n24784), .IN4(n257), .IN5(
        n2358), .Q(n2355) );
  OA22X1 U2293 ( .IN1(n24792), .IN2(n300), .IN3(n24800), .IN4(n343), .Q(n2358)
         );
  OA221X1 U2294 ( .IN1(n24744), .IN2(n386), .IN3(n24752), .IN4(n429), .IN5(
        n2359), .Q(n2354) );
  OA22X1 U2295 ( .IN1(n24760), .IN2(n472), .IN3(n24768), .IN4(n515), .Q(n2359)
         );
  OA221X1 U2296 ( .IN1(n24712), .IN2(n558), .IN3(n24720), .IN4(n601), .IN5(
        n2360), .Q(n2353) );
  OA22X1 U2297 ( .IN1(n24728), .IN2(n644), .IN3(n24736), .IN4(n687), .Q(n2360)
         );
  NAND4X0 U2298 ( .IN1(n2361), .IN2(n2362), .IN3(n2363), .IN4(n2364), .QN(
        n2329) );
  OA221X1 U2299 ( .IN1(n24680), .IN2(n42), .IN3(n24688), .IN4(n85), .IN5(n2365), .Q(n2364) );
  OA22X1 U2300 ( .IN1(n24696), .IN2(n128), .IN3(n24704), .IN4(n171), .Q(n2365)
         );
  OA221X1 U2301 ( .IN1(n24648), .IN2(n214), .IN3(n24656), .IN4(n257), .IN5(
        n2366), .Q(n2363) );
  OA22X1 U2302 ( .IN1(n24664), .IN2(n300), .IN3(n24672), .IN4(n343), .Q(n2366)
         );
  OA221X1 U2303 ( .IN1(n24616), .IN2(n386), .IN3(n24624), .IN4(n429), .IN5(
        n2367), .Q(n2362) );
  OA22X1 U2304 ( .IN1(n24632), .IN2(n472), .IN3(n24640), .IN4(n515), .Q(n2367)
         );
  OA221X1 U2305 ( .IN1(n24584), .IN2(n558), .IN3(n24592), .IN4(n601), .IN5(
        n2368), .Q(n2361) );
  OA22X1 U2306 ( .IN1(n24600), .IN2(n644), .IN3(n24608), .IN4(n687), .Q(n2368)
         );
  OR4X1 U2307 ( .IN1(n2369), .IN2(n2370), .IN3(n2371), .IN4(n2372), .Q(n2202)
         );
  AO221X1 U2308 ( .IN1(n2157), .IN2(n2373), .IN3(n2159), .IN4(n2374), .IN5(
        n2375), .Q(n2372) );
  AO22X1 U2309 ( .IN1(n2162), .IN2(n2376), .IN3(n2164), .IN4(n2377), .Q(n2375)
         );
  NAND4X0 U2310 ( .IN1(n2378), .IN2(n2379), .IN3(n2380), .IN4(n2381), .QN(
        n2377) );
  OA221X1 U2311 ( .IN1(n24551), .IN2(n42), .IN3(n24559), .IN4(n85), .IN5(n2382), .Q(n2381) );
  OA22X1 U2312 ( .IN1(n24567), .IN2(n128), .IN3(n24575), .IN4(n171), .Q(n2382)
         );
  OA221X1 U2313 ( .IN1(n24519), .IN2(n214), .IN3(n24527), .IN4(n257), .IN5(
        n2383), .Q(n2380) );
  OA22X1 U2314 ( .IN1(n24535), .IN2(n300), .IN3(n24543), .IN4(n343), .Q(n2383)
         );
  OA221X1 U2315 ( .IN1(n24487), .IN2(n386), .IN3(n24495), .IN4(n429), .IN5(
        n2384), .Q(n2379) );
  OA22X1 U2316 ( .IN1(n24503), .IN2(n472), .IN3(n24511), .IN4(n515), .Q(n2384)
         );
  OA221X1 U2317 ( .IN1(n24455), .IN2(n558), .IN3(n24463), .IN4(n601), .IN5(
        n2385), .Q(n2378) );
  OA22X1 U2318 ( .IN1(n24471), .IN2(n644), .IN3(n24479), .IN4(n687), .Q(n2385)
         );
  NAND4X0 U2319 ( .IN1(n2386), .IN2(n2387), .IN3(n2388), .IN4(n2389), .QN(
        n2376) );
  OA221X1 U2320 ( .IN1(n24423), .IN2(n42), .IN3(n24431), .IN4(n85), .IN5(n2390), .Q(n2389) );
  OA22X1 U2321 ( .IN1(n24439), .IN2(n128), .IN3(n24447), .IN4(n171), .Q(n2390)
         );
  OA221X1 U2322 ( .IN1(n24391), .IN2(n214), .IN3(n24399), .IN4(n257), .IN5(
        n2391), .Q(n2388) );
  OA22X1 U2323 ( .IN1(n24407), .IN2(n300), .IN3(n24415), .IN4(n343), .Q(n2391)
         );
  OA221X1 U2324 ( .IN1(n24359), .IN2(n386), .IN3(n24367), .IN4(n429), .IN5(
        n2392), .Q(n2387) );
  OA22X1 U2325 ( .IN1(n24375), .IN2(n472), .IN3(n24383), .IN4(n515), .Q(n2392)
         );
  OA221X1 U2326 ( .IN1(n24327), .IN2(n558), .IN3(n24335), .IN4(n601), .IN5(
        n2393), .Q(n2386) );
  OA22X1 U2327 ( .IN1(n24343), .IN2(n644), .IN3(n24351), .IN4(n687), .Q(n2393)
         );
  NAND4X0 U2328 ( .IN1(n2394), .IN2(n2395), .IN3(n2396), .IN4(n2397), .QN(
        n2374) );
  OA221X1 U2329 ( .IN1(n24295), .IN2(n42), .IN3(n24303), .IN4(n85), .IN5(n2398), .Q(n2397) );
  OA22X1 U2330 ( .IN1(n24311), .IN2(n128), .IN3(n24319), .IN4(n171), .Q(n2398)
         );
  OA221X1 U2331 ( .IN1(n24263), .IN2(n214), .IN3(n24271), .IN4(n257), .IN5(
        n2399), .Q(n2396) );
  OA22X1 U2332 ( .IN1(n24279), .IN2(n300), .IN3(n24287), .IN4(n343), .Q(n2399)
         );
  OA221X1 U2333 ( .IN1(n24231), .IN2(n386), .IN3(n24239), .IN4(n429), .IN5(
        n2400), .Q(n2395) );
  OA22X1 U2334 ( .IN1(n24247), .IN2(n472), .IN3(n24255), .IN4(n515), .Q(n2400)
         );
  OA221X1 U2335 ( .IN1(n24199), .IN2(n558), .IN3(n24207), .IN4(n601), .IN5(
        n2401), .Q(n2394) );
  OA22X1 U2336 ( .IN1(n24215), .IN2(n644), .IN3(n24223), .IN4(n687), .Q(n2401)
         );
  NAND4X0 U2337 ( .IN1(n2402), .IN2(n2403), .IN3(n2404), .IN4(n2405), .QN(
        n2373) );
  OA221X1 U2338 ( .IN1(n24167), .IN2(n42), .IN3(n24175), .IN4(n85), .IN5(n2406), .Q(n2405) );
  OA22X1 U2339 ( .IN1(n24183), .IN2(n128), .IN3(n24191), .IN4(n171), .Q(n2406)
         );
  OA221X1 U2340 ( .IN1(n24135), .IN2(n214), .IN3(n24143), .IN4(n257), .IN5(
        n2407), .Q(n2404) );
  OA22X1 U2341 ( .IN1(n24151), .IN2(n300), .IN3(n24159), .IN4(n343), .Q(n2407)
         );
  OA221X1 U2342 ( .IN1(n24103), .IN2(n386), .IN3(n24111), .IN4(n429), .IN5(
        n2408), .Q(n2403) );
  OA22X1 U2343 ( .IN1(n24119), .IN2(n472), .IN3(n24127), .IN4(n515), .Q(n2408)
         );
  OA221X1 U2344 ( .IN1(n24071), .IN2(n558), .IN3(n24079), .IN4(n601), .IN5(
        n2409), .Q(n2402) );
  OA22X1 U2345 ( .IN1(n24087), .IN2(n644), .IN3(n24095), .IN4(n687), .Q(n2409)
         );
  AO221X1 U2346 ( .IN1(n2246), .IN2(n2410), .IN3(n2248), .IN4(n2411), .IN5(
        n2412), .Q(n2371) );
  AO22X1 U2347 ( .IN1(n2251), .IN2(n2413), .IN3(n2253), .IN4(n2414), .Q(n2412)
         );
  NAND4X0 U2348 ( .IN1(n2415), .IN2(n2416), .IN3(n2417), .IN4(n2418), .QN(
        n2414) );
  OA221X1 U2349 ( .IN1(n24039), .IN2(n41), .IN3(n24047), .IN4(n84), .IN5(n2419), .Q(n2418) );
  OA22X1 U2350 ( .IN1(n24055), .IN2(n127), .IN3(n24063), .IN4(n170), .Q(n2419)
         );
  OA221X1 U2351 ( .IN1(n24007), .IN2(n213), .IN3(n24015), .IN4(n256), .IN5(
        n2420), .Q(n2417) );
  OA22X1 U2352 ( .IN1(n24023), .IN2(n299), .IN3(n24031), .IN4(n342), .Q(n2420)
         );
  OA221X1 U2353 ( .IN1(n23975), .IN2(n385), .IN3(n23983), .IN4(n428), .IN5(
        n2421), .Q(n2416) );
  OA22X1 U2354 ( .IN1(n23991), .IN2(n471), .IN3(n23999), .IN4(n514), .Q(n2421)
         );
  OA221X1 U2355 ( .IN1(n23943), .IN2(n557), .IN3(n23951), .IN4(n600), .IN5(
        n2422), .Q(n2415) );
  OA22X1 U2356 ( .IN1(n23959), .IN2(n643), .IN3(n23967), .IN4(n686), .Q(n2422)
         );
  NAND4X0 U2357 ( .IN1(n2423), .IN2(n2424), .IN3(n2425), .IN4(n2426), .QN(
        n2413) );
  OA221X1 U2358 ( .IN1(n23911), .IN2(n41), .IN3(n23919), .IN4(n84), .IN5(n2427), .Q(n2426) );
  OA22X1 U2359 ( .IN1(n23927), .IN2(n127), .IN3(n23935), .IN4(n170), .Q(n2427)
         );
  OA221X1 U2360 ( .IN1(n23879), .IN2(n213), .IN3(n23887), .IN4(n256), .IN5(
        n2428), .Q(n2425) );
  OA22X1 U2361 ( .IN1(n23895), .IN2(n299), .IN3(n23903), .IN4(n342), .Q(n2428)
         );
  OA221X1 U2362 ( .IN1(n23847), .IN2(n385), .IN3(n23855), .IN4(n428), .IN5(
        n2429), .Q(n2424) );
  OA22X1 U2363 ( .IN1(n23863), .IN2(n471), .IN3(n23871), .IN4(n514), .Q(n2429)
         );
  OA221X1 U2364 ( .IN1(n23815), .IN2(n557), .IN3(n23823), .IN4(n600), .IN5(
        n2430), .Q(n2423) );
  OA22X1 U2365 ( .IN1(n23831), .IN2(n643), .IN3(n23839), .IN4(n686), .Q(n2430)
         );
  NAND4X0 U2366 ( .IN1(n2431), .IN2(n2432), .IN3(n2433), .IN4(n2434), .QN(
        n2411) );
  OA221X1 U2367 ( .IN1(n23783), .IN2(n41), .IN3(n23791), .IN4(n84), .IN5(n2435), .Q(n2434) );
  OA22X1 U2368 ( .IN1(n23799), .IN2(n127), .IN3(n23807), .IN4(n170), .Q(n2435)
         );
  OA221X1 U2369 ( .IN1(n23751), .IN2(n213), .IN3(n23759), .IN4(n256), .IN5(
        n2436), .Q(n2433) );
  OA22X1 U2370 ( .IN1(n23767), .IN2(n299), .IN3(n23775), .IN4(n342), .Q(n2436)
         );
  OA221X1 U2371 ( .IN1(n23719), .IN2(n385), .IN3(n23727), .IN4(n428), .IN5(
        n2437), .Q(n2432) );
  OA22X1 U2372 ( .IN1(n23735), .IN2(n471), .IN3(n23743), .IN4(n514), .Q(n2437)
         );
  OA221X1 U2373 ( .IN1(n23687), .IN2(n557), .IN3(n23695), .IN4(n600), .IN5(
        n2438), .Q(n2431) );
  OA22X1 U2374 ( .IN1(n23703), .IN2(n643), .IN3(n23711), .IN4(n686), .Q(n2438)
         );
  NAND4X0 U2375 ( .IN1(n2439), .IN2(n2440), .IN3(n2441), .IN4(n2442), .QN(
        n2410) );
  OA221X1 U2376 ( .IN1(n23655), .IN2(n41), .IN3(n23663), .IN4(n84), .IN5(n2443), .Q(n2442) );
  OA22X1 U2377 ( .IN1(n23671), .IN2(n127), .IN3(n23679), .IN4(n170), .Q(n2443)
         );
  OA221X1 U2378 ( .IN1(n23623), .IN2(n213), .IN3(n23631), .IN4(n256), .IN5(
        n2444), .Q(n2441) );
  OA22X1 U2379 ( .IN1(n23639), .IN2(n299), .IN3(n23647), .IN4(n342), .Q(n2444)
         );
  OA221X1 U2380 ( .IN1(n23591), .IN2(n385), .IN3(n23599), .IN4(n428), .IN5(
        n2445), .Q(n2440) );
  OA22X1 U2381 ( .IN1(n23607), .IN2(n471), .IN3(n23615), .IN4(n514), .Q(n2445)
         );
  OA221X1 U2382 ( .IN1(n23559), .IN2(n557), .IN3(n23567), .IN4(n600), .IN5(
        n2446), .Q(n2439) );
  OA22X1 U2383 ( .IN1(n23575), .IN2(n643), .IN3(n23583), .IN4(n686), .Q(n2446)
         );
  AO221X1 U2384 ( .IN1(n2287), .IN2(n2447), .IN3(n2289), .IN4(n2448), .IN5(
        n2449), .Q(n2370) );
  AO22X1 U2385 ( .IN1(n2292), .IN2(n2450), .IN3(n2294), .IN4(n2451), .Q(n2449)
         );
  NAND4X0 U2386 ( .IN1(n2452), .IN2(n2453), .IN3(n2454), .IN4(n2455), .QN(
        n2451) );
  OA221X1 U2387 ( .IN1(n25575), .IN2(n41), .IN3(n25583), .IN4(n84), .IN5(n2456), .Q(n2455) );
  OA22X1 U2388 ( .IN1(n25591), .IN2(n127), .IN3(n25599), .IN4(n170), .Q(n2456)
         );
  OA221X1 U2389 ( .IN1(n25543), .IN2(n213), .IN3(n25551), .IN4(n256), .IN5(
        n2457), .Q(n2454) );
  OA22X1 U2390 ( .IN1(n25559), .IN2(n299), .IN3(n25567), .IN4(n342), .Q(n2457)
         );
  OA221X1 U2391 ( .IN1(n25511), .IN2(n385), .IN3(n25519), .IN4(n428), .IN5(
        n2458), .Q(n2453) );
  OA22X1 U2392 ( .IN1(n25527), .IN2(n471), .IN3(n25535), .IN4(n514), .Q(n2458)
         );
  OA221X1 U2393 ( .IN1(n25479), .IN2(n557), .IN3(n25487), .IN4(n600), .IN5(
        n2459), .Q(n2452) );
  OA22X1 U2394 ( .IN1(n25495), .IN2(n643), .IN3(n25503), .IN4(n686), .Q(n2459)
         );
  NAND4X0 U2395 ( .IN1(n2460), .IN2(n2461), .IN3(n2462), .IN4(n2463), .QN(
        n2450) );
  OA221X1 U2396 ( .IN1(n25447), .IN2(n41), .IN3(n25455), .IN4(n84), .IN5(n2464), .Q(n2463) );
  OA22X1 U2397 ( .IN1(n25463), .IN2(n127), .IN3(n25471), .IN4(n170), .Q(n2464)
         );
  OA221X1 U2398 ( .IN1(n25415), .IN2(n213), .IN3(n25423), .IN4(n256), .IN5(
        n2465), .Q(n2462) );
  OA22X1 U2399 ( .IN1(n25431), .IN2(n299), .IN3(n25439), .IN4(n342), .Q(n2465)
         );
  OA221X1 U2400 ( .IN1(n25383), .IN2(n385), .IN3(n25391), .IN4(n428), .IN5(
        n2466), .Q(n2461) );
  OA22X1 U2401 ( .IN1(n25399), .IN2(n471), .IN3(n25407), .IN4(n514), .Q(n2466)
         );
  OA221X1 U2402 ( .IN1(n25351), .IN2(n557), .IN3(n25359), .IN4(n600), .IN5(
        n2467), .Q(n2460) );
  OA22X1 U2403 ( .IN1(n25367), .IN2(n643), .IN3(n25375), .IN4(n686), .Q(n2467)
         );
  NAND4X0 U2404 ( .IN1(n2468), .IN2(n2469), .IN3(n2470), .IN4(n2471), .QN(
        n2448) );
  OA221X1 U2405 ( .IN1(n25319), .IN2(n41), .IN3(n25327), .IN4(n84), .IN5(n2472), .Q(n2471) );
  OA22X1 U2406 ( .IN1(n25335), .IN2(n127), .IN3(n25343), .IN4(n170), .Q(n2472)
         );
  OA221X1 U2407 ( .IN1(n25287), .IN2(n213), .IN3(n25295), .IN4(n256), .IN5(
        n2473), .Q(n2470) );
  OA22X1 U2408 ( .IN1(n25303), .IN2(n299), .IN3(n25311), .IN4(n342), .Q(n2473)
         );
  OA221X1 U2409 ( .IN1(n25255), .IN2(n385), .IN3(n25263), .IN4(n428), .IN5(
        n2474), .Q(n2469) );
  OA22X1 U2410 ( .IN1(n25271), .IN2(n471), .IN3(n25279), .IN4(n514), .Q(n2474)
         );
  OA221X1 U2411 ( .IN1(n25223), .IN2(n557), .IN3(n25231), .IN4(n600), .IN5(
        n2475), .Q(n2468) );
  OA22X1 U2412 ( .IN1(n25239), .IN2(n643), .IN3(n25247), .IN4(n686), .Q(n2475)
         );
  NAND4X0 U2413 ( .IN1(n2476), .IN2(n2477), .IN3(n2478), .IN4(n2479), .QN(
        n2447) );
  OA221X1 U2414 ( .IN1(n25191), .IN2(n41), .IN3(n25199), .IN4(n84), .IN5(n2480), .Q(n2479) );
  OA22X1 U2415 ( .IN1(n25207), .IN2(n127), .IN3(n25215), .IN4(n170), .Q(n2480)
         );
  OA221X1 U2416 ( .IN1(n25159), .IN2(n213), .IN3(n25167), .IN4(n256), .IN5(
        n2481), .Q(n2478) );
  OA22X1 U2417 ( .IN1(n25175), .IN2(n299), .IN3(n25183), .IN4(n342), .Q(n2481)
         );
  OA221X1 U2418 ( .IN1(n25127), .IN2(n385), .IN3(n25135), .IN4(n428), .IN5(
        n2482), .Q(n2477) );
  OA22X1 U2419 ( .IN1(n25143), .IN2(n471), .IN3(n25151), .IN4(n514), .Q(n2482)
         );
  OA221X1 U2420 ( .IN1(n25095), .IN2(n557), .IN3(n25103), .IN4(n600), .IN5(
        n2483), .Q(n2476) );
  OA22X1 U2421 ( .IN1(n25111), .IN2(n643), .IN3(n25119), .IN4(n686), .Q(n2483)
         );
  AO221X1 U2422 ( .IN1(n2328), .IN2(n2484), .IN3(n2330), .IN4(n2485), .IN5(
        n2486), .Q(n2369) );
  AO22X1 U2423 ( .IN1(n2333), .IN2(n2487), .IN3(n2335), .IN4(n2488), .Q(n2486)
         );
  NAND4X0 U2424 ( .IN1(n2489), .IN2(n2490), .IN3(n2491), .IN4(n2492), .QN(
        n2488) );
  OA221X1 U2425 ( .IN1(n25063), .IN2(n41), .IN3(n25071), .IN4(n84), .IN5(n2493), .Q(n2492) );
  OA22X1 U2426 ( .IN1(n25079), .IN2(n127), .IN3(n25087), .IN4(n170), .Q(n2493)
         );
  OA221X1 U2427 ( .IN1(n25031), .IN2(n213), .IN3(n25039), .IN4(n256), .IN5(
        n2494), .Q(n2491) );
  OA22X1 U2428 ( .IN1(n25047), .IN2(n299), .IN3(n25055), .IN4(n342), .Q(n2494)
         );
  OA221X1 U2429 ( .IN1(n24999), .IN2(n385), .IN3(n25007), .IN4(n428), .IN5(
        n2495), .Q(n2490) );
  OA22X1 U2430 ( .IN1(n25015), .IN2(n471), .IN3(n25023), .IN4(n514), .Q(n2495)
         );
  OA221X1 U2431 ( .IN1(n24967), .IN2(n557), .IN3(n24975), .IN4(n600), .IN5(
        n2496), .Q(n2489) );
  OA22X1 U2432 ( .IN1(n24983), .IN2(n643), .IN3(n24991), .IN4(n686), .Q(n2496)
         );
  NAND4X0 U2433 ( .IN1(n2497), .IN2(n2498), .IN3(n2499), .IN4(n2500), .QN(
        n2487) );
  OA221X1 U2434 ( .IN1(n24935), .IN2(n41), .IN3(n24943), .IN4(n84), .IN5(n2501), .Q(n2500) );
  OA22X1 U2435 ( .IN1(n24951), .IN2(n127), .IN3(n24959), .IN4(n170), .Q(n2501)
         );
  OA221X1 U2436 ( .IN1(n24903), .IN2(n213), .IN3(n24911), .IN4(n256), .IN5(
        n2502), .Q(n2499) );
  OA22X1 U2437 ( .IN1(n24919), .IN2(n299), .IN3(n24927), .IN4(n342), .Q(n2502)
         );
  OA221X1 U2438 ( .IN1(n24871), .IN2(n385), .IN3(n24879), .IN4(n428), .IN5(
        n2503), .Q(n2498) );
  OA22X1 U2439 ( .IN1(n24887), .IN2(n471), .IN3(n24895), .IN4(n514), .Q(n2503)
         );
  OA221X1 U2440 ( .IN1(n24839), .IN2(n557), .IN3(n24847), .IN4(n600), .IN5(
        n2504), .Q(n2497) );
  OA22X1 U2441 ( .IN1(n24855), .IN2(n643), .IN3(n24863), .IN4(n686), .Q(n2504)
         );
  NAND4X0 U2442 ( .IN1(n2505), .IN2(n2506), .IN3(n2507), .IN4(n2508), .QN(
        n2485) );
  OA221X1 U2443 ( .IN1(n24807), .IN2(n41), .IN3(n24815), .IN4(n84), .IN5(n2509), .Q(n2508) );
  OA22X1 U2444 ( .IN1(n24823), .IN2(n127), .IN3(n24831), .IN4(n170), .Q(n2509)
         );
  OA221X1 U2445 ( .IN1(n24775), .IN2(n213), .IN3(n24783), .IN4(n256), .IN5(
        n2510), .Q(n2507) );
  OA22X1 U2446 ( .IN1(n24791), .IN2(n299), .IN3(n24799), .IN4(n342), .Q(n2510)
         );
  OA221X1 U2447 ( .IN1(n24743), .IN2(n385), .IN3(n24751), .IN4(n428), .IN5(
        n2511), .Q(n2506) );
  OA22X1 U2448 ( .IN1(n24759), .IN2(n471), .IN3(n24767), .IN4(n514), .Q(n2511)
         );
  OA221X1 U2449 ( .IN1(n24711), .IN2(n557), .IN3(n24719), .IN4(n600), .IN5(
        n2512), .Q(n2505) );
  OA22X1 U2450 ( .IN1(n24727), .IN2(n643), .IN3(n24735), .IN4(n686), .Q(n2512)
         );
  NAND4X0 U2451 ( .IN1(n2513), .IN2(n2514), .IN3(n2515), .IN4(n2516), .QN(
        n2484) );
  OA221X1 U2452 ( .IN1(n24679), .IN2(n41), .IN3(n24687), .IN4(n84), .IN5(n2517), .Q(n2516) );
  OA22X1 U2453 ( .IN1(n24695), .IN2(n127), .IN3(n24703), .IN4(n170), .Q(n2517)
         );
  OA221X1 U2454 ( .IN1(n24647), .IN2(n213), .IN3(n24655), .IN4(n256), .IN5(
        n2518), .Q(n2515) );
  OA22X1 U2455 ( .IN1(n24663), .IN2(n299), .IN3(n24671), .IN4(n342), .Q(n2518)
         );
  OA221X1 U2456 ( .IN1(n24615), .IN2(n385), .IN3(n24623), .IN4(n428), .IN5(
        n2519), .Q(n2514) );
  OA22X1 U2457 ( .IN1(n24631), .IN2(n471), .IN3(n24639), .IN4(n514), .Q(n2519)
         );
  OA221X1 U2458 ( .IN1(n24583), .IN2(n557), .IN3(n24591), .IN4(n600), .IN5(
        n2520), .Q(n2513) );
  OA22X1 U2459 ( .IN1(n24599), .IN2(n643), .IN3(n24607), .IN4(n686), .Q(n2520)
         );
  OR4X1 U2460 ( .IN1(n2521), .IN2(n2522), .IN3(n2523), .IN4(n2524), .Q(n2201)
         );
  AO221X1 U2461 ( .IN1(n2157), .IN2(n2525), .IN3(n2159), .IN4(n2526), .IN5(
        n2527), .Q(n2524) );
  AO22X1 U2462 ( .IN1(n2162), .IN2(n2528), .IN3(n2164), .IN4(n2529), .Q(n2527)
         );
  NAND4X0 U2463 ( .IN1(n2530), .IN2(n2531), .IN3(n2532), .IN4(n2533), .QN(
        n2529) );
  OA221X1 U2464 ( .IN1(n24550), .IN2(n40), .IN3(n24558), .IN4(n83), .IN5(n2534), .Q(n2533) );
  OA22X1 U2465 ( .IN1(n24566), .IN2(n126), .IN3(n24574), .IN4(n169), .Q(n2534)
         );
  OA221X1 U2466 ( .IN1(n24518), .IN2(n212), .IN3(n24526), .IN4(n255), .IN5(
        n2535), .Q(n2532) );
  OA22X1 U2467 ( .IN1(n24534), .IN2(n298), .IN3(n24542), .IN4(n341), .Q(n2535)
         );
  OA221X1 U2468 ( .IN1(n24486), .IN2(n384), .IN3(n24494), .IN4(n427), .IN5(
        n2536), .Q(n2531) );
  OA22X1 U2469 ( .IN1(n24502), .IN2(n470), .IN3(n24510), .IN4(n513), .Q(n2536)
         );
  OA221X1 U2470 ( .IN1(n24454), .IN2(n556), .IN3(n24462), .IN4(n599), .IN5(
        n2537), .Q(n2530) );
  OA22X1 U2471 ( .IN1(n24470), .IN2(n642), .IN3(n24478), .IN4(n685), .Q(n2537)
         );
  NAND4X0 U2472 ( .IN1(n2538), .IN2(n2539), .IN3(n2540), .IN4(n2541), .QN(
        n2528) );
  OA221X1 U2473 ( .IN1(n24422), .IN2(n40), .IN3(n24430), .IN4(n83), .IN5(n2542), .Q(n2541) );
  OA22X1 U2474 ( .IN1(n24438), .IN2(n126), .IN3(n24446), .IN4(n169), .Q(n2542)
         );
  OA221X1 U2475 ( .IN1(n24390), .IN2(n212), .IN3(n24398), .IN4(n255), .IN5(
        n2543), .Q(n2540) );
  OA22X1 U2476 ( .IN1(n24406), .IN2(n298), .IN3(n24414), .IN4(n341), .Q(n2543)
         );
  OA221X1 U2477 ( .IN1(n24358), .IN2(n384), .IN3(n24366), .IN4(n427), .IN5(
        n2544), .Q(n2539) );
  OA22X1 U2478 ( .IN1(n24374), .IN2(n470), .IN3(n24382), .IN4(n513), .Q(n2544)
         );
  OA221X1 U2479 ( .IN1(n24326), .IN2(n556), .IN3(n24334), .IN4(n599), .IN5(
        n2545), .Q(n2538) );
  OA22X1 U2480 ( .IN1(n24342), .IN2(n642), .IN3(n24350), .IN4(n685), .Q(n2545)
         );
  NAND4X0 U2481 ( .IN1(n2546), .IN2(n2547), .IN3(n2548), .IN4(n2549), .QN(
        n2526) );
  OA221X1 U2482 ( .IN1(n24294), .IN2(n40), .IN3(n24302), .IN4(n83), .IN5(n2550), .Q(n2549) );
  OA22X1 U2483 ( .IN1(n24310), .IN2(n126), .IN3(n24318), .IN4(n169), .Q(n2550)
         );
  OA221X1 U2484 ( .IN1(n24262), .IN2(n212), .IN3(n24270), .IN4(n255), .IN5(
        n2551), .Q(n2548) );
  OA22X1 U2485 ( .IN1(n24278), .IN2(n298), .IN3(n24286), .IN4(n341), .Q(n2551)
         );
  OA221X1 U2486 ( .IN1(n24230), .IN2(n384), .IN3(n24238), .IN4(n427), .IN5(
        n2552), .Q(n2547) );
  OA22X1 U2487 ( .IN1(n24246), .IN2(n470), .IN3(n24254), .IN4(n513), .Q(n2552)
         );
  OA221X1 U2488 ( .IN1(n24198), .IN2(n556), .IN3(n24206), .IN4(n599), .IN5(
        n2553), .Q(n2546) );
  OA22X1 U2489 ( .IN1(n24214), .IN2(n642), .IN3(n24222), .IN4(n685), .Q(n2553)
         );
  NAND4X0 U2490 ( .IN1(n2554), .IN2(n2555), .IN3(n2556), .IN4(n2557), .QN(
        n2525) );
  OA221X1 U2491 ( .IN1(n24166), .IN2(n40), .IN3(n24174), .IN4(n83), .IN5(n2558), .Q(n2557) );
  OA22X1 U2492 ( .IN1(n24182), .IN2(n126), .IN3(n24190), .IN4(n169), .Q(n2558)
         );
  OA221X1 U2493 ( .IN1(n24134), .IN2(n212), .IN3(n24142), .IN4(n255), .IN5(
        n2559), .Q(n2556) );
  OA22X1 U2494 ( .IN1(n24150), .IN2(n298), .IN3(n24158), .IN4(n341), .Q(n2559)
         );
  OA221X1 U2495 ( .IN1(n24102), .IN2(n384), .IN3(n24110), .IN4(n427), .IN5(
        n2560), .Q(n2555) );
  OA22X1 U2496 ( .IN1(n24118), .IN2(n470), .IN3(n24126), .IN4(n513), .Q(n2560)
         );
  OA221X1 U2497 ( .IN1(n24070), .IN2(n556), .IN3(n24078), .IN4(n599), .IN5(
        n2561), .Q(n2554) );
  OA22X1 U2498 ( .IN1(n24086), .IN2(n642), .IN3(n24094), .IN4(n685), .Q(n2561)
         );
  AO221X1 U2499 ( .IN1(n2246), .IN2(n2562), .IN3(n2248), .IN4(n2563), .IN5(
        n2564), .Q(n2523) );
  AO22X1 U2500 ( .IN1(n2251), .IN2(n2565), .IN3(n2253), .IN4(n2566), .Q(n2564)
         );
  NAND4X0 U2501 ( .IN1(n2567), .IN2(n2568), .IN3(n2569), .IN4(n2570), .QN(
        n2566) );
  OA221X1 U2502 ( .IN1(n24038), .IN2(n40), .IN3(n24046), .IN4(n83), .IN5(n2571), .Q(n2570) );
  OA22X1 U2503 ( .IN1(n24054), .IN2(n126), .IN3(n24062), .IN4(n169), .Q(n2571)
         );
  OA221X1 U2504 ( .IN1(n24006), .IN2(n212), .IN3(n24014), .IN4(n255), .IN5(
        n2572), .Q(n2569) );
  OA22X1 U2505 ( .IN1(n24022), .IN2(n298), .IN3(n24030), .IN4(n341), .Q(n2572)
         );
  OA221X1 U2506 ( .IN1(n23974), .IN2(n384), .IN3(n23982), .IN4(n427), .IN5(
        n2573), .Q(n2568) );
  OA22X1 U2507 ( .IN1(n23990), .IN2(n470), .IN3(n23998), .IN4(n513), .Q(n2573)
         );
  OA221X1 U2508 ( .IN1(n23942), .IN2(n556), .IN3(n23950), .IN4(n599), .IN5(
        n2574), .Q(n2567) );
  OA22X1 U2509 ( .IN1(n23958), .IN2(n642), .IN3(n23966), .IN4(n685), .Q(n2574)
         );
  NAND4X0 U2510 ( .IN1(n2575), .IN2(n2576), .IN3(n2577), .IN4(n2578), .QN(
        n2565) );
  OA221X1 U2511 ( .IN1(n23910), .IN2(n40), .IN3(n23918), .IN4(n83), .IN5(n2579), .Q(n2578) );
  OA22X1 U2512 ( .IN1(n23926), .IN2(n126), .IN3(n23934), .IN4(n169), .Q(n2579)
         );
  OA221X1 U2513 ( .IN1(n23878), .IN2(n212), .IN3(n23886), .IN4(n255), .IN5(
        n2580), .Q(n2577) );
  OA22X1 U2514 ( .IN1(n23894), .IN2(n298), .IN3(n23902), .IN4(n341), .Q(n2580)
         );
  OA221X1 U2515 ( .IN1(n23846), .IN2(n384), .IN3(n23854), .IN4(n427), .IN5(
        n2581), .Q(n2576) );
  OA22X1 U2516 ( .IN1(n23862), .IN2(n470), .IN3(n23870), .IN4(n513), .Q(n2581)
         );
  OA221X1 U2517 ( .IN1(n23814), .IN2(n556), .IN3(n23822), .IN4(n599), .IN5(
        n2582), .Q(n2575) );
  OA22X1 U2518 ( .IN1(n23830), .IN2(n642), .IN3(n23838), .IN4(n685), .Q(n2582)
         );
  NAND4X0 U2519 ( .IN1(n2583), .IN2(n2584), .IN3(n2585), .IN4(n2586), .QN(
        n2563) );
  OA221X1 U2520 ( .IN1(n23782), .IN2(n40), .IN3(n23790), .IN4(n83), .IN5(n2587), .Q(n2586) );
  OA22X1 U2521 ( .IN1(n23798), .IN2(n126), .IN3(n23806), .IN4(n169), .Q(n2587)
         );
  OA221X1 U2522 ( .IN1(n23750), .IN2(n212), .IN3(n23758), .IN4(n255), .IN5(
        n2588), .Q(n2585) );
  OA22X1 U2523 ( .IN1(n23766), .IN2(n298), .IN3(n23774), .IN4(n341), .Q(n2588)
         );
  OA221X1 U2524 ( .IN1(n23718), .IN2(n384), .IN3(n23726), .IN4(n427), .IN5(
        n2589), .Q(n2584) );
  OA22X1 U2525 ( .IN1(n23734), .IN2(n470), .IN3(n23742), .IN4(n513), .Q(n2589)
         );
  OA221X1 U2526 ( .IN1(n23686), .IN2(n556), .IN3(n23694), .IN4(n599), .IN5(
        n2590), .Q(n2583) );
  OA22X1 U2527 ( .IN1(n23702), .IN2(n642), .IN3(n23710), .IN4(n685), .Q(n2590)
         );
  NAND4X0 U2528 ( .IN1(n2591), .IN2(n2592), .IN3(n2593), .IN4(n2594), .QN(
        n2562) );
  OA221X1 U2529 ( .IN1(n23654), .IN2(n40), .IN3(n23662), .IN4(n83), .IN5(n2595), .Q(n2594) );
  OA22X1 U2530 ( .IN1(n23670), .IN2(n126), .IN3(n23678), .IN4(n169), .Q(n2595)
         );
  OA221X1 U2531 ( .IN1(n23622), .IN2(n212), .IN3(n23630), .IN4(n255), .IN5(
        n2596), .Q(n2593) );
  OA22X1 U2532 ( .IN1(n23638), .IN2(n298), .IN3(n23646), .IN4(n341), .Q(n2596)
         );
  OA221X1 U2533 ( .IN1(n23590), .IN2(n384), .IN3(n23598), .IN4(n427), .IN5(
        n2597), .Q(n2592) );
  OA22X1 U2534 ( .IN1(n23606), .IN2(n470), .IN3(n23614), .IN4(n513), .Q(n2597)
         );
  OA221X1 U2535 ( .IN1(n23558), .IN2(n556), .IN3(n23566), .IN4(n599), .IN5(
        n2598), .Q(n2591) );
  OA22X1 U2536 ( .IN1(n23574), .IN2(n642), .IN3(n23582), .IN4(n685), .Q(n2598)
         );
  AO221X1 U2537 ( .IN1(n2287), .IN2(n2599), .IN3(n2289), .IN4(n2600), .IN5(
        n2601), .Q(n2522) );
  AO22X1 U2538 ( .IN1(n2292), .IN2(n2602), .IN3(n2294), .IN4(n2603), .Q(n2601)
         );
  NAND4X0 U2539 ( .IN1(n2604), .IN2(n2605), .IN3(n2606), .IN4(n2607), .QN(
        n2603) );
  OA221X1 U2540 ( .IN1(n25574), .IN2(n40), .IN3(n25582), .IN4(n83), .IN5(n2608), .Q(n2607) );
  OA22X1 U2541 ( .IN1(n25590), .IN2(n126), .IN3(n25598), .IN4(n169), .Q(n2608)
         );
  OA221X1 U2542 ( .IN1(n25542), .IN2(n212), .IN3(n25550), .IN4(n255), .IN5(
        n2609), .Q(n2606) );
  OA22X1 U2543 ( .IN1(n25558), .IN2(n298), .IN3(n25566), .IN4(n341), .Q(n2609)
         );
  OA221X1 U2544 ( .IN1(n25510), .IN2(n384), .IN3(n25518), .IN4(n427), .IN5(
        n2610), .Q(n2605) );
  OA22X1 U2545 ( .IN1(n25526), .IN2(n470), .IN3(n25534), .IN4(n513), .Q(n2610)
         );
  OA221X1 U2546 ( .IN1(n25478), .IN2(n556), .IN3(n25486), .IN4(n599), .IN5(
        n2611), .Q(n2604) );
  OA22X1 U2547 ( .IN1(n25494), .IN2(n642), .IN3(n25502), .IN4(n685), .Q(n2611)
         );
  NAND4X0 U2548 ( .IN1(n2612), .IN2(n2613), .IN3(n2614), .IN4(n2615), .QN(
        n2602) );
  OA221X1 U2549 ( .IN1(n25446), .IN2(n40), .IN3(n25454), .IN4(n83), .IN5(n2616), .Q(n2615) );
  OA22X1 U2550 ( .IN1(n25462), .IN2(n126), .IN3(n25470), .IN4(n169), .Q(n2616)
         );
  OA221X1 U2551 ( .IN1(n25414), .IN2(n212), .IN3(n25422), .IN4(n255), .IN5(
        n2617), .Q(n2614) );
  OA22X1 U2552 ( .IN1(n25430), .IN2(n298), .IN3(n25438), .IN4(n341), .Q(n2617)
         );
  OA221X1 U2553 ( .IN1(n25382), .IN2(n384), .IN3(n25390), .IN4(n427), .IN5(
        n2618), .Q(n2613) );
  OA22X1 U2554 ( .IN1(n25398), .IN2(n470), .IN3(n25406), .IN4(n513), .Q(n2618)
         );
  OA221X1 U2555 ( .IN1(n25350), .IN2(n556), .IN3(n25358), .IN4(n599), .IN5(
        n2619), .Q(n2612) );
  OA22X1 U2556 ( .IN1(n25366), .IN2(n642), .IN3(n25374), .IN4(n685), .Q(n2619)
         );
  NAND4X0 U2557 ( .IN1(n2620), .IN2(n2621), .IN3(n2622), .IN4(n2623), .QN(
        n2600) );
  OA221X1 U2558 ( .IN1(n25318), .IN2(n40), .IN3(n25326), .IN4(n83), .IN5(n2624), .Q(n2623) );
  OA22X1 U2559 ( .IN1(n25334), .IN2(n126), .IN3(n25342), .IN4(n169), .Q(n2624)
         );
  OA221X1 U2560 ( .IN1(n25286), .IN2(n212), .IN3(n25294), .IN4(n255), .IN5(
        n2625), .Q(n2622) );
  OA22X1 U2561 ( .IN1(n25302), .IN2(n298), .IN3(n25310), .IN4(n341), .Q(n2625)
         );
  OA221X1 U2562 ( .IN1(n25254), .IN2(n384), .IN3(n25262), .IN4(n427), .IN5(
        n2626), .Q(n2621) );
  OA22X1 U2563 ( .IN1(n25270), .IN2(n470), .IN3(n25278), .IN4(n513), .Q(n2626)
         );
  OA221X1 U2564 ( .IN1(n25222), .IN2(n556), .IN3(n25230), .IN4(n599), .IN5(
        n2627), .Q(n2620) );
  OA22X1 U2565 ( .IN1(n25238), .IN2(n642), .IN3(n25246), .IN4(n685), .Q(n2627)
         );
  NAND4X0 U2566 ( .IN1(n2628), .IN2(n2629), .IN3(n2630), .IN4(n2631), .QN(
        n2599) );
  OA221X1 U2567 ( .IN1(n25190), .IN2(n40), .IN3(n25198), .IN4(n83), .IN5(n2632), .Q(n2631) );
  OA22X1 U2568 ( .IN1(n25206), .IN2(n126), .IN3(n25214), .IN4(n169), .Q(n2632)
         );
  OA221X1 U2569 ( .IN1(n25158), .IN2(n212), .IN3(n25166), .IN4(n255), .IN5(
        n2633), .Q(n2630) );
  OA22X1 U2570 ( .IN1(n25174), .IN2(n298), .IN3(n25182), .IN4(n341), .Q(n2633)
         );
  OA221X1 U2571 ( .IN1(n25126), .IN2(n384), .IN3(n25134), .IN4(n427), .IN5(
        n2634), .Q(n2629) );
  OA22X1 U2572 ( .IN1(n25142), .IN2(n470), .IN3(n25150), .IN4(n513), .Q(n2634)
         );
  OA221X1 U2573 ( .IN1(n25094), .IN2(n556), .IN3(n25102), .IN4(n599), .IN5(
        n2635), .Q(n2628) );
  OA22X1 U2574 ( .IN1(n25110), .IN2(n642), .IN3(n25118), .IN4(n685), .Q(n2635)
         );
  AO221X1 U2575 ( .IN1(n2328), .IN2(n2636), .IN3(n2330), .IN4(n2637), .IN5(
        n2638), .Q(n2521) );
  AO22X1 U2576 ( .IN1(n2333), .IN2(n2639), .IN3(n2335), .IN4(n2640), .Q(n2638)
         );
  NAND4X0 U2577 ( .IN1(n2641), .IN2(n2642), .IN3(n2643), .IN4(n2644), .QN(
        n2640) );
  OA221X1 U2578 ( .IN1(n25062), .IN2(n39), .IN3(n25070), .IN4(n82), .IN5(n2645), .Q(n2644) );
  OA22X1 U2579 ( .IN1(n25078), .IN2(n125), .IN3(n25086), .IN4(n168), .Q(n2645)
         );
  OA221X1 U2580 ( .IN1(n25030), .IN2(n211), .IN3(n25038), .IN4(n254), .IN5(
        n2646), .Q(n2643) );
  OA22X1 U2581 ( .IN1(n25046), .IN2(n297), .IN3(n25054), .IN4(n340), .Q(n2646)
         );
  OA221X1 U2582 ( .IN1(n24998), .IN2(n383), .IN3(n25006), .IN4(n426), .IN5(
        n2647), .Q(n2642) );
  OA22X1 U2583 ( .IN1(n25014), .IN2(n469), .IN3(n25022), .IN4(n512), .Q(n2647)
         );
  OA221X1 U2584 ( .IN1(n24966), .IN2(n555), .IN3(n24974), .IN4(n598), .IN5(
        n2648), .Q(n2641) );
  OA22X1 U2585 ( .IN1(n24982), .IN2(n641), .IN3(n24990), .IN4(n684), .Q(n2648)
         );
  NAND4X0 U2586 ( .IN1(n2649), .IN2(n2650), .IN3(n2651), .IN4(n2652), .QN(
        n2639) );
  OA221X1 U2587 ( .IN1(n24934), .IN2(n39), .IN3(n24942), .IN4(n82), .IN5(n2653), .Q(n2652) );
  OA22X1 U2588 ( .IN1(n24950), .IN2(n125), .IN3(n24958), .IN4(n168), .Q(n2653)
         );
  OA221X1 U2589 ( .IN1(n24902), .IN2(n211), .IN3(n24910), .IN4(n254), .IN5(
        n2654), .Q(n2651) );
  OA22X1 U2590 ( .IN1(n24918), .IN2(n297), .IN3(n24926), .IN4(n340), .Q(n2654)
         );
  OA221X1 U2591 ( .IN1(n24870), .IN2(n383), .IN3(n24878), .IN4(n426), .IN5(
        n2655), .Q(n2650) );
  OA22X1 U2592 ( .IN1(n24886), .IN2(n469), .IN3(n24894), .IN4(n512), .Q(n2655)
         );
  OA221X1 U2593 ( .IN1(n24838), .IN2(n555), .IN3(n24846), .IN4(n598), .IN5(
        n2656), .Q(n2649) );
  OA22X1 U2594 ( .IN1(n24854), .IN2(n641), .IN3(n24862), .IN4(n684), .Q(n2656)
         );
  NAND4X0 U2595 ( .IN1(n2657), .IN2(n2658), .IN3(n2659), .IN4(n2660), .QN(
        n2637) );
  OA221X1 U2596 ( .IN1(n24806), .IN2(n39), .IN3(n24814), .IN4(n82), .IN5(n2661), .Q(n2660) );
  OA22X1 U2597 ( .IN1(n24822), .IN2(n125), .IN3(n24830), .IN4(n168), .Q(n2661)
         );
  OA221X1 U2598 ( .IN1(n24774), .IN2(n211), .IN3(n24782), .IN4(n254), .IN5(
        n2662), .Q(n2659) );
  OA22X1 U2599 ( .IN1(n24790), .IN2(n297), .IN3(n24798), .IN4(n340), .Q(n2662)
         );
  OA221X1 U2600 ( .IN1(n24742), .IN2(n383), .IN3(n24750), .IN4(n426), .IN5(
        n2663), .Q(n2658) );
  OA22X1 U2601 ( .IN1(n24758), .IN2(n469), .IN3(n24766), .IN4(n512), .Q(n2663)
         );
  OA221X1 U2602 ( .IN1(n24710), .IN2(n555), .IN3(n24718), .IN4(n598), .IN5(
        n2664), .Q(n2657) );
  OA22X1 U2603 ( .IN1(n24726), .IN2(n641), .IN3(n24734), .IN4(n684), .Q(n2664)
         );
  NAND4X0 U2604 ( .IN1(n2665), .IN2(n2666), .IN3(n2667), .IN4(n2668), .QN(
        n2636) );
  OA221X1 U2605 ( .IN1(n24678), .IN2(n39), .IN3(n24686), .IN4(n82), .IN5(n2669), .Q(n2668) );
  OA22X1 U2606 ( .IN1(n24694), .IN2(n125), .IN3(n24702), .IN4(n168), .Q(n2669)
         );
  OA221X1 U2607 ( .IN1(n24646), .IN2(n211), .IN3(n24654), .IN4(n254), .IN5(
        n2670), .Q(n2667) );
  OA22X1 U2608 ( .IN1(n24662), .IN2(n297), .IN3(n24670), .IN4(n340), .Q(n2670)
         );
  OA221X1 U2609 ( .IN1(n24614), .IN2(n383), .IN3(n24622), .IN4(n426), .IN5(
        n2671), .Q(n2666) );
  OA22X1 U2610 ( .IN1(n24630), .IN2(n469), .IN3(n24638), .IN4(n512), .Q(n2671)
         );
  OA221X1 U2611 ( .IN1(n24582), .IN2(n555), .IN3(n24590), .IN4(n598), .IN5(
        n2672), .Q(n2665) );
  OA22X1 U2612 ( .IN1(n24598), .IN2(n641), .IN3(n24606), .IN4(n684), .Q(n2672)
         );
  OR4X1 U2613 ( .IN1(n2673), .IN2(n2674), .IN3(n2675), .IN4(n2676), .Q(n2200)
         );
  AO221X1 U2614 ( .IN1(n2157), .IN2(n2677), .IN3(n2159), .IN4(n2678), .IN5(
        n2679), .Q(n2676) );
  AO22X1 U2615 ( .IN1(n2162), .IN2(n2680), .IN3(n2164), .IN4(n2681), .Q(n2679)
         );
  NAND4X0 U2616 ( .IN1(n2682), .IN2(n2683), .IN3(n2684), .IN4(n2685), .QN(
        n2681) );
  OA221X1 U2617 ( .IN1(n24549), .IN2(n39), .IN3(n24557), .IN4(n82), .IN5(n2686), .Q(n2685) );
  OA22X1 U2618 ( .IN1(n24565), .IN2(n125), .IN3(n24573), .IN4(n168), .Q(n2686)
         );
  OA221X1 U2619 ( .IN1(n24517), .IN2(n211), .IN3(n24525), .IN4(n254), .IN5(
        n2687), .Q(n2684) );
  OA22X1 U2620 ( .IN1(n24533), .IN2(n297), .IN3(n24541), .IN4(n340), .Q(n2687)
         );
  OA221X1 U2621 ( .IN1(n24485), .IN2(n383), .IN3(n24493), .IN4(n426), .IN5(
        n2688), .Q(n2683) );
  OA22X1 U2622 ( .IN1(n24501), .IN2(n469), .IN3(n24509), .IN4(n512), .Q(n2688)
         );
  OA221X1 U2623 ( .IN1(n24453), .IN2(n555), .IN3(n24461), .IN4(n598), .IN5(
        n2689), .Q(n2682) );
  OA22X1 U2624 ( .IN1(n24469), .IN2(n641), .IN3(n24477), .IN4(n684), .Q(n2689)
         );
  NAND4X0 U2625 ( .IN1(n2690), .IN2(n2691), .IN3(n2692), .IN4(n2693), .QN(
        n2680) );
  OA221X1 U2626 ( .IN1(n24421), .IN2(n39), .IN3(n24429), .IN4(n82), .IN5(n2694), .Q(n2693) );
  OA22X1 U2627 ( .IN1(n24437), .IN2(n125), .IN3(n24445), .IN4(n168), .Q(n2694)
         );
  OA221X1 U2628 ( .IN1(n24389), .IN2(n211), .IN3(n24397), .IN4(n254), .IN5(
        n2695), .Q(n2692) );
  OA22X1 U2629 ( .IN1(n24405), .IN2(n297), .IN3(n24413), .IN4(n340), .Q(n2695)
         );
  OA221X1 U2630 ( .IN1(n24357), .IN2(n383), .IN3(n24365), .IN4(n426), .IN5(
        n2696), .Q(n2691) );
  OA22X1 U2631 ( .IN1(n24373), .IN2(n469), .IN3(n24381), .IN4(n512), .Q(n2696)
         );
  OA221X1 U2632 ( .IN1(n24325), .IN2(n555), .IN3(n24333), .IN4(n598), .IN5(
        n2697), .Q(n2690) );
  OA22X1 U2633 ( .IN1(n24341), .IN2(n641), .IN3(n24349), .IN4(n684), .Q(n2697)
         );
  NAND4X0 U2634 ( .IN1(n2698), .IN2(n2699), .IN3(n2700), .IN4(n2701), .QN(
        n2678) );
  OA221X1 U2635 ( .IN1(n24293), .IN2(n39), .IN3(n24301), .IN4(n82), .IN5(n2702), .Q(n2701) );
  OA22X1 U2636 ( .IN1(n24309), .IN2(n125), .IN3(n24317), .IN4(n168), .Q(n2702)
         );
  OA221X1 U2637 ( .IN1(n24261), .IN2(n211), .IN3(n24269), .IN4(n254), .IN5(
        n2703), .Q(n2700) );
  OA22X1 U2638 ( .IN1(n24277), .IN2(n297), .IN3(n24285), .IN4(n340), .Q(n2703)
         );
  OA221X1 U2639 ( .IN1(n24229), .IN2(n383), .IN3(n24237), .IN4(n426), .IN5(
        n2704), .Q(n2699) );
  OA22X1 U2640 ( .IN1(n24245), .IN2(n469), .IN3(n24253), .IN4(n512), .Q(n2704)
         );
  OA221X1 U2641 ( .IN1(n24197), .IN2(n555), .IN3(n24205), .IN4(n598), .IN5(
        n2705), .Q(n2698) );
  OA22X1 U2642 ( .IN1(n24213), .IN2(n641), .IN3(n24221), .IN4(n684), .Q(n2705)
         );
  NAND4X0 U2643 ( .IN1(n2706), .IN2(n2707), .IN3(n2708), .IN4(n2709), .QN(
        n2677) );
  OA221X1 U2644 ( .IN1(n24165), .IN2(n39), .IN3(n24173), .IN4(n82), .IN5(n2710), .Q(n2709) );
  OA22X1 U2645 ( .IN1(n24181), .IN2(n125), .IN3(n24189), .IN4(n168), .Q(n2710)
         );
  OA221X1 U2646 ( .IN1(n24133), .IN2(n211), .IN3(n24141), .IN4(n254), .IN5(
        n2711), .Q(n2708) );
  OA22X1 U2647 ( .IN1(n24149), .IN2(n297), .IN3(n24157), .IN4(n340), .Q(n2711)
         );
  OA221X1 U2648 ( .IN1(n24101), .IN2(n383), .IN3(n24109), .IN4(n426), .IN5(
        n2712), .Q(n2707) );
  OA22X1 U2649 ( .IN1(n24117), .IN2(n469), .IN3(n24125), .IN4(n512), .Q(n2712)
         );
  OA221X1 U2650 ( .IN1(n24069), .IN2(n555), .IN3(n24077), .IN4(n598), .IN5(
        n2713), .Q(n2706) );
  OA22X1 U2651 ( .IN1(n24085), .IN2(n641), .IN3(n24093), .IN4(n684), .Q(n2713)
         );
  AO221X1 U2652 ( .IN1(n2246), .IN2(n2714), .IN3(n2248), .IN4(n2715), .IN5(
        n2716), .Q(n2675) );
  AO22X1 U2653 ( .IN1(n2251), .IN2(n2717), .IN3(n2253), .IN4(n2718), .Q(n2716)
         );
  NAND4X0 U2654 ( .IN1(n2719), .IN2(n2720), .IN3(n2721), .IN4(n2722), .QN(
        n2718) );
  OA221X1 U2655 ( .IN1(n24037), .IN2(n39), .IN3(n24045), .IN4(n82), .IN5(n2723), .Q(n2722) );
  OA22X1 U2656 ( .IN1(n24053), .IN2(n125), .IN3(n24061), .IN4(n168), .Q(n2723)
         );
  OA221X1 U2657 ( .IN1(n24005), .IN2(n211), .IN3(n24013), .IN4(n254), .IN5(
        n2724), .Q(n2721) );
  OA22X1 U2658 ( .IN1(n24021), .IN2(n297), .IN3(n24029), .IN4(n340), .Q(n2724)
         );
  OA221X1 U2659 ( .IN1(n23973), .IN2(n383), .IN3(n23981), .IN4(n426), .IN5(
        n2725), .Q(n2720) );
  OA22X1 U2660 ( .IN1(n23989), .IN2(n469), .IN3(n23997), .IN4(n512), .Q(n2725)
         );
  OA221X1 U2661 ( .IN1(n23941), .IN2(n555), .IN3(n23949), .IN4(n598), .IN5(
        n2726), .Q(n2719) );
  OA22X1 U2662 ( .IN1(n23957), .IN2(n641), .IN3(n23965), .IN4(n684), .Q(n2726)
         );
  NAND4X0 U2663 ( .IN1(n2727), .IN2(n2728), .IN3(n2729), .IN4(n2730), .QN(
        n2717) );
  OA221X1 U2664 ( .IN1(n23909), .IN2(n39), .IN3(n23917), .IN4(n82), .IN5(n2731), .Q(n2730) );
  OA22X1 U2665 ( .IN1(n23925), .IN2(n125), .IN3(n23933), .IN4(n168), .Q(n2731)
         );
  OA221X1 U2666 ( .IN1(n23877), .IN2(n211), .IN3(n23885), .IN4(n254), .IN5(
        n2732), .Q(n2729) );
  OA22X1 U2667 ( .IN1(n23893), .IN2(n297), .IN3(n23901), .IN4(n340), .Q(n2732)
         );
  OA221X1 U2668 ( .IN1(n23845), .IN2(n383), .IN3(n23853), .IN4(n426), .IN5(
        n2733), .Q(n2728) );
  OA22X1 U2669 ( .IN1(n23861), .IN2(n469), .IN3(n23869), .IN4(n512), .Q(n2733)
         );
  OA221X1 U2670 ( .IN1(n23813), .IN2(n555), .IN3(n23821), .IN4(n598), .IN5(
        n2734), .Q(n2727) );
  OA22X1 U2671 ( .IN1(n23829), .IN2(n641), .IN3(n23837), .IN4(n684), .Q(n2734)
         );
  NAND4X0 U2672 ( .IN1(n2735), .IN2(n2736), .IN3(n2737), .IN4(n2738), .QN(
        n2715) );
  OA221X1 U2673 ( .IN1(n23781), .IN2(n39), .IN3(n23789), .IN4(n82), .IN5(n2739), .Q(n2738) );
  OA22X1 U2674 ( .IN1(n23797), .IN2(n125), .IN3(n23805), .IN4(n168), .Q(n2739)
         );
  OA221X1 U2675 ( .IN1(n23749), .IN2(n211), .IN3(n23757), .IN4(n254), .IN5(
        n2740), .Q(n2737) );
  OA22X1 U2676 ( .IN1(n23765), .IN2(n297), .IN3(n23773), .IN4(n340), .Q(n2740)
         );
  OA221X1 U2677 ( .IN1(n23717), .IN2(n383), .IN3(n23725), .IN4(n426), .IN5(
        n2741), .Q(n2736) );
  OA22X1 U2678 ( .IN1(n23733), .IN2(n469), .IN3(n23741), .IN4(n512), .Q(n2741)
         );
  OA221X1 U2679 ( .IN1(n23685), .IN2(n555), .IN3(n23693), .IN4(n598), .IN5(
        n2742), .Q(n2735) );
  OA22X1 U2680 ( .IN1(n23701), .IN2(n641), .IN3(n23709), .IN4(n684), .Q(n2742)
         );
  NAND4X0 U2681 ( .IN1(n2743), .IN2(n2744), .IN3(n2745), .IN4(n2746), .QN(
        n2714) );
  OA221X1 U2682 ( .IN1(n23653), .IN2(n39), .IN3(n23661), .IN4(n82), .IN5(n2747), .Q(n2746) );
  OA22X1 U2683 ( .IN1(n23669), .IN2(n125), .IN3(n23677), .IN4(n168), .Q(n2747)
         );
  OA221X1 U2684 ( .IN1(n23621), .IN2(n211), .IN3(n23629), .IN4(n254), .IN5(
        n2748), .Q(n2745) );
  OA22X1 U2685 ( .IN1(n23637), .IN2(n297), .IN3(n23645), .IN4(n340), .Q(n2748)
         );
  OA221X1 U2686 ( .IN1(n23589), .IN2(n383), .IN3(n23597), .IN4(n426), .IN5(
        n2749), .Q(n2744) );
  OA22X1 U2687 ( .IN1(n23605), .IN2(n469), .IN3(n23613), .IN4(n512), .Q(n2749)
         );
  OA221X1 U2688 ( .IN1(n23557), .IN2(n555), .IN3(n23565), .IN4(n598), .IN5(
        n2750), .Q(n2743) );
  OA22X1 U2689 ( .IN1(n23573), .IN2(n641), .IN3(n23581), .IN4(n684), .Q(n2750)
         );
  AO221X1 U2690 ( .IN1(n2287), .IN2(n2751), .IN3(n2289), .IN4(n2752), .IN5(
        n2753), .Q(n2674) );
  AO22X1 U2691 ( .IN1(n2292), .IN2(n2754), .IN3(n2294), .IN4(n2755), .Q(n2753)
         );
  NAND4X0 U2692 ( .IN1(n2756), .IN2(n2757), .IN3(n2758), .IN4(n2759), .QN(
        n2755) );
  OA221X1 U2693 ( .IN1(n25573), .IN2(n38), .IN3(n25581), .IN4(n81), .IN5(n2760), .Q(n2759) );
  OA22X1 U2694 ( .IN1(n25589), .IN2(n124), .IN3(n25597), .IN4(n167), .Q(n2760)
         );
  OA221X1 U2695 ( .IN1(n25541), .IN2(n210), .IN3(n25549), .IN4(n253), .IN5(
        n2761), .Q(n2758) );
  OA22X1 U2696 ( .IN1(n25557), .IN2(n296), .IN3(n25565), .IN4(n339), .Q(n2761)
         );
  OA221X1 U2697 ( .IN1(n25509), .IN2(n382), .IN3(n25517), .IN4(n425), .IN5(
        n2762), .Q(n2757) );
  OA22X1 U2698 ( .IN1(n25525), .IN2(n468), .IN3(n25533), .IN4(n511), .Q(n2762)
         );
  OA221X1 U2699 ( .IN1(n25477), .IN2(n554), .IN3(n25485), .IN4(n597), .IN5(
        n2763), .Q(n2756) );
  OA22X1 U2700 ( .IN1(n25493), .IN2(n640), .IN3(n25501), .IN4(n683), .Q(n2763)
         );
  NAND4X0 U2701 ( .IN1(n2764), .IN2(n2765), .IN3(n2766), .IN4(n2767), .QN(
        n2754) );
  OA221X1 U2702 ( .IN1(n25445), .IN2(n38), .IN3(n25453), .IN4(n81), .IN5(n2768), .Q(n2767) );
  OA22X1 U2703 ( .IN1(n25461), .IN2(n124), .IN3(n25469), .IN4(n167), .Q(n2768)
         );
  OA221X1 U2704 ( .IN1(n25413), .IN2(n210), .IN3(n25421), .IN4(n253), .IN5(
        n2769), .Q(n2766) );
  OA22X1 U2705 ( .IN1(n25429), .IN2(n296), .IN3(n25437), .IN4(n339), .Q(n2769)
         );
  OA221X1 U2706 ( .IN1(n25381), .IN2(n382), .IN3(n25389), .IN4(n425), .IN5(
        n2770), .Q(n2765) );
  OA22X1 U2707 ( .IN1(n25397), .IN2(n468), .IN3(n25405), .IN4(n511), .Q(n2770)
         );
  OA221X1 U2708 ( .IN1(n25349), .IN2(n554), .IN3(n25357), .IN4(n597), .IN5(
        n2771), .Q(n2764) );
  OA22X1 U2709 ( .IN1(n25365), .IN2(n640), .IN3(n25373), .IN4(n683), .Q(n2771)
         );
  NAND4X0 U2710 ( .IN1(n2772), .IN2(n2773), .IN3(n2774), .IN4(n2775), .QN(
        n2752) );
  OA221X1 U2711 ( .IN1(n25317), .IN2(n38), .IN3(n25325), .IN4(n81), .IN5(n2776), .Q(n2775) );
  OA22X1 U2712 ( .IN1(n25333), .IN2(n124), .IN3(n25341), .IN4(n167), .Q(n2776)
         );
  OA221X1 U2713 ( .IN1(n25285), .IN2(n210), .IN3(n25293), .IN4(n253), .IN5(
        n2777), .Q(n2774) );
  OA22X1 U2714 ( .IN1(n25301), .IN2(n296), .IN3(n25309), .IN4(n339), .Q(n2777)
         );
  OA221X1 U2715 ( .IN1(n25253), .IN2(n382), .IN3(n25261), .IN4(n425), .IN5(
        n2778), .Q(n2773) );
  OA22X1 U2716 ( .IN1(n25269), .IN2(n468), .IN3(n25277), .IN4(n511), .Q(n2778)
         );
  OA221X1 U2717 ( .IN1(n25221), .IN2(n554), .IN3(n25229), .IN4(n597), .IN5(
        n2779), .Q(n2772) );
  OA22X1 U2718 ( .IN1(n25237), .IN2(n640), .IN3(n25245), .IN4(n683), .Q(n2779)
         );
  NAND4X0 U2719 ( .IN1(n2780), .IN2(n2781), .IN3(n2782), .IN4(n2783), .QN(
        n2751) );
  OA221X1 U2720 ( .IN1(n25189), .IN2(n38), .IN3(n25197), .IN4(n81), .IN5(n2784), .Q(n2783) );
  OA22X1 U2721 ( .IN1(n25205), .IN2(n124), .IN3(n25213), .IN4(n167), .Q(n2784)
         );
  OA221X1 U2722 ( .IN1(n25157), .IN2(n210), .IN3(n25165), .IN4(n253), .IN5(
        n2785), .Q(n2782) );
  OA22X1 U2723 ( .IN1(n25173), .IN2(n296), .IN3(n25181), .IN4(n339), .Q(n2785)
         );
  OA221X1 U2724 ( .IN1(n25125), .IN2(n382), .IN3(n25133), .IN4(n425), .IN5(
        n2786), .Q(n2781) );
  OA22X1 U2725 ( .IN1(n25141), .IN2(n468), .IN3(n25149), .IN4(n511), .Q(n2786)
         );
  OA221X1 U2726 ( .IN1(n25093), .IN2(n554), .IN3(n25101), .IN4(n597), .IN5(
        n2787), .Q(n2780) );
  OA22X1 U2727 ( .IN1(n25109), .IN2(n640), .IN3(n25117), .IN4(n683), .Q(n2787)
         );
  AO221X1 U2728 ( .IN1(n2328), .IN2(n2788), .IN3(n2330), .IN4(n2789), .IN5(
        n2790), .Q(n2673) );
  AO22X1 U2729 ( .IN1(n2333), .IN2(n2791), .IN3(n2335), .IN4(n2792), .Q(n2790)
         );
  NAND4X0 U2730 ( .IN1(n2793), .IN2(n2794), .IN3(n2795), .IN4(n2796), .QN(
        n2792) );
  OA221X1 U2731 ( .IN1(n25061), .IN2(n38), .IN3(n25069), .IN4(n81), .IN5(n2797), .Q(n2796) );
  OA22X1 U2732 ( .IN1(n25077), .IN2(n124), .IN3(n25085), .IN4(n167), .Q(n2797)
         );
  OA221X1 U2733 ( .IN1(n25029), .IN2(n210), .IN3(n25037), .IN4(n253), .IN5(
        n2798), .Q(n2795) );
  OA22X1 U2734 ( .IN1(n25045), .IN2(n296), .IN3(n25053), .IN4(n339), .Q(n2798)
         );
  OA221X1 U2735 ( .IN1(n24997), .IN2(n382), .IN3(n25005), .IN4(n425), .IN5(
        n2799), .Q(n2794) );
  OA22X1 U2736 ( .IN1(n25013), .IN2(n468), .IN3(n25021), .IN4(n511), .Q(n2799)
         );
  OA221X1 U2737 ( .IN1(n24965), .IN2(n554), .IN3(n24973), .IN4(n597), .IN5(
        n2800), .Q(n2793) );
  OA22X1 U2738 ( .IN1(n24981), .IN2(n640), .IN3(n24989), .IN4(n683), .Q(n2800)
         );
  NAND4X0 U2739 ( .IN1(n2801), .IN2(n2802), .IN3(n2803), .IN4(n2804), .QN(
        n2791) );
  OA221X1 U2740 ( .IN1(n24933), .IN2(n38), .IN3(n24941), .IN4(n81), .IN5(n2805), .Q(n2804) );
  OA22X1 U2741 ( .IN1(n24949), .IN2(n124), .IN3(n24957), .IN4(n167), .Q(n2805)
         );
  OA221X1 U2742 ( .IN1(n24901), .IN2(n210), .IN3(n24909), .IN4(n253), .IN5(
        n2806), .Q(n2803) );
  OA22X1 U2743 ( .IN1(n24917), .IN2(n296), .IN3(n24925), .IN4(n339), .Q(n2806)
         );
  OA221X1 U2744 ( .IN1(n24869), .IN2(n382), .IN3(n24877), .IN4(n425), .IN5(
        n2807), .Q(n2802) );
  OA22X1 U2745 ( .IN1(n24885), .IN2(n468), .IN3(n24893), .IN4(n511), .Q(n2807)
         );
  OA221X1 U2746 ( .IN1(n24837), .IN2(n554), .IN3(n24845), .IN4(n597), .IN5(
        n2808), .Q(n2801) );
  OA22X1 U2747 ( .IN1(n24853), .IN2(n640), .IN3(n24861), .IN4(n683), .Q(n2808)
         );
  NAND4X0 U2748 ( .IN1(n2809), .IN2(n2810), .IN3(n2811), .IN4(n2812), .QN(
        n2789) );
  OA221X1 U2749 ( .IN1(n24805), .IN2(n38), .IN3(n24813), .IN4(n81), .IN5(n2813), .Q(n2812) );
  OA22X1 U2750 ( .IN1(n24821), .IN2(n124), .IN3(n24829), .IN4(n167), .Q(n2813)
         );
  OA221X1 U2751 ( .IN1(n24773), .IN2(n210), .IN3(n24781), .IN4(n253), .IN5(
        n2814), .Q(n2811) );
  OA22X1 U2752 ( .IN1(n24789), .IN2(n296), .IN3(n24797), .IN4(n339), .Q(n2814)
         );
  OA221X1 U2753 ( .IN1(n24741), .IN2(n382), .IN3(n24749), .IN4(n425), .IN5(
        n2815), .Q(n2810) );
  OA22X1 U2754 ( .IN1(n24757), .IN2(n468), .IN3(n24765), .IN4(n511), .Q(n2815)
         );
  OA221X1 U2755 ( .IN1(n24709), .IN2(n554), .IN3(n24717), .IN4(n597), .IN5(
        n2816), .Q(n2809) );
  OA22X1 U2756 ( .IN1(n24725), .IN2(n640), .IN3(n24733), .IN4(n683), .Q(n2816)
         );
  NAND4X0 U2757 ( .IN1(n2817), .IN2(n2818), .IN3(n2819), .IN4(n2820), .QN(
        n2788) );
  OA221X1 U2758 ( .IN1(n24677), .IN2(n38), .IN3(n24685), .IN4(n81), .IN5(n2821), .Q(n2820) );
  OA22X1 U2759 ( .IN1(n24693), .IN2(n124), .IN3(n24701), .IN4(n167), .Q(n2821)
         );
  OA221X1 U2760 ( .IN1(n24645), .IN2(n210), .IN3(n24653), .IN4(n253), .IN5(
        n2822), .Q(n2819) );
  OA22X1 U2761 ( .IN1(n24661), .IN2(n296), .IN3(n24669), .IN4(n339), .Q(n2822)
         );
  OA221X1 U2762 ( .IN1(n24613), .IN2(n382), .IN3(n24621), .IN4(n425), .IN5(
        n2823), .Q(n2818) );
  OA22X1 U2763 ( .IN1(n24629), .IN2(n468), .IN3(n24637), .IN4(n511), .Q(n2823)
         );
  OA221X1 U2764 ( .IN1(n24581), .IN2(n554), .IN3(n24589), .IN4(n597), .IN5(
        n2824), .Q(n2817) );
  OA22X1 U2765 ( .IN1(n24597), .IN2(n640), .IN3(n24605), .IN4(n683), .Q(n2824)
         );
  OR4X1 U2766 ( .IN1(n2825), .IN2(n2826), .IN3(n2827), .IN4(n2828), .Q(n2199)
         );
  AO221X1 U2767 ( .IN1(n2157), .IN2(n2829), .IN3(n2159), .IN4(n2830), .IN5(
        n2831), .Q(n2828) );
  AO22X1 U2768 ( .IN1(n2162), .IN2(n2832), .IN3(n2164), .IN4(n2833), .Q(n2831)
         );
  NAND4X0 U2769 ( .IN1(n2834), .IN2(n2835), .IN3(n2836), .IN4(n2837), .QN(
        n2833) );
  OA221X1 U2770 ( .IN1(n24548), .IN2(n38), .IN3(n24556), .IN4(n81), .IN5(n2838), .Q(n2837) );
  OA22X1 U2771 ( .IN1(n24564), .IN2(n124), .IN3(n24572), .IN4(n167), .Q(n2838)
         );
  OA221X1 U2772 ( .IN1(n24516), .IN2(n210), .IN3(n24524), .IN4(n253), .IN5(
        n2839), .Q(n2836) );
  OA22X1 U2773 ( .IN1(n24532), .IN2(n296), .IN3(n24540), .IN4(n339), .Q(n2839)
         );
  OA221X1 U2774 ( .IN1(n24484), .IN2(n382), .IN3(n24492), .IN4(n425), .IN5(
        n2840), .Q(n2835) );
  OA22X1 U2775 ( .IN1(n24500), .IN2(n468), .IN3(n24508), .IN4(n511), .Q(n2840)
         );
  OA221X1 U2776 ( .IN1(n24452), .IN2(n554), .IN3(n24460), .IN4(n597), .IN5(
        n2841), .Q(n2834) );
  OA22X1 U2777 ( .IN1(n24468), .IN2(n640), .IN3(n24476), .IN4(n683), .Q(n2841)
         );
  NAND4X0 U2778 ( .IN1(n2842), .IN2(n2843), .IN3(n2844), .IN4(n2845), .QN(
        n2832) );
  OA221X1 U2779 ( .IN1(n24420), .IN2(n38), .IN3(n24428), .IN4(n81), .IN5(n2846), .Q(n2845) );
  OA22X1 U2780 ( .IN1(n24436), .IN2(n124), .IN3(n24444), .IN4(n167), .Q(n2846)
         );
  OA221X1 U2781 ( .IN1(n24388), .IN2(n210), .IN3(n24396), .IN4(n253), .IN5(
        n2847), .Q(n2844) );
  OA22X1 U2782 ( .IN1(n24404), .IN2(n296), .IN3(n24412), .IN4(n339), .Q(n2847)
         );
  OA221X1 U2783 ( .IN1(n24356), .IN2(n382), .IN3(n24364), .IN4(n425), .IN5(
        n2848), .Q(n2843) );
  OA22X1 U2784 ( .IN1(n24372), .IN2(n468), .IN3(n24380), .IN4(n511), .Q(n2848)
         );
  OA221X1 U2785 ( .IN1(n24324), .IN2(n554), .IN3(n24332), .IN4(n597), .IN5(
        n2849), .Q(n2842) );
  OA22X1 U2786 ( .IN1(n24340), .IN2(n640), .IN3(n24348), .IN4(n683), .Q(n2849)
         );
  NAND4X0 U2787 ( .IN1(n2850), .IN2(n2851), .IN3(n2852), .IN4(n2853), .QN(
        n2830) );
  OA221X1 U2788 ( .IN1(n24292), .IN2(n38), .IN3(n24300), .IN4(n81), .IN5(n2854), .Q(n2853) );
  OA22X1 U2789 ( .IN1(n24308), .IN2(n124), .IN3(n24316), .IN4(n167), .Q(n2854)
         );
  OA221X1 U2790 ( .IN1(n24260), .IN2(n210), .IN3(n24268), .IN4(n253), .IN5(
        n2855), .Q(n2852) );
  OA22X1 U2791 ( .IN1(n24276), .IN2(n296), .IN3(n24284), .IN4(n339), .Q(n2855)
         );
  OA221X1 U2792 ( .IN1(n24228), .IN2(n382), .IN3(n24236), .IN4(n425), .IN5(
        n2856), .Q(n2851) );
  OA22X1 U2793 ( .IN1(n24244), .IN2(n468), .IN3(n24252), .IN4(n511), .Q(n2856)
         );
  OA221X1 U2794 ( .IN1(n24196), .IN2(n554), .IN3(n24204), .IN4(n597), .IN5(
        n2857), .Q(n2850) );
  OA22X1 U2795 ( .IN1(n24212), .IN2(n640), .IN3(n24220), .IN4(n683), .Q(n2857)
         );
  NAND4X0 U2796 ( .IN1(n2858), .IN2(n2859), .IN3(n2860), .IN4(n2861), .QN(
        n2829) );
  OA221X1 U2797 ( .IN1(n24164), .IN2(n38), .IN3(n24172), .IN4(n81), .IN5(n2862), .Q(n2861) );
  OA22X1 U2798 ( .IN1(n24180), .IN2(n124), .IN3(n24188), .IN4(n167), .Q(n2862)
         );
  OA221X1 U2799 ( .IN1(n24132), .IN2(n210), .IN3(n24140), .IN4(n253), .IN5(
        n2863), .Q(n2860) );
  OA22X1 U2800 ( .IN1(n24148), .IN2(n296), .IN3(n24156), .IN4(n339), .Q(n2863)
         );
  OA221X1 U2801 ( .IN1(n24100), .IN2(n382), .IN3(n24108), .IN4(n425), .IN5(
        n2864), .Q(n2859) );
  OA22X1 U2802 ( .IN1(n24116), .IN2(n468), .IN3(n24124), .IN4(n511), .Q(n2864)
         );
  OA221X1 U2803 ( .IN1(n24068), .IN2(n554), .IN3(n24076), .IN4(n597), .IN5(
        n2865), .Q(n2858) );
  OA22X1 U2804 ( .IN1(n24084), .IN2(n640), .IN3(n24092), .IN4(n683), .Q(n2865)
         );
  AO221X1 U2805 ( .IN1(n2246), .IN2(n2866), .IN3(n2248), .IN4(n2867), .IN5(
        n2868), .Q(n2827) );
  AO22X1 U2806 ( .IN1(n2251), .IN2(n2869), .IN3(n2253), .IN4(n2870), .Q(n2868)
         );
  NAND4X0 U2807 ( .IN1(n2871), .IN2(n2872), .IN3(n2873), .IN4(n2874), .QN(
        n2870) );
  OA221X1 U2808 ( .IN1(n24036), .IN2(n37), .IN3(n24044), .IN4(n80), .IN5(n2875), .Q(n2874) );
  OA22X1 U2809 ( .IN1(n24052), .IN2(n123), .IN3(n24060), .IN4(n166), .Q(n2875)
         );
  OA221X1 U2810 ( .IN1(n24004), .IN2(n209), .IN3(n24012), .IN4(n252), .IN5(
        n2876), .Q(n2873) );
  OA22X1 U2811 ( .IN1(n24020), .IN2(n295), .IN3(n24028), .IN4(n338), .Q(n2876)
         );
  OA221X1 U2812 ( .IN1(n23972), .IN2(n381), .IN3(n23980), .IN4(n424), .IN5(
        n2877), .Q(n2872) );
  OA22X1 U2813 ( .IN1(n23988), .IN2(n467), .IN3(n23996), .IN4(n510), .Q(n2877)
         );
  OA221X1 U2814 ( .IN1(n23940), .IN2(n553), .IN3(n23948), .IN4(n596), .IN5(
        n2878), .Q(n2871) );
  OA22X1 U2815 ( .IN1(n23956), .IN2(n639), .IN3(n23964), .IN4(n682), .Q(n2878)
         );
  NAND4X0 U2816 ( .IN1(n2879), .IN2(n2880), .IN3(n2881), .IN4(n2882), .QN(
        n2869) );
  OA221X1 U2817 ( .IN1(n23908), .IN2(n37), .IN3(n23916), .IN4(n80), .IN5(n2883), .Q(n2882) );
  OA22X1 U2818 ( .IN1(n23924), .IN2(n123), .IN3(n23932), .IN4(n166), .Q(n2883)
         );
  OA221X1 U2819 ( .IN1(n23876), .IN2(n209), .IN3(n23884), .IN4(n252), .IN5(
        n2884), .Q(n2881) );
  OA22X1 U2820 ( .IN1(n23892), .IN2(n295), .IN3(n23900), .IN4(n338), .Q(n2884)
         );
  OA221X1 U2821 ( .IN1(n23844), .IN2(n381), .IN3(n23852), .IN4(n424), .IN5(
        n2885), .Q(n2880) );
  OA22X1 U2822 ( .IN1(n23860), .IN2(n467), .IN3(n23868), .IN4(n510), .Q(n2885)
         );
  OA221X1 U2823 ( .IN1(n23812), .IN2(n553), .IN3(n23820), .IN4(n596), .IN5(
        n2886), .Q(n2879) );
  OA22X1 U2824 ( .IN1(n23828), .IN2(n639), .IN3(n23836), .IN4(n682), .Q(n2886)
         );
  NAND4X0 U2825 ( .IN1(n2887), .IN2(n2888), .IN3(n2889), .IN4(n2890), .QN(
        n2867) );
  OA221X1 U2826 ( .IN1(n23780), .IN2(n37), .IN3(n23788), .IN4(n80), .IN5(n2891), .Q(n2890) );
  OA22X1 U2827 ( .IN1(n23796), .IN2(n123), .IN3(n23804), .IN4(n166), .Q(n2891)
         );
  OA221X1 U2828 ( .IN1(n23748), .IN2(n209), .IN3(n23756), .IN4(n252), .IN5(
        n2892), .Q(n2889) );
  OA22X1 U2829 ( .IN1(n23764), .IN2(n295), .IN3(n23772), .IN4(n338), .Q(n2892)
         );
  OA221X1 U2830 ( .IN1(n23716), .IN2(n381), .IN3(n23724), .IN4(n424), .IN5(
        n2893), .Q(n2888) );
  OA22X1 U2831 ( .IN1(n23732), .IN2(n467), .IN3(n23740), .IN4(n510), .Q(n2893)
         );
  OA221X1 U2832 ( .IN1(n23684), .IN2(n553), .IN3(n23692), .IN4(n596), .IN5(
        n2894), .Q(n2887) );
  OA22X1 U2833 ( .IN1(n23700), .IN2(n639), .IN3(n23708), .IN4(n682), .Q(n2894)
         );
  NAND4X0 U2834 ( .IN1(n2895), .IN2(n2896), .IN3(n2897), .IN4(n2898), .QN(
        n2866) );
  OA221X1 U2835 ( .IN1(n23652), .IN2(n37), .IN3(n23660), .IN4(n80), .IN5(n2899), .Q(n2898) );
  OA22X1 U2836 ( .IN1(n23668), .IN2(n123), .IN3(n23676), .IN4(n166), .Q(n2899)
         );
  OA221X1 U2837 ( .IN1(n23620), .IN2(n209), .IN3(n23628), .IN4(n252), .IN5(
        n2900), .Q(n2897) );
  OA22X1 U2838 ( .IN1(n23636), .IN2(n295), .IN3(n23644), .IN4(n338), .Q(n2900)
         );
  OA221X1 U2839 ( .IN1(n23588), .IN2(n381), .IN3(n23596), .IN4(n424), .IN5(
        n2901), .Q(n2896) );
  OA22X1 U2840 ( .IN1(n23604), .IN2(n467), .IN3(n23612), .IN4(n510), .Q(n2901)
         );
  OA221X1 U2841 ( .IN1(n23556), .IN2(n553), .IN3(n23564), .IN4(n596), .IN5(
        n2902), .Q(n2895) );
  OA22X1 U2842 ( .IN1(n23572), .IN2(n639), .IN3(n23580), .IN4(n682), .Q(n2902)
         );
  AO221X1 U2843 ( .IN1(n2287), .IN2(n2903), .IN3(n2289), .IN4(n2904), .IN5(
        n2905), .Q(n2826) );
  AO22X1 U2844 ( .IN1(n2292), .IN2(n2906), .IN3(n2294), .IN4(n2907), .Q(n2905)
         );
  NAND4X0 U2845 ( .IN1(n2908), .IN2(n2909), .IN3(n2910), .IN4(n2911), .QN(
        n2907) );
  OA221X1 U2846 ( .IN1(n25572), .IN2(n37), .IN3(n25580), .IN4(n80), .IN5(n2912), .Q(n2911) );
  OA22X1 U2847 ( .IN1(n25588), .IN2(n123), .IN3(n25596), .IN4(n166), .Q(n2912)
         );
  OA221X1 U2848 ( .IN1(n25540), .IN2(n209), .IN3(n25548), .IN4(n252), .IN5(
        n2913), .Q(n2910) );
  OA22X1 U2849 ( .IN1(n25556), .IN2(n295), .IN3(n25564), .IN4(n338), .Q(n2913)
         );
  OA221X1 U2850 ( .IN1(n25508), .IN2(n381), .IN3(n25516), .IN4(n424), .IN5(
        n2914), .Q(n2909) );
  OA22X1 U2851 ( .IN1(n25524), .IN2(n467), .IN3(n25532), .IN4(n510), .Q(n2914)
         );
  OA221X1 U2852 ( .IN1(n25476), .IN2(n553), .IN3(n25484), .IN4(n596), .IN5(
        n2915), .Q(n2908) );
  OA22X1 U2853 ( .IN1(n25492), .IN2(n639), .IN3(n25500), .IN4(n682), .Q(n2915)
         );
  NAND4X0 U2854 ( .IN1(n2916), .IN2(n2917), .IN3(n2918), .IN4(n2919), .QN(
        n2906) );
  OA221X1 U2855 ( .IN1(n25444), .IN2(n37), .IN3(n25452), .IN4(n80), .IN5(n2920), .Q(n2919) );
  OA22X1 U2856 ( .IN1(n25460), .IN2(n123), .IN3(n25468), .IN4(n166), .Q(n2920)
         );
  OA221X1 U2857 ( .IN1(n25412), .IN2(n209), .IN3(n25420), .IN4(n252), .IN5(
        n2921), .Q(n2918) );
  OA22X1 U2858 ( .IN1(n25428), .IN2(n295), .IN3(n25436), .IN4(n338), .Q(n2921)
         );
  OA221X1 U2859 ( .IN1(n25380), .IN2(n381), .IN3(n25388), .IN4(n424), .IN5(
        n2922), .Q(n2917) );
  OA22X1 U2860 ( .IN1(n25396), .IN2(n467), .IN3(n25404), .IN4(n510), .Q(n2922)
         );
  OA221X1 U2861 ( .IN1(n25348), .IN2(n553), .IN3(n25356), .IN4(n596), .IN5(
        n2923), .Q(n2916) );
  OA22X1 U2862 ( .IN1(n25364), .IN2(n639), .IN3(n25372), .IN4(n682), .Q(n2923)
         );
  NAND4X0 U2863 ( .IN1(n2924), .IN2(n2925), .IN3(n2926), .IN4(n2927), .QN(
        n2904) );
  OA221X1 U2864 ( .IN1(n25316), .IN2(n37), .IN3(n25324), .IN4(n80), .IN5(n2928), .Q(n2927) );
  OA22X1 U2865 ( .IN1(n25332), .IN2(n123), .IN3(n25340), .IN4(n166), .Q(n2928)
         );
  OA221X1 U2866 ( .IN1(n25284), .IN2(n209), .IN3(n25292), .IN4(n252), .IN5(
        n2929), .Q(n2926) );
  OA22X1 U2867 ( .IN1(n25300), .IN2(n295), .IN3(n25308), .IN4(n338), .Q(n2929)
         );
  OA221X1 U2868 ( .IN1(n25252), .IN2(n381), .IN3(n25260), .IN4(n424), .IN5(
        n2930), .Q(n2925) );
  OA22X1 U2869 ( .IN1(n25268), .IN2(n467), .IN3(n25276), .IN4(n510), .Q(n2930)
         );
  OA221X1 U2870 ( .IN1(n25220), .IN2(n553), .IN3(n25228), .IN4(n596), .IN5(
        n2931), .Q(n2924) );
  OA22X1 U2871 ( .IN1(n25236), .IN2(n639), .IN3(n25244), .IN4(n682), .Q(n2931)
         );
  NAND4X0 U2872 ( .IN1(n2932), .IN2(n2933), .IN3(n2934), .IN4(n2935), .QN(
        n2903) );
  OA221X1 U2873 ( .IN1(n25188), .IN2(n37), .IN3(n25196), .IN4(n80), .IN5(n2936), .Q(n2935) );
  OA22X1 U2874 ( .IN1(n25204), .IN2(n123), .IN3(n25212), .IN4(n166), .Q(n2936)
         );
  OA221X1 U2875 ( .IN1(n25156), .IN2(n209), .IN3(n25164), .IN4(n252), .IN5(
        n2937), .Q(n2934) );
  OA22X1 U2876 ( .IN1(n25172), .IN2(n295), .IN3(n25180), .IN4(n338), .Q(n2937)
         );
  OA221X1 U2877 ( .IN1(n25124), .IN2(n381), .IN3(n25132), .IN4(n424), .IN5(
        n2938), .Q(n2933) );
  OA22X1 U2878 ( .IN1(n25140), .IN2(n467), .IN3(n25148), .IN4(n510), .Q(n2938)
         );
  OA221X1 U2879 ( .IN1(n25092), .IN2(n553), .IN3(n25100), .IN4(n596), .IN5(
        n2939), .Q(n2932) );
  OA22X1 U2880 ( .IN1(n25108), .IN2(n639), .IN3(n25116), .IN4(n682), .Q(n2939)
         );
  AO221X1 U2881 ( .IN1(n2328), .IN2(n2940), .IN3(n2330), .IN4(n2941), .IN5(
        n2942), .Q(n2825) );
  AO22X1 U2882 ( .IN1(n2333), .IN2(n2943), .IN3(n2335), .IN4(n2944), .Q(n2942)
         );
  NAND4X0 U2883 ( .IN1(n2945), .IN2(n2946), .IN3(n2947), .IN4(n2948), .QN(
        n2944) );
  OA221X1 U2884 ( .IN1(n25060), .IN2(n37), .IN3(n25068), .IN4(n80), .IN5(n2949), .Q(n2948) );
  OA22X1 U2885 ( .IN1(n25076), .IN2(n123), .IN3(n25084), .IN4(n166), .Q(n2949)
         );
  OA221X1 U2886 ( .IN1(n25028), .IN2(n209), .IN3(n25036), .IN4(n252), .IN5(
        n2950), .Q(n2947) );
  OA22X1 U2887 ( .IN1(n25044), .IN2(n295), .IN3(n25052), .IN4(n338), .Q(n2950)
         );
  OA221X1 U2888 ( .IN1(n24996), .IN2(n381), .IN3(n25004), .IN4(n424), .IN5(
        n2951), .Q(n2946) );
  OA22X1 U2889 ( .IN1(n25012), .IN2(n467), .IN3(n25020), .IN4(n510), .Q(n2951)
         );
  OA221X1 U2890 ( .IN1(n24964), .IN2(n553), .IN3(n24972), .IN4(n596), .IN5(
        n2952), .Q(n2945) );
  OA22X1 U2891 ( .IN1(n24980), .IN2(n639), .IN3(n24988), .IN4(n682), .Q(n2952)
         );
  NAND4X0 U2892 ( .IN1(n2953), .IN2(n2954), .IN3(n2955), .IN4(n2956), .QN(
        n2943) );
  OA221X1 U2893 ( .IN1(n24932), .IN2(n37), .IN3(n24940), .IN4(n80), .IN5(n2957), .Q(n2956) );
  OA22X1 U2894 ( .IN1(n24948), .IN2(n123), .IN3(n24956), .IN4(n166), .Q(n2957)
         );
  OA221X1 U2895 ( .IN1(n24900), .IN2(n209), .IN3(n24908), .IN4(n252), .IN5(
        n2958), .Q(n2955) );
  OA22X1 U2896 ( .IN1(n24916), .IN2(n295), .IN3(n24924), .IN4(n338), .Q(n2958)
         );
  OA221X1 U2897 ( .IN1(n24868), .IN2(n381), .IN3(n24876), .IN4(n424), .IN5(
        n2959), .Q(n2954) );
  OA22X1 U2898 ( .IN1(n24884), .IN2(n467), .IN3(n24892), .IN4(n510), .Q(n2959)
         );
  OA221X1 U2899 ( .IN1(n24836), .IN2(n553), .IN3(n24844), .IN4(n596), .IN5(
        n2960), .Q(n2953) );
  OA22X1 U2900 ( .IN1(n24852), .IN2(n639), .IN3(n24860), .IN4(n682), .Q(n2960)
         );
  NAND4X0 U2901 ( .IN1(n2961), .IN2(n2962), .IN3(n2963), .IN4(n2964), .QN(
        n2941) );
  OA221X1 U2902 ( .IN1(n24804), .IN2(n37), .IN3(n24812), .IN4(n80), .IN5(n2965), .Q(n2964) );
  OA22X1 U2903 ( .IN1(n24820), .IN2(n123), .IN3(n24828), .IN4(n166), .Q(n2965)
         );
  OA221X1 U2904 ( .IN1(n24772), .IN2(n209), .IN3(n24780), .IN4(n252), .IN5(
        n2966), .Q(n2963) );
  OA22X1 U2905 ( .IN1(n24788), .IN2(n295), .IN3(n24796), .IN4(n338), .Q(n2966)
         );
  OA221X1 U2906 ( .IN1(n24740), .IN2(n381), .IN3(n24748), .IN4(n424), .IN5(
        n2967), .Q(n2962) );
  OA22X1 U2907 ( .IN1(n24756), .IN2(n467), .IN3(n24764), .IN4(n510), .Q(n2967)
         );
  OA221X1 U2908 ( .IN1(n24708), .IN2(n553), .IN3(n24716), .IN4(n596), .IN5(
        n2968), .Q(n2961) );
  OA22X1 U2909 ( .IN1(n24724), .IN2(n639), .IN3(n24732), .IN4(n682), .Q(n2968)
         );
  NAND4X0 U2910 ( .IN1(n2969), .IN2(n2970), .IN3(n2971), .IN4(n2972), .QN(
        n2940) );
  OA221X1 U2911 ( .IN1(n24676), .IN2(n37), .IN3(n24684), .IN4(n80), .IN5(n2973), .Q(n2972) );
  OA22X1 U2912 ( .IN1(n24692), .IN2(n123), .IN3(n24700), .IN4(n166), .Q(n2973)
         );
  OA221X1 U2913 ( .IN1(n24644), .IN2(n209), .IN3(n24652), .IN4(n252), .IN5(
        n2974), .Q(n2971) );
  OA22X1 U2914 ( .IN1(n24660), .IN2(n295), .IN3(n24668), .IN4(n338), .Q(n2974)
         );
  OA221X1 U2915 ( .IN1(n24612), .IN2(n381), .IN3(n24620), .IN4(n424), .IN5(
        n2975), .Q(n2970) );
  OA22X1 U2916 ( .IN1(n24628), .IN2(n467), .IN3(n24636), .IN4(n510), .Q(n2975)
         );
  OA221X1 U2917 ( .IN1(n24580), .IN2(n553), .IN3(n24588), .IN4(n596), .IN5(
        n2976), .Q(n2969) );
  OA22X1 U2918 ( .IN1(n24596), .IN2(n639), .IN3(n24604), .IN4(n682), .Q(n2976)
         );
  OR4X1 U2919 ( .IN1(n2977), .IN2(n2978), .IN3(n2979), .IN4(n2980), .Q(n2198)
         );
  AO221X1 U2920 ( .IN1(n2157), .IN2(n2981), .IN3(n2159), .IN4(n2982), .IN5(
        n2983), .Q(n2980) );
  AO22X1 U2921 ( .IN1(n2162), .IN2(n2984), .IN3(n2164), .IN4(n2985), .Q(n2983)
         );
  NAND4X0 U2922 ( .IN1(n2986), .IN2(n2987), .IN3(n2988), .IN4(n2989), .QN(
        n2985) );
  OA221X1 U2923 ( .IN1(n24547), .IN2(n36), .IN3(n24555), .IN4(n79), .IN5(n2990), .Q(n2989) );
  OA22X1 U2924 ( .IN1(n24563), .IN2(n122), .IN3(n24571), .IN4(n165), .Q(n2990)
         );
  OA221X1 U2925 ( .IN1(n24515), .IN2(n208), .IN3(n24523), .IN4(n251), .IN5(
        n2991), .Q(n2988) );
  OA22X1 U2926 ( .IN1(n24531), .IN2(n294), .IN3(n24539), .IN4(n337), .Q(n2991)
         );
  OA221X1 U2927 ( .IN1(n24483), .IN2(n380), .IN3(n24491), .IN4(n423), .IN5(
        n2992), .Q(n2987) );
  OA22X1 U2928 ( .IN1(n24499), .IN2(n466), .IN3(n24507), .IN4(n509), .Q(n2992)
         );
  OA221X1 U2929 ( .IN1(n24451), .IN2(n552), .IN3(n24459), .IN4(n595), .IN5(
        n2993), .Q(n2986) );
  OA22X1 U2930 ( .IN1(n24467), .IN2(n638), .IN3(n24475), .IN4(n681), .Q(n2993)
         );
  NAND4X0 U2931 ( .IN1(n2994), .IN2(n2995), .IN3(n2996), .IN4(n2997), .QN(
        n2984) );
  OA221X1 U2932 ( .IN1(n24419), .IN2(n36), .IN3(n24427), .IN4(n79), .IN5(n2998), .Q(n2997) );
  OA22X1 U2933 ( .IN1(n24435), .IN2(n122), .IN3(n24443), .IN4(n165), .Q(n2998)
         );
  OA221X1 U2934 ( .IN1(n24387), .IN2(n208), .IN3(n24395), .IN4(n251), .IN5(
        n2999), .Q(n2996) );
  OA22X1 U2935 ( .IN1(n24403), .IN2(n294), .IN3(n24411), .IN4(n337), .Q(n2999)
         );
  OA221X1 U2936 ( .IN1(n24355), .IN2(n380), .IN3(n24363), .IN4(n423), .IN5(
        n3000), .Q(n2995) );
  OA22X1 U2937 ( .IN1(n24371), .IN2(n466), .IN3(n24379), .IN4(n509), .Q(n3000)
         );
  OA221X1 U2938 ( .IN1(n24323), .IN2(n552), .IN3(n24331), .IN4(n595), .IN5(
        n3001), .Q(n2994) );
  OA22X1 U2939 ( .IN1(n24339), .IN2(n638), .IN3(n24347), .IN4(n681), .Q(n3001)
         );
  NAND4X0 U2940 ( .IN1(n3002), .IN2(n3003), .IN3(n3004), .IN4(n3005), .QN(
        n2982) );
  OA221X1 U2941 ( .IN1(n24291), .IN2(n36), .IN3(n24299), .IN4(n79), .IN5(n3006), .Q(n3005) );
  OA22X1 U2942 ( .IN1(n24307), .IN2(n122), .IN3(n24315), .IN4(n165), .Q(n3006)
         );
  OA221X1 U2943 ( .IN1(n24259), .IN2(n208), .IN3(n24267), .IN4(n251), .IN5(
        n3007), .Q(n3004) );
  OA22X1 U2944 ( .IN1(n24275), .IN2(n294), .IN3(n24283), .IN4(n337), .Q(n3007)
         );
  OA221X1 U2945 ( .IN1(n24227), .IN2(n380), .IN3(n24235), .IN4(n423), .IN5(
        n3008), .Q(n3003) );
  OA22X1 U2946 ( .IN1(n24243), .IN2(n466), .IN3(n24251), .IN4(n509), .Q(n3008)
         );
  OA221X1 U2947 ( .IN1(n24195), .IN2(n552), .IN3(n24203), .IN4(n595), .IN5(
        n3009), .Q(n3002) );
  OA22X1 U2948 ( .IN1(n24211), .IN2(n638), .IN3(n24219), .IN4(n681), .Q(n3009)
         );
  NAND4X0 U2949 ( .IN1(n3010), .IN2(n3011), .IN3(n3012), .IN4(n3013), .QN(
        n2981) );
  OA221X1 U2950 ( .IN1(n24163), .IN2(n36), .IN3(n24171), .IN4(n79), .IN5(n3014), .Q(n3013) );
  OA22X1 U2951 ( .IN1(n24179), .IN2(n122), .IN3(n24187), .IN4(n165), .Q(n3014)
         );
  OA221X1 U2952 ( .IN1(n24131), .IN2(n208), .IN3(n24139), .IN4(n251), .IN5(
        n3015), .Q(n3012) );
  OA22X1 U2953 ( .IN1(n24147), .IN2(n294), .IN3(n24155), .IN4(n337), .Q(n3015)
         );
  OA221X1 U2954 ( .IN1(n24099), .IN2(n380), .IN3(n24107), .IN4(n423), .IN5(
        n3016), .Q(n3011) );
  OA22X1 U2955 ( .IN1(n24115), .IN2(n466), .IN3(n24123), .IN4(n509), .Q(n3016)
         );
  OA221X1 U2956 ( .IN1(n24067), .IN2(n552), .IN3(n24075), .IN4(n595), .IN5(
        n3017), .Q(n3010) );
  OA22X1 U2957 ( .IN1(n24083), .IN2(n638), .IN3(n24091), .IN4(n681), .Q(n3017)
         );
  AO221X1 U2958 ( .IN1(n2246), .IN2(n3018), .IN3(n2248), .IN4(n3019), .IN5(
        n3020), .Q(n2979) );
  AO22X1 U2959 ( .IN1(n2251), .IN2(n3021), .IN3(n2253), .IN4(n3022), .Q(n3020)
         );
  NAND4X0 U2960 ( .IN1(n3023), .IN2(n3024), .IN3(n3025), .IN4(n3026), .QN(
        n3022) );
  OA221X1 U2961 ( .IN1(n24035), .IN2(n36), .IN3(n24043), .IN4(n79), .IN5(n3027), .Q(n3026) );
  OA22X1 U2962 ( .IN1(n24051), .IN2(n122), .IN3(n24059), .IN4(n165), .Q(n3027)
         );
  OA221X1 U2963 ( .IN1(n24003), .IN2(n208), .IN3(n24011), .IN4(n251), .IN5(
        n3028), .Q(n3025) );
  OA22X1 U2964 ( .IN1(n24019), .IN2(n294), .IN3(n24027), .IN4(n337), .Q(n3028)
         );
  OA221X1 U2965 ( .IN1(n23971), .IN2(n380), .IN3(n23979), .IN4(n423), .IN5(
        n3029), .Q(n3024) );
  OA22X1 U2966 ( .IN1(n23987), .IN2(n466), .IN3(n23995), .IN4(n509), .Q(n3029)
         );
  OA221X1 U2967 ( .IN1(n23939), .IN2(n552), .IN3(n23947), .IN4(n595), .IN5(
        n3030), .Q(n3023) );
  OA22X1 U2968 ( .IN1(n23955), .IN2(n638), .IN3(n23963), .IN4(n681), .Q(n3030)
         );
  NAND4X0 U2969 ( .IN1(n3031), .IN2(n3032), .IN3(n3033), .IN4(n3034), .QN(
        n3021) );
  OA221X1 U2970 ( .IN1(n23907), .IN2(n36), .IN3(n23915), .IN4(n79), .IN5(n3035), .Q(n3034) );
  OA22X1 U2971 ( .IN1(n23923), .IN2(n122), .IN3(n23931), .IN4(n165), .Q(n3035)
         );
  OA221X1 U2972 ( .IN1(n23875), .IN2(n208), .IN3(n23883), .IN4(n251), .IN5(
        n3036), .Q(n3033) );
  OA22X1 U2973 ( .IN1(n23891), .IN2(n294), .IN3(n23899), .IN4(n337), .Q(n3036)
         );
  OA221X1 U2974 ( .IN1(n23843), .IN2(n380), .IN3(n23851), .IN4(n423), .IN5(
        n3037), .Q(n3032) );
  OA22X1 U2975 ( .IN1(n23859), .IN2(n466), .IN3(n23867), .IN4(n509), .Q(n3037)
         );
  OA221X1 U2976 ( .IN1(n23811), .IN2(n552), .IN3(n23819), .IN4(n595), .IN5(
        n3038), .Q(n3031) );
  OA22X1 U2977 ( .IN1(n23827), .IN2(n638), .IN3(n23835), .IN4(n681), .Q(n3038)
         );
  NAND4X0 U2978 ( .IN1(n3039), .IN2(n3040), .IN3(n3041), .IN4(n3042), .QN(
        n3019) );
  OA221X1 U2979 ( .IN1(n23779), .IN2(n36), .IN3(n23787), .IN4(n79), .IN5(n3043), .Q(n3042) );
  OA22X1 U2980 ( .IN1(n23795), .IN2(n122), .IN3(n23803), .IN4(n165), .Q(n3043)
         );
  OA221X1 U2981 ( .IN1(n23747), .IN2(n208), .IN3(n23755), .IN4(n251), .IN5(
        n3044), .Q(n3041) );
  OA22X1 U2982 ( .IN1(n23763), .IN2(n294), .IN3(n23771), .IN4(n337), .Q(n3044)
         );
  OA221X1 U2983 ( .IN1(n23715), .IN2(n380), .IN3(n23723), .IN4(n423), .IN5(
        n3045), .Q(n3040) );
  OA22X1 U2984 ( .IN1(n23731), .IN2(n466), .IN3(n23739), .IN4(n509), .Q(n3045)
         );
  OA221X1 U2985 ( .IN1(n23683), .IN2(n552), .IN3(n23691), .IN4(n595), .IN5(
        n3046), .Q(n3039) );
  OA22X1 U2986 ( .IN1(n23699), .IN2(n638), .IN3(n23707), .IN4(n681), .Q(n3046)
         );
  NAND4X0 U2987 ( .IN1(n3047), .IN2(n3048), .IN3(n3049), .IN4(n3050), .QN(
        n3018) );
  OA221X1 U2988 ( .IN1(n23651), .IN2(n36), .IN3(n23659), .IN4(n79), .IN5(n3051), .Q(n3050) );
  OA22X1 U2989 ( .IN1(n23667), .IN2(n122), .IN3(n23675), .IN4(n165), .Q(n3051)
         );
  OA221X1 U2990 ( .IN1(n23619), .IN2(n208), .IN3(n23627), .IN4(n251), .IN5(
        n3052), .Q(n3049) );
  OA22X1 U2991 ( .IN1(n23635), .IN2(n294), .IN3(n23643), .IN4(n337), .Q(n3052)
         );
  OA221X1 U2992 ( .IN1(n23587), .IN2(n380), .IN3(n23595), .IN4(n423), .IN5(
        n3053), .Q(n3048) );
  OA22X1 U2993 ( .IN1(n23603), .IN2(n466), .IN3(n23611), .IN4(n509), .Q(n3053)
         );
  OA221X1 U2994 ( .IN1(n23555), .IN2(n552), .IN3(n23563), .IN4(n595), .IN5(
        n3054), .Q(n3047) );
  OA22X1 U2995 ( .IN1(n23571), .IN2(n638), .IN3(n23579), .IN4(n681), .Q(n3054)
         );
  AO221X1 U2996 ( .IN1(n2287), .IN2(n3055), .IN3(n2289), .IN4(n3056), .IN5(
        n3057), .Q(n2978) );
  AO22X1 U2997 ( .IN1(n2292), .IN2(n3058), .IN3(n2294), .IN4(n3059), .Q(n3057)
         );
  NAND4X0 U2998 ( .IN1(n3060), .IN2(n3061), .IN3(n3062), .IN4(n3063), .QN(
        n3059) );
  OA221X1 U2999 ( .IN1(n25571), .IN2(n36), .IN3(n25579), .IN4(n79), .IN5(n3064), .Q(n3063) );
  OA22X1 U3000 ( .IN1(n25587), .IN2(n122), .IN3(n25595), .IN4(n165), .Q(n3064)
         );
  OA221X1 U3001 ( .IN1(n25539), .IN2(n208), .IN3(n25547), .IN4(n251), .IN5(
        n3065), .Q(n3062) );
  OA22X1 U3002 ( .IN1(n25555), .IN2(n294), .IN3(n25563), .IN4(n337), .Q(n3065)
         );
  OA221X1 U3003 ( .IN1(n25507), .IN2(n380), .IN3(n25515), .IN4(n423), .IN5(
        n3066), .Q(n3061) );
  OA22X1 U3004 ( .IN1(n25523), .IN2(n466), .IN3(n25531), .IN4(n509), .Q(n3066)
         );
  OA221X1 U3005 ( .IN1(n25475), .IN2(n552), .IN3(n25483), .IN4(n595), .IN5(
        n3067), .Q(n3060) );
  OA22X1 U3006 ( .IN1(n25491), .IN2(n638), .IN3(n25499), .IN4(n681), .Q(n3067)
         );
  NAND4X0 U3007 ( .IN1(n3068), .IN2(n3069), .IN3(n3070), .IN4(n3071), .QN(
        n3058) );
  OA221X1 U3008 ( .IN1(n25443), .IN2(n36), .IN3(n25451), .IN4(n79), .IN5(n3072), .Q(n3071) );
  OA22X1 U3009 ( .IN1(n25459), .IN2(n122), .IN3(n25467), .IN4(n165), .Q(n3072)
         );
  OA221X1 U3010 ( .IN1(n25411), .IN2(n208), .IN3(n25419), .IN4(n251), .IN5(
        n3073), .Q(n3070) );
  OA22X1 U3011 ( .IN1(n25427), .IN2(n294), .IN3(n25435), .IN4(n337), .Q(n3073)
         );
  OA221X1 U3012 ( .IN1(n25379), .IN2(n380), .IN3(n25387), .IN4(n423), .IN5(
        n3074), .Q(n3069) );
  OA22X1 U3013 ( .IN1(n25395), .IN2(n466), .IN3(n25403), .IN4(n509), .Q(n3074)
         );
  OA221X1 U3014 ( .IN1(n25347), .IN2(n552), .IN3(n25355), .IN4(n595), .IN5(
        n3075), .Q(n3068) );
  OA22X1 U3015 ( .IN1(n25363), .IN2(n638), .IN3(n25371), .IN4(n681), .Q(n3075)
         );
  NAND4X0 U3016 ( .IN1(n3076), .IN2(n3077), .IN3(n3078), .IN4(n3079), .QN(
        n3056) );
  OA221X1 U3017 ( .IN1(n25315), .IN2(n36), .IN3(n25323), .IN4(n79), .IN5(n3080), .Q(n3079) );
  OA22X1 U3018 ( .IN1(n25331), .IN2(n122), .IN3(n25339), .IN4(n165), .Q(n3080)
         );
  OA221X1 U3019 ( .IN1(n25283), .IN2(n208), .IN3(n25291), .IN4(n251), .IN5(
        n3081), .Q(n3078) );
  OA22X1 U3020 ( .IN1(n25299), .IN2(n294), .IN3(n25307), .IN4(n337), .Q(n3081)
         );
  OA221X1 U3021 ( .IN1(n25251), .IN2(n380), .IN3(n25259), .IN4(n423), .IN5(
        n3082), .Q(n3077) );
  OA22X1 U3022 ( .IN1(n25267), .IN2(n466), .IN3(n25275), .IN4(n509), .Q(n3082)
         );
  OA221X1 U3023 ( .IN1(n25219), .IN2(n552), .IN3(n25227), .IN4(n595), .IN5(
        n3083), .Q(n3076) );
  OA22X1 U3024 ( .IN1(n25235), .IN2(n638), .IN3(n25243), .IN4(n681), .Q(n3083)
         );
  NAND4X0 U3025 ( .IN1(n3084), .IN2(n3085), .IN3(n3086), .IN4(n3087), .QN(
        n3055) );
  OA221X1 U3026 ( .IN1(n25187), .IN2(n36), .IN3(n25195), .IN4(n79), .IN5(n3088), .Q(n3087) );
  OA22X1 U3027 ( .IN1(n25203), .IN2(n122), .IN3(n25211), .IN4(n165), .Q(n3088)
         );
  OA221X1 U3028 ( .IN1(n25155), .IN2(n208), .IN3(n25163), .IN4(n251), .IN5(
        n3089), .Q(n3086) );
  OA22X1 U3029 ( .IN1(n25171), .IN2(n294), .IN3(n25179), .IN4(n337), .Q(n3089)
         );
  OA221X1 U3030 ( .IN1(n25123), .IN2(n380), .IN3(n25131), .IN4(n423), .IN5(
        n3090), .Q(n3085) );
  OA22X1 U3031 ( .IN1(n25139), .IN2(n466), .IN3(n25147), .IN4(n509), .Q(n3090)
         );
  OA221X1 U3032 ( .IN1(n25091), .IN2(n552), .IN3(n25099), .IN4(n595), .IN5(
        n3091), .Q(n3084) );
  OA22X1 U3033 ( .IN1(n25107), .IN2(n638), .IN3(n25115), .IN4(n681), .Q(n3091)
         );
  AO221X1 U3034 ( .IN1(n2328), .IN2(n3092), .IN3(n2330), .IN4(n3093), .IN5(
        n3094), .Q(n2977) );
  AO22X1 U3035 ( .IN1(n2333), .IN2(n3095), .IN3(n2335), .IN4(n3096), .Q(n3094)
         );
  NAND4X0 U3036 ( .IN1(n3097), .IN2(n3098), .IN3(n3099), .IN4(n3100), .QN(
        n3096) );
  OA221X1 U3037 ( .IN1(n25059), .IN2(n35), .IN3(n25067), .IN4(n78), .IN5(n3101), .Q(n3100) );
  OA22X1 U3038 ( .IN1(n25075), .IN2(n121), .IN3(n25083), .IN4(n164), .Q(n3101)
         );
  OA221X1 U3039 ( .IN1(n25027), .IN2(n207), .IN3(n25035), .IN4(n250), .IN5(
        n3102), .Q(n3099) );
  OA22X1 U3040 ( .IN1(n25043), .IN2(n293), .IN3(n25051), .IN4(n336), .Q(n3102)
         );
  OA221X1 U3041 ( .IN1(n24995), .IN2(n379), .IN3(n25003), .IN4(n422), .IN5(
        n3103), .Q(n3098) );
  OA22X1 U3042 ( .IN1(n25011), .IN2(n465), .IN3(n25019), .IN4(n508), .Q(n3103)
         );
  OA221X1 U3043 ( .IN1(n24963), .IN2(n551), .IN3(n24971), .IN4(n594), .IN5(
        n3104), .Q(n3097) );
  OA22X1 U3044 ( .IN1(n24979), .IN2(n637), .IN3(n24987), .IN4(n680), .Q(n3104)
         );
  NAND4X0 U3045 ( .IN1(n3105), .IN2(n3106), .IN3(n3107), .IN4(n3108), .QN(
        n3095) );
  OA221X1 U3046 ( .IN1(n24931), .IN2(n35), .IN3(n24939), .IN4(n78), .IN5(n3109), .Q(n3108) );
  OA22X1 U3047 ( .IN1(n24947), .IN2(n121), .IN3(n24955), .IN4(n164), .Q(n3109)
         );
  OA221X1 U3048 ( .IN1(n24899), .IN2(n207), .IN3(n24907), .IN4(n250), .IN5(
        n3110), .Q(n3107) );
  OA22X1 U3049 ( .IN1(n24915), .IN2(n293), .IN3(n24923), .IN4(n336), .Q(n3110)
         );
  OA221X1 U3050 ( .IN1(n24867), .IN2(n379), .IN3(n24875), .IN4(n422), .IN5(
        n3111), .Q(n3106) );
  OA22X1 U3051 ( .IN1(n24883), .IN2(n465), .IN3(n24891), .IN4(n508), .Q(n3111)
         );
  OA221X1 U3052 ( .IN1(n24835), .IN2(n551), .IN3(n24843), .IN4(n594), .IN5(
        n3112), .Q(n3105) );
  OA22X1 U3053 ( .IN1(n24851), .IN2(n637), .IN3(n24859), .IN4(n680), .Q(n3112)
         );
  NAND4X0 U3054 ( .IN1(n3113), .IN2(n3114), .IN3(n3115), .IN4(n3116), .QN(
        n3093) );
  OA221X1 U3055 ( .IN1(n24803), .IN2(n35), .IN3(n24811), .IN4(n78), .IN5(n3117), .Q(n3116) );
  OA22X1 U3056 ( .IN1(n24819), .IN2(n121), .IN3(n24827), .IN4(n164), .Q(n3117)
         );
  OA221X1 U3057 ( .IN1(n24771), .IN2(n207), .IN3(n24779), .IN4(n250), .IN5(
        n3118), .Q(n3115) );
  OA22X1 U3058 ( .IN1(n24787), .IN2(n293), .IN3(n24795), .IN4(n336), .Q(n3118)
         );
  OA221X1 U3059 ( .IN1(n24739), .IN2(n379), .IN3(n24747), .IN4(n422), .IN5(
        n3119), .Q(n3114) );
  OA22X1 U3060 ( .IN1(n24755), .IN2(n465), .IN3(n24763), .IN4(n508), .Q(n3119)
         );
  OA221X1 U3061 ( .IN1(n24707), .IN2(n551), .IN3(n24715), .IN4(n594), .IN5(
        n3120), .Q(n3113) );
  OA22X1 U3062 ( .IN1(n24723), .IN2(n637), .IN3(n24731), .IN4(n680), .Q(n3120)
         );
  NAND4X0 U3063 ( .IN1(n3121), .IN2(n3122), .IN3(n3123), .IN4(n3124), .QN(
        n3092) );
  OA221X1 U3064 ( .IN1(n24675), .IN2(n35), .IN3(n24683), .IN4(n78), .IN5(n3125), .Q(n3124) );
  OA22X1 U3065 ( .IN1(n24691), .IN2(n121), .IN3(n24699), .IN4(n164), .Q(n3125)
         );
  OA221X1 U3066 ( .IN1(n24643), .IN2(n207), .IN3(n24651), .IN4(n250), .IN5(
        n3126), .Q(n3123) );
  OA22X1 U3067 ( .IN1(n24659), .IN2(n293), .IN3(n24667), .IN4(n336), .Q(n3126)
         );
  OA221X1 U3068 ( .IN1(n24611), .IN2(n379), .IN3(n24619), .IN4(n422), .IN5(
        n3127), .Q(n3122) );
  OA22X1 U3069 ( .IN1(n24627), .IN2(n465), .IN3(n24635), .IN4(n508), .Q(n3127)
         );
  OA221X1 U3070 ( .IN1(n24579), .IN2(n551), .IN3(n24587), .IN4(n594), .IN5(
        n3128), .Q(n3121) );
  OA22X1 U3071 ( .IN1(n24595), .IN2(n637), .IN3(n24603), .IN4(n680), .Q(n3128)
         );
  OR4X1 U3072 ( .IN1(n3129), .IN2(n3130), .IN3(n3131), .IN4(n3132), .Q(n2197)
         );
  AO221X1 U3073 ( .IN1(n2157), .IN2(n3133), .IN3(n2159), .IN4(n3134), .IN5(
        n3135), .Q(n3132) );
  AO22X1 U3074 ( .IN1(n2162), .IN2(n3136), .IN3(n2164), .IN4(n3137), .Q(n3135)
         );
  NAND4X0 U3075 ( .IN1(n3138), .IN2(n3139), .IN3(n3140), .IN4(n3141), .QN(
        n3137) );
  OA221X1 U3076 ( .IN1(n24546), .IN2(n35), .IN3(n24554), .IN4(n78), .IN5(n3142), .Q(n3141) );
  OA22X1 U3077 ( .IN1(n24562), .IN2(n121), .IN3(n24570), .IN4(n164), .Q(n3142)
         );
  OA221X1 U3078 ( .IN1(n24514), .IN2(n207), .IN3(n24522), .IN4(n250), .IN5(
        n3143), .Q(n3140) );
  OA22X1 U3079 ( .IN1(n24530), .IN2(n293), .IN3(n24538), .IN4(n336), .Q(n3143)
         );
  OA221X1 U3080 ( .IN1(n24482), .IN2(n379), .IN3(n24490), .IN4(n422), .IN5(
        n3144), .Q(n3139) );
  OA22X1 U3081 ( .IN1(n24498), .IN2(n465), .IN3(n24506), .IN4(n508), .Q(n3144)
         );
  OA221X1 U3082 ( .IN1(n24450), .IN2(n551), .IN3(n24458), .IN4(n594), .IN5(
        n3145), .Q(n3138) );
  OA22X1 U3083 ( .IN1(n24466), .IN2(n637), .IN3(n24474), .IN4(n680), .Q(n3145)
         );
  NAND4X0 U3084 ( .IN1(n3146), .IN2(n3147), .IN3(n3148), .IN4(n3149), .QN(
        n3136) );
  OA221X1 U3085 ( .IN1(n24418), .IN2(n35), .IN3(n24426), .IN4(n78), .IN5(n3150), .Q(n3149) );
  OA22X1 U3086 ( .IN1(n24434), .IN2(n121), .IN3(n24442), .IN4(n164), .Q(n3150)
         );
  OA221X1 U3087 ( .IN1(n24386), .IN2(n207), .IN3(n24394), .IN4(n250), .IN5(
        n3151), .Q(n3148) );
  OA22X1 U3088 ( .IN1(n24402), .IN2(n293), .IN3(n24410), .IN4(n336), .Q(n3151)
         );
  OA221X1 U3089 ( .IN1(n24354), .IN2(n379), .IN3(n24362), .IN4(n422), .IN5(
        n3152), .Q(n3147) );
  OA22X1 U3090 ( .IN1(n24370), .IN2(n465), .IN3(n24378), .IN4(n508), .Q(n3152)
         );
  OA221X1 U3091 ( .IN1(n24322), .IN2(n551), .IN3(n24330), .IN4(n594), .IN5(
        n3153), .Q(n3146) );
  OA22X1 U3092 ( .IN1(n24338), .IN2(n637), .IN3(n24346), .IN4(n680), .Q(n3153)
         );
  NAND4X0 U3093 ( .IN1(n3154), .IN2(n3155), .IN3(n3156), .IN4(n3157), .QN(
        n3134) );
  OA221X1 U3094 ( .IN1(n24290), .IN2(n35), .IN3(n24298), .IN4(n78), .IN5(n3158), .Q(n3157) );
  OA22X1 U3095 ( .IN1(n24306), .IN2(n121), .IN3(n24314), .IN4(n164), .Q(n3158)
         );
  OA221X1 U3096 ( .IN1(n24258), .IN2(n207), .IN3(n24266), .IN4(n250), .IN5(
        n3159), .Q(n3156) );
  OA22X1 U3097 ( .IN1(n24274), .IN2(n293), .IN3(n24282), .IN4(n336), .Q(n3159)
         );
  OA221X1 U3098 ( .IN1(n24226), .IN2(n379), .IN3(n24234), .IN4(n422), .IN5(
        n3160), .Q(n3155) );
  OA22X1 U3099 ( .IN1(n24242), .IN2(n465), .IN3(n24250), .IN4(n508), .Q(n3160)
         );
  OA221X1 U3100 ( .IN1(n24194), .IN2(n551), .IN3(n24202), .IN4(n594), .IN5(
        n3161), .Q(n3154) );
  OA22X1 U3101 ( .IN1(n24210), .IN2(n637), .IN3(n24218), .IN4(n680), .Q(n3161)
         );
  NAND4X0 U3102 ( .IN1(n3162), .IN2(n3163), .IN3(n3164), .IN4(n3165), .QN(
        n3133) );
  OA221X1 U3103 ( .IN1(n24162), .IN2(n35), .IN3(n24170), .IN4(n78), .IN5(n3166), .Q(n3165) );
  OA22X1 U3104 ( .IN1(n24178), .IN2(n121), .IN3(n24186), .IN4(n164), .Q(n3166)
         );
  OA221X1 U3105 ( .IN1(n24130), .IN2(n207), .IN3(n24138), .IN4(n250), .IN5(
        n3167), .Q(n3164) );
  OA22X1 U3106 ( .IN1(n24146), .IN2(n293), .IN3(n24154), .IN4(n336), .Q(n3167)
         );
  OA221X1 U3107 ( .IN1(n24098), .IN2(n379), .IN3(n24106), .IN4(n422), .IN5(
        n3168), .Q(n3163) );
  OA22X1 U3108 ( .IN1(n24114), .IN2(n465), .IN3(n24122), .IN4(n508), .Q(n3168)
         );
  OA221X1 U3109 ( .IN1(n24066), .IN2(n551), .IN3(n24074), .IN4(n594), .IN5(
        n3169), .Q(n3162) );
  OA22X1 U3110 ( .IN1(n24082), .IN2(n637), .IN3(n24090), .IN4(n680), .Q(n3169)
         );
  AO221X1 U3111 ( .IN1(n2246), .IN2(n3170), .IN3(n2248), .IN4(n3171), .IN5(
        n3172), .Q(n3131) );
  AO22X1 U3112 ( .IN1(n2251), .IN2(n3173), .IN3(n2253), .IN4(n3174), .Q(n3172)
         );
  NAND4X0 U3113 ( .IN1(n3175), .IN2(n3176), .IN3(n3177), .IN4(n3178), .QN(
        n3174) );
  OA221X1 U3114 ( .IN1(n24034), .IN2(n35), .IN3(n24042), .IN4(n78), .IN5(n3179), .Q(n3178) );
  OA22X1 U3115 ( .IN1(n24050), .IN2(n121), .IN3(n24058), .IN4(n164), .Q(n3179)
         );
  OA221X1 U3116 ( .IN1(n24002), .IN2(n207), .IN3(n24010), .IN4(n250), .IN5(
        n3180), .Q(n3177) );
  OA22X1 U3117 ( .IN1(n24018), .IN2(n293), .IN3(n24026), .IN4(n336), .Q(n3180)
         );
  OA221X1 U3118 ( .IN1(n23970), .IN2(n379), .IN3(n23978), .IN4(n422), .IN5(
        n3181), .Q(n3176) );
  OA22X1 U3119 ( .IN1(n23986), .IN2(n465), .IN3(n23994), .IN4(n508), .Q(n3181)
         );
  OA221X1 U3120 ( .IN1(n23938), .IN2(n551), .IN3(n23946), .IN4(n594), .IN5(
        n3182), .Q(n3175) );
  OA22X1 U3121 ( .IN1(n23954), .IN2(n637), .IN3(n23962), .IN4(n680), .Q(n3182)
         );
  NAND4X0 U3122 ( .IN1(n3183), .IN2(n3184), .IN3(n3185), .IN4(n3186), .QN(
        n3173) );
  OA221X1 U3123 ( .IN1(n23906), .IN2(n35), .IN3(n23914), .IN4(n78), .IN5(n3187), .Q(n3186) );
  OA22X1 U3124 ( .IN1(n23922), .IN2(n121), .IN3(n23930), .IN4(n164), .Q(n3187)
         );
  OA221X1 U3125 ( .IN1(n23874), .IN2(n207), .IN3(n23882), .IN4(n250), .IN5(
        n3188), .Q(n3185) );
  OA22X1 U3126 ( .IN1(n23890), .IN2(n293), .IN3(n23898), .IN4(n336), .Q(n3188)
         );
  OA221X1 U3127 ( .IN1(n23842), .IN2(n379), .IN3(n23850), .IN4(n422), .IN5(
        n3189), .Q(n3184) );
  OA22X1 U3128 ( .IN1(n23858), .IN2(n465), .IN3(n23866), .IN4(n508), .Q(n3189)
         );
  OA221X1 U3129 ( .IN1(n23810), .IN2(n551), .IN3(n23818), .IN4(n594), .IN5(
        n3190), .Q(n3183) );
  OA22X1 U3130 ( .IN1(n23826), .IN2(n637), .IN3(n23834), .IN4(n680), .Q(n3190)
         );
  NAND4X0 U3131 ( .IN1(n3191), .IN2(n3192), .IN3(n3193), .IN4(n3194), .QN(
        n3171) );
  OA221X1 U3132 ( .IN1(n23778), .IN2(n35), .IN3(n23786), .IN4(n78), .IN5(n3195), .Q(n3194) );
  OA22X1 U3133 ( .IN1(n23794), .IN2(n121), .IN3(n23802), .IN4(n164), .Q(n3195)
         );
  OA221X1 U3134 ( .IN1(n23746), .IN2(n207), .IN3(n23754), .IN4(n250), .IN5(
        n3196), .Q(n3193) );
  OA22X1 U3135 ( .IN1(n23762), .IN2(n293), .IN3(n23770), .IN4(n336), .Q(n3196)
         );
  OA221X1 U3136 ( .IN1(n23714), .IN2(n379), .IN3(n23722), .IN4(n422), .IN5(
        n3197), .Q(n3192) );
  OA22X1 U3137 ( .IN1(n23730), .IN2(n465), .IN3(n23738), .IN4(n508), .Q(n3197)
         );
  OA221X1 U3138 ( .IN1(n23682), .IN2(n551), .IN3(n23690), .IN4(n594), .IN5(
        n3198), .Q(n3191) );
  OA22X1 U3139 ( .IN1(n23698), .IN2(n637), .IN3(n23706), .IN4(n680), .Q(n3198)
         );
  NAND4X0 U3140 ( .IN1(n3199), .IN2(n3200), .IN3(n3201), .IN4(n3202), .QN(
        n3170) );
  OA221X1 U3141 ( .IN1(n23650), .IN2(n35), .IN3(n23658), .IN4(n78), .IN5(n3203), .Q(n3202) );
  OA22X1 U3142 ( .IN1(n23666), .IN2(n121), .IN3(n23674), .IN4(n164), .Q(n3203)
         );
  OA221X1 U3143 ( .IN1(n23618), .IN2(n207), .IN3(n23626), .IN4(n250), .IN5(
        n3204), .Q(n3201) );
  OA22X1 U3144 ( .IN1(n23634), .IN2(n293), .IN3(n23642), .IN4(n336), .Q(n3204)
         );
  OA221X1 U3145 ( .IN1(n23586), .IN2(n379), .IN3(n23594), .IN4(n422), .IN5(
        n3205), .Q(n3200) );
  OA22X1 U3146 ( .IN1(n23602), .IN2(n465), .IN3(n23610), .IN4(n508), .Q(n3205)
         );
  OA221X1 U3147 ( .IN1(n23554), .IN2(n551), .IN3(n23562), .IN4(n594), .IN5(
        n3206), .Q(n3199) );
  OA22X1 U3148 ( .IN1(n23570), .IN2(n637), .IN3(n23578), .IN4(n680), .Q(n3206)
         );
  AO221X1 U3149 ( .IN1(n2287), .IN2(n3207), .IN3(n2289), .IN4(n3208), .IN5(
        n3209), .Q(n3130) );
  AO22X1 U3150 ( .IN1(n2292), .IN2(n3210), .IN3(n2294), .IN4(n3211), .Q(n3209)
         );
  NAND4X0 U3151 ( .IN1(n3212), .IN2(n3213), .IN3(n3214), .IN4(n3215), .QN(
        n3211) );
  OA221X1 U3152 ( .IN1(n25570), .IN2(n34), .IN3(n25578), .IN4(n77), .IN5(n3216), .Q(n3215) );
  OA22X1 U3153 ( .IN1(n25586), .IN2(n120), .IN3(n25594), .IN4(n163), .Q(n3216)
         );
  OA221X1 U3154 ( .IN1(n25538), .IN2(n206), .IN3(n25546), .IN4(n249), .IN5(
        n3217), .Q(n3214) );
  OA22X1 U3155 ( .IN1(n25554), .IN2(n292), .IN3(n25562), .IN4(n335), .Q(n3217)
         );
  OA221X1 U3156 ( .IN1(n25506), .IN2(n378), .IN3(n25514), .IN4(n421), .IN5(
        n3218), .Q(n3213) );
  OA22X1 U3157 ( .IN1(n25522), .IN2(n464), .IN3(n25530), .IN4(n507), .Q(n3218)
         );
  OA221X1 U3158 ( .IN1(n25474), .IN2(n550), .IN3(n25482), .IN4(n593), .IN5(
        n3219), .Q(n3212) );
  OA22X1 U3159 ( .IN1(n25490), .IN2(n636), .IN3(n25498), .IN4(n679), .Q(n3219)
         );
  NAND4X0 U3160 ( .IN1(n3220), .IN2(n3221), .IN3(n3222), .IN4(n3223), .QN(
        n3210) );
  OA221X1 U3161 ( .IN1(n25442), .IN2(n34), .IN3(n25450), .IN4(n77), .IN5(n3224), .Q(n3223) );
  OA22X1 U3162 ( .IN1(n25458), .IN2(n120), .IN3(n25466), .IN4(n163), .Q(n3224)
         );
  OA221X1 U3163 ( .IN1(n25410), .IN2(n206), .IN3(n25418), .IN4(n249), .IN5(
        n3225), .Q(n3222) );
  OA22X1 U3164 ( .IN1(n25426), .IN2(n292), .IN3(n25434), .IN4(n335), .Q(n3225)
         );
  OA221X1 U3165 ( .IN1(n25378), .IN2(n378), .IN3(n25386), .IN4(n421), .IN5(
        n3226), .Q(n3221) );
  OA22X1 U3166 ( .IN1(n25394), .IN2(n464), .IN3(n25402), .IN4(n507), .Q(n3226)
         );
  OA221X1 U3167 ( .IN1(n25346), .IN2(n550), .IN3(n25354), .IN4(n593), .IN5(
        n3227), .Q(n3220) );
  OA22X1 U3168 ( .IN1(n25362), .IN2(n636), .IN3(n25370), .IN4(n679), .Q(n3227)
         );
  NAND4X0 U3169 ( .IN1(n3228), .IN2(n3229), .IN3(n3230), .IN4(n3231), .QN(
        n3208) );
  OA221X1 U3170 ( .IN1(n25314), .IN2(n34), .IN3(n25322), .IN4(n77), .IN5(n3232), .Q(n3231) );
  OA22X1 U3171 ( .IN1(n25330), .IN2(n120), .IN3(n25338), .IN4(n163), .Q(n3232)
         );
  OA221X1 U3172 ( .IN1(n25282), .IN2(n206), .IN3(n25290), .IN4(n249), .IN5(
        n3233), .Q(n3230) );
  OA22X1 U3173 ( .IN1(n25298), .IN2(n292), .IN3(n25306), .IN4(n335), .Q(n3233)
         );
  OA221X1 U3174 ( .IN1(n25250), .IN2(n378), .IN3(n25258), .IN4(n421), .IN5(
        n3234), .Q(n3229) );
  OA22X1 U3175 ( .IN1(n25266), .IN2(n464), .IN3(n25274), .IN4(n507), .Q(n3234)
         );
  OA221X1 U3176 ( .IN1(n25218), .IN2(n550), .IN3(n25226), .IN4(n593), .IN5(
        n3235), .Q(n3228) );
  OA22X1 U3177 ( .IN1(n25234), .IN2(n636), .IN3(n25242), .IN4(n679), .Q(n3235)
         );
  NAND4X0 U3178 ( .IN1(n3236), .IN2(n3237), .IN3(n3238), .IN4(n3239), .QN(
        n3207) );
  OA221X1 U3179 ( .IN1(n25186), .IN2(n34), .IN3(n25194), .IN4(n77), .IN5(n3240), .Q(n3239) );
  OA22X1 U3180 ( .IN1(n25202), .IN2(n120), .IN3(n25210), .IN4(n163), .Q(n3240)
         );
  OA221X1 U3181 ( .IN1(n25154), .IN2(n206), .IN3(n25162), .IN4(n249), .IN5(
        n3241), .Q(n3238) );
  OA22X1 U3182 ( .IN1(n25170), .IN2(n292), .IN3(n25178), .IN4(n335), .Q(n3241)
         );
  OA221X1 U3183 ( .IN1(n25122), .IN2(n378), .IN3(n25130), .IN4(n421), .IN5(
        n3242), .Q(n3237) );
  OA22X1 U3184 ( .IN1(n25138), .IN2(n464), .IN3(n25146), .IN4(n507), .Q(n3242)
         );
  OA221X1 U3185 ( .IN1(n25090), .IN2(n550), .IN3(n25098), .IN4(n593), .IN5(
        n3243), .Q(n3236) );
  OA22X1 U3186 ( .IN1(n25106), .IN2(n636), .IN3(n25114), .IN4(n679), .Q(n3243)
         );
  AO221X1 U3187 ( .IN1(n2328), .IN2(n3244), .IN3(n2330), .IN4(n3245), .IN5(
        n3246), .Q(n3129) );
  AO22X1 U3188 ( .IN1(n2333), .IN2(n3247), .IN3(n2335), .IN4(n3248), .Q(n3246)
         );
  NAND4X0 U3189 ( .IN1(n3249), .IN2(n3250), .IN3(n3251), .IN4(n3252), .QN(
        n3248) );
  OA221X1 U3190 ( .IN1(n25058), .IN2(n34), .IN3(n25066), .IN4(n77), .IN5(n3253), .Q(n3252) );
  OA22X1 U3191 ( .IN1(n25074), .IN2(n120), .IN3(n25082), .IN4(n163), .Q(n3253)
         );
  OA221X1 U3192 ( .IN1(n25026), .IN2(n206), .IN3(n25034), .IN4(n249), .IN5(
        n3254), .Q(n3251) );
  OA22X1 U3193 ( .IN1(n25042), .IN2(n292), .IN3(n25050), .IN4(n335), .Q(n3254)
         );
  OA221X1 U3194 ( .IN1(n24994), .IN2(n378), .IN3(n25002), .IN4(n421), .IN5(
        n3255), .Q(n3250) );
  OA22X1 U3195 ( .IN1(n25010), .IN2(n464), .IN3(n25018), .IN4(n507), .Q(n3255)
         );
  OA221X1 U3196 ( .IN1(n24962), .IN2(n550), .IN3(n24970), .IN4(n593), .IN5(
        n3256), .Q(n3249) );
  OA22X1 U3197 ( .IN1(n24978), .IN2(n636), .IN3(n24986), .IN4(n679), .Q(n3256)
         );
  NAND4X0 U3198 ( .IN1(n3257), .IN2(n3258), .IN3(n3259), .IN4(n3260), .QN(
        n3247) );
  OA221X1 U3199 ( .IN1(n24930), .IN2(n34), .IN3(n24938), .IN4(n77), .IN5(n3261), .Q(n3260) );
  OA22X1 U3200 ( .IN1(n24946), .IN2(n120), .IN3(n24954), .IN4(n163), .Q(n3261)
         );
  OA221X1 U3201 ( .IN1(n24898), .IN2(n206), .IN3(n24906), .IN4(n249), .IN5(
        n3262), .Q(n3259) );
  OA22X1 U3202 ( .IN1(n24914), .IN2(n292), .IN3(n24922), .IN4(n335), .Q(n3262)
         );
  OA221X1 U3203 ( .IN1(n24866), .IN2(n378), .IN3(n24874), .IN4(n421), .IN5(
        n3263), .Q(n3258) );
  OA22X1 U3204 ( .IN1(n24882), .IN2(n464), .IN3(n24890), .IN4(n507), .Q(n3263)
         );
  OA221X1 U3205 ( .IN1(n24834), .IN2(n550), .IN3(n24842), .IN4(n593), .IN5(
        n3264), .Q(n3257) );
  OA22X1 U3206 ( .IN1(n24850), .IN2(n636), .IN3(n24858), .IN4(n679), .Q(n3264)
         );
  NAND4X0 U3207 ( .IN1(n3265), .IN2(n3266), .IN3(n3267), .IN4(n3268), .QN(
        n3245) );
  OA221X1 U3208 ( .IN1(n24802), .IN2(n34), .IN3(n24810), .IN4(n77), .IN5(n3269), .Q(n3268) );
  OA22X1 U3209 ( .IN1(n24818), .IN2(n120), .IN3(n24826), .IN4(n163), .Q(n3269)
         );
  OA221X1 U3210 ( .IN1(n24770), .IN2(n206), .IN3(n24778), .IN4(n249), .IN5(
        n3270), .Q(n3267) );
  OA22X1 U3211 ( .IN1(n24786), .IN2(n292), .IN3(n24794), .IN4(n335), .Q(n3270)
         );
  OA221X1 U3212 ( .IN1(n24738), .IN2(n378), .IN3(n24746), .IN4(n421), .IN5(
        n3271), .Q(n3266) );
  OA22X1 U3213 ( .IN1(n24754), .IN2(n464), .IN3(n24762), .IN4(n507), .Q(n3271)
         );
  OA221X1 U3214 ( .IN1(n24706), .IN2(n550), .IN3(n24714), .IN4(n593), .IN5(
        n3272), .Q(n3265) );
  OA22X1 U3215 ( .IN1(n24722), .IN2(n636), .IN3(n24730), .IN4(n679), .Q(n3272)
         );
  NAND4X0 U3216 ( .IN1(n3273), .IN2(n3274), .IN3(n3275), .IN4(n3276), .QN(
        n3244) );
  OA221X1 U3217 ( .IN1(n24674), .IN2(n34), .IN3(n24682), .IN4(n77), .IN5(n3277), .Q(n3276) );
  OA22X1 U3218 ( .IN1(n24690), .IN2(n120), .IN3(n24698), .IN4(n163), .Q(n3277)
         );
  OA221X1 U3219 ( .IN1(n24642), .IN2(n206), .IN3(n24650), .IN4(n249), .IN5(
        n3278), .Q(n3275) );
  OA22X1 U3220 ( .IN1(n24658), .IN2(n292), .IN3(n24666), .IN4(n335), .Q(n3278)
         );
  OA221X1 U3221 ( .IN1(n24610), .IN2(n378), .IN3(n24618), .IN4(n421), .IN5(
        n3279), .Q(n3274) );
  OA22X1 U3222 ( .IN1(n24626), .IN2(n464), .IN3(n24634), .IN4(n507), .Q(n3279)
         );
  OA221X1 U3223 ( .IN1(n24578), .IN2(n550), .IN3(n24586), .IN4(n593), .IN5(
        n3280), .Q(n3273) );
  OA22X1 U3224 ( .IN1(n24594), .IN2(n636), .IN3(n24602), .IN4(n679), .Q(n3280)
         );
  OR4X1 U3225 ( .IN1(n3281), .IN2(n3282), .IN3(n3283), .IN4(n3284), .Q(n2196)
         );
  AO221X1 U3226 ( .IN1(n2157), .IN2(n3285), .IN3(n2159), .IN4(n3286), .IN5(
        n3287), .Q(n3284) );
  AO22X1 U3227 ( .IN1(n2162), .IN2(n3288), .IN3(n2164), .IN4(n3289), .Q(n3287)
         );
  NAND4X0 U3228 ( .IN1(n3290), .IN2(n3291), .IN3(n3292), .IN4(n3293), .QN(
        n3289) );
  OA221X1 U3229 ( .IN1(n24545), .IN2(n34), .IN3(n24553), .IN4(n77), .IN5(n3294), .Q(n3293) );
  OA22X1 U3230 ( .IN1(n24561), .IN2(n120), .IN3(n24569), .IN4(n163), .Q(n3294)
         );
  OA221X1 U3231 ( .IN1(n24513), .IN2(n206), .IN3(n24521), .IN4(n249), .IN5(
        n3295), .Q(n3292) );
  OA22X1 U3232 ( .IN1(n24529), .IN2(n292), .IN3(n24537), .IN4(n335), .Q(n3295)
         );
  OA221X1 U3233 ( .IN1(n24481), .IN2(n378), .IN3(n24489), .IN4(n421), .IN5(
        n3296), .Q(n3291) );
  OA22X1 U3234 ( .IN1(n24497), .IN2(n464), .IN3(n24505), .IN4(n507), .Q(n3296)
         );
  OA221X1 U3235 ( .IN1(n24449), .IN2(n550), .IN3(n24457), .IN4(n593), .IN5(
        n3297), .Q(n3290) );
  OA22X1 U3236 ( .IN1(n24465), .IN2(n636), .IN3(n24473), .IN4(n679), .Q(n3297)
         );
  NAND4X0 U3237 ( .IN1(n3298), .IN2(n3299), .IN3(n3300), .IN4(n3301), .QN(
        n3288) );
  OA221X1 U3238 ( .IN1(n24417), .IN2(n34), .IN3(n24425), .IN4(n77), .IN5(n3302), .Q(n3301) );
  OA22X1 U3239 ( .IN1(n24433), .IN2(n120), .IN3(n24441), .IN4(n163), .Q(n3302)
         );
  OA221X1 U3240 ( .IN1(n24385), .IN2(n206), .IN3(n24393), .IN4(n249), .IN5(
        n3303), .Q(n3300) );
  OA22X1 U3241 ( .IN1(n24401), .IN2(n292), .IN3(n24409), .IN4(n335), .Q(n3303)
         );
  OA221X1 U3242 ( .IN1(n24353), .IN2(n378), .IN3(n24361), .IN4(n421), .IN5(
        n3304), .Q(n3299) );
  OA22X1 U3243 ( .IN1(n24369), .IN2(n464), .IN3(n24377), .IN4(n507), .Q(n3304)
         );
  OA221X1 U3244 ( .IN1(n24321), .IN2(n550), .IN3(n24329), .IN4(n593), .IN5(
        n3305), .Q(n3298) );
  OA22X1 U3245 ( .IN1(n24337), .IN2(n636), .IN3(n24345), .IN4(n679), .Q(n3305)
         );
  NAND4X0 U3246 ( .IN1(n3306), .IN2(n3307), .IN3(n3308), .IN4(n3309), .QN(
        n3286) );
  OA221X1 U3247 ( .IN1(n24289), .IN2(n34), .IN3(n24297), .IN4(n77), .IN5(n3310), .Q(n3309) );
  OA22X1 U3248 ( .IN1(n24305), .IN2(n120), .IN3(n24313), .IN4(n163), .Q(n3310)
         );
  OA221X1 U3249 ( .IN1(n24257), .IN2(n206), .IN3(n24265), .IN4(n249), .IN5(
        n3311), .Q(n3308) );
  OA22X1 U3250 ( .IN1(n24273), .IN2(n292), .IN3(n24281), .IN4(n335), .Q(n3311)
         );
  OA221X1 U3251 ( .IN1(n24225), .IN2(n378), .IN3(n24233), .IN4(n421), .IN5(
        n3312), .Q(n3307) );
  OA22X1 U3252 ( .IN1(n24241), .IN2(n464), .IN3(n24249), .IN4(n507), .Q(n3312)
         );
  OA221X1 U3253 ( .IN1(n24193), .IN2(n550), .IN3(n24201), .IN4(n593), .IN5(
        n3313), .Q(n3306) );
  OA22X1 U3254 ( .IN1(n24209), .IN2(n636), .IN3(n24217), .IN4(n679), .Q(n3313)
         );
  NAND4X0 U3255 ( .IN1(n3314), .IN2(n3315), .IN3(n3316), .IN4(n3317), .QN(
        n3285) );
  OA221X1 U3256 ( .IN1(n24161), .IN2(n34), .IN3(n24169), .IN4(n77), .IN5(n3318), .Q(n3317) );
  OA22X1 U3257 ( .IN1(n24177), .IN2(n120), .IN3(n24185), .IN4(n163), .Q(n3318)
         );
  OA221X1 U3258 ( .IN1(n24129), .IN2(n206), .IN3(n24137), .IN4(n249), .IN5(
        n3319), .Q(n3316) );
  OA22X1 U3259 ( .IN1(n24145), .IN2(n292), .IN3(n24153), .IN4(n335), .Q(n3319)
         );
  OA221X1 U3260 ( .IN1(n24097), .IN2(n378), .IN3(n24105), .IN4(n421), .IN5(
        n3320), .Q(n3315) );
  OA22X1 U3261 ( .IN1(n24113), .IN2(n464), .IN3(n24121), .IN4(n507), .Q(n3320)
         );
  OA221X1 U3262 ( .IN1(n24065), .IN2(n550), .IN3(n24073), .IN4(n593), .IN5(
        n3321), .Q(n3314) );
  OA22X1 U3263 ( .IN1(n24081), .IN2(n636), .IN3(n24089), .IN4(n679), .Q(n3321)
         );
  AO221X1 U3264 ( .IN1(n2246), .IN2(n3322), .IN3(n2248), .IN4(n3323), .IN5(
        n3324), .Q(n3283) );
  AO22X1 U3265 ( .IN1(n2251), .IN2(n3325), .IN3(n2253), .IN4(n3326), .Q(n3324)
         );
  NAND4X0 U3266 ( .IN1(n3327), .IN2(n3328), .IN3(n3329), .IN4(n3330), .QN(
        n3326) );
  OA221X1 U3267 ( .IN1(n24033), .IN2(n33), .IN3(n24041), .IN4(n76), .IN5(n3331), .Q(n3330) );
  OA22X1 U3268 ( .IN1(n24049), .IN2(n119), .IN3(n24057), .IN4(n162), .Q(n3331)
         );
  OA221X1 U3269 ( .IN1(n24001), .IN2(n205), .IN3(n24009), .IN4(n248), .IN5(
        n3332), .Q(n3329) );
  OA22X1 U3270 ( .IN1(n24017), .IN2(n291), .IN3(n24025), .IN4(n334), .Q(n3332)
         );
  OA221X1 U3271 ( .IN1(n23969), .IN2(n377), .IN3(n23977), .IN4(n420), .IN5(
        n3333), .Q(n3328) );
  OA22X1 U3272 ( .IN1(n23985), .IN2(n463), .IN3(n23993), .IN4(n506), .Q(n3333)
         );
  OA221X1 U3273 ( .IN1(n23937), .IN2(n549), .IN3(n23945), .IN4(n592), .IN5(
        n3334), .Q(n3327) );
  OA22X1 U3274 ( .IN1(n23953), .IN2(n635), .IN3(n23961), .IN4(n678), .Q(n3334)
         );
  NAND4X0 U3275 ( .IN1(n3335), .IN2(n3336), .IN3(n3337), .IN4(n3338), .QN(
        n3325) );
  OA221X1 U3276 ( .IN1(n23905), .IN2(n33), .IN3(n23913), .IN4(n76), .IN5(n3339), .Q(n3338) );
  OA22X1 U3277 ( .IN1(n23921), .IN2(n119), .IN3(n23929), .IN4(n162), .Q(n3339)
         );
  OA221X1 U3278 ( .IN1(n23873), .IN2(n205), .IN3(n23881), .IN4(n248), .IN5(
        n3340), .Q(n3337) );
  OA22X1 U3279 ( .IN1(n23889), .IN2(n291), .IN3(n23897), .IN4(n334), .Q(n3340)
         );
  OA221X1 U3280 ( .IN1(n23841), .IN2(n377), .IN3(n23849), .IN4(n420), .IN5(
        n3341), .Q(n3336) );
  OA22X1 U3281 ( .IN1(n23857), .IN2(n463), .IN3(n23865), .IN4(n506), .Q(n3341)
         );
  OA221X1 U3282 ( .IN1(n23809), .IN2(n549), .IN3(n23817), .IN4(n592), .IN5(
        n3342), .Q(n3335) );
  OA22X1 U3283 ( .IN1(n23825), .IN2(n635), .IN3(n23833), .IN4(n678), .Q(n3342)
         );
  NAND4X0 U3284 ( .IN1(n3343), .IN2(n3344), .IN3(n3345), .IN4(n3346), .QN(
        n3323) );
  OA221X1 U3285 ( .IN1(n23777), .IN2(n33), .IN3(n23785), .IN4(n76), .IN5(n3347), .Q(n3346) );
  OA22X1 U3286 ( .IN1(n23793), .IN2(n119), .IN3(n23801), .IN4(n162), .Q(n3347)
         );
  OA221X1 U3287 ( .IN1(n23745), .IN2(n205), .IN3(n23753), .IN4(n248), .IN5(
        n3348), .Q(n3345) );
  OA22X1 U3288 ( .IN1(n23761), .IN2(n291), .IN3(n23769), .IN4(n334), .Q(n3348)
         );
  OA221X1 U3289 ( .IN1(n23713), .IN2(n377), .IN3(n23721), .IN4(n420), .IN5(
        n3349), .Q(n3344) );
  OA22X1 U3290 ( .IN1(n23729), .IN2(n463), .IN3(n23737), .IN4(n506), .Q(n3349)
         );
  OA221X1 U3291 ( .IN1(n23681), .IN2(n549), .IN3(n23689), .IN4(n592), .IN5(
        n3350), .Q(n3343) );
  OA22X1 U3292 ( .IN1(n23697), .IN2(n635), .IN3(n23705), .IN4(n678), .Q(n3350)
         );
  NAND4X0 U3293 ( .IN1(n3351), .IN2(n3352), .IN3(n3353), .IN4(n3354), .QN(
        n3322) );
  OA221X1 U3294 ( .IN1(n23649), .IN2(n33), .IN3(n23657), .IN4(n76), .IN5(n3355), .Q(n3354) );
  OA22X1 U3295 ( .IN1(n23665), .IN2(n119), .IN3(n23673), .IN4(n162), .Q(n3355)
         );
  OA221X1 U3296 ( .IN1(n23617), .IN2(n205), .IN3(n23625), .IN4(n248), .IN5(
        n3356), .Q(n3353) );
  OA22X1 U3297 ( .IN1(n23633), .IN2(n291), .IN3(n23641), .IN4(n334), .Q(n3356)
         );
  OA221X1 U3298 ( .IN1(n23585), .IN2(n377), .IN3(n23593), .IN4(n420), .IN5(
        n3357), .Q(n3352) );
  OA22X1 U3299 ( .IN1(n23601), .IN2(n463), .IN3(n23609), .IN4(n506), .Q(n3357)
         );
  OA221X1 U3300 ( .IN1(n23553), .IN2(n549), .IN3(n23561), .IN4(n592), .IN5(
        n3358), .Q(n3351) );
  OA22X1 U3301 ( .IN1(n23569), .IN2(n635), .IN3(n23577), .IN4(n678), .Q(n3358)
         );
  AO221X1 U3302 ( .IN1(n2287), .IN2(n3359), .IN3(n2289), .IN4(n3360), .IN5(
        n3361), .Q(n3282) );
  AO22X1 U3303 ( .IN1(n2292), .IN2(n3362), .IN3(n2294), .IN4(n3363), .Q(n3361)
         );
  NAND4X0 U3304 ( .IN1(n3364), .IN2(n3365), .IN3(n3366), .IN4(n3367), .QN(
        n3363) );
  OA221X1 U3305 ( .IN1(n25569), .IN2(n33), .IN3(n25577), .IN4(n76), .IN5(n3368), .Q(n3367) );
  OA22X1 U3306 ( .IN1(n25585), .IN2(n119), .IN3(n25593), .IN4(n162), .Q(n3368)
         );
  OA221X1 U3307 ( .IN1(n25537), .IN2(n205), .IN3(n25545), .IN4(n248), .IN5(
        n3369), .Q(n3366) );
  OA22X1 U3308 ( .IN1(n25553), .IN2(n291), .IN3(n25561), .IN4(n334), .Q(n3369)
         );
  OA221X1 U3309 ( .IN1(n25505), .IN2(n377), .IN3(n25513), .IN4(n420), .IN5(
        n3370), .Q(n3365) );
  OA22X1 U3310 ( .IN1(n25521), .IN2(n463), .IN3(n25529), .IN4(n506), .Q(n3370)
         );
  OA221X1 U3311 ( .IN1(n25473), .IN2(n549), .IN3(n25481), .IN4(n592), .IN5(
        n3371), .Q(n3364) );
  OA22X1 U3312 ( .IN1(n25489), .IN2(n635), .IN3(n25497), .IN4(n678), .Q(n3371)
         );
  NAND4X0 U3313 ( .IN1(n3372), .IN2(n3373), .IN3(n3374), .IN4(n3375), .QN(
        n3362) );
  OA221X1 U3314 ( .IN1(n25441), .IN2(n33), .IN3(n25449), .IN4(n76), .IN5(n3376), .Q(n3375) );
  OA22X1 U3315 ( .IN1(n25457), .IN2(n119), .IN3(n25465), .IN4(n162), .Q(n3376)
         );
  OA221X1 U3316 ( .IN1(n25409), .IN2(n205), .IN3(n25417), .IN4(n248), .IN5(
        n3377), .Q(n3374) );
  OA22X1 U3317 ( .IN1(n25425), .IN2(n291), .IN3(n25433), .IN4(n334), .Q(n3377)
         );
  OA221X1 U3318 ( .IN1(n25377), .IN2(n377), .IN3(n25385), .IN4(n420), .IN5(
        n3378), .Q(n3373) );
  OA22X1 U3319 ( .IN1(n25393), .IN2(n463), .IN3(n25401), .IN4(n506), .Q(n3378)
         );
  OA221X1 U3320 ( .IN1(n25345), .IN2(n549), .IN3(n25353), .IN4(n592), .IN5(
        n3379), .Q(n3372) );
  OA22X1 U3321 ( .IN1(n25361), .IN2(n635), .IN3(n25369), .IN4(n678), .Q(n3379)
         );
  NAND4X0 U3322 ( .IN1(n3380), .IN2(n3381), .IN3(n3382), .IN4(n3383), .QN(
        n3360) );
  OA221X1 U3323 ( .IN1(n25313), .IN2(n33), .IN3(n25321), .IN4(n76), .IN5(n3384), .Q(n3383) );
  OA22X1 U3324 ( .IN1(n25329), .IN2(n119), .IN3(n25337), .IN4(n162), .Q(n3384)
         );
  OA221X1 U3325 ( .IN1(n25281), .IN2(n205), .IN3(n25289), .IN4(n248), .IN5(
        n3385), .Q(n3382) );
  OA22X1 U3326 ( .IN1(n25297), .IN2(n291), .IN3(n25305), .IN4(n334), .Q(n3385)
         );
  OA221X1 U3327 ( .IN1(n25249), .IN2(n377), .IN3(n25257), .IN4(n420), .IN5(
        n3386), .Q(n3381) );
  OA22X1 U3328 ( .IN1(n25265), .IN2(n463), .IN3(n25273), .IN4(n506), .Q(n3386)
         );
  OA221X1 U3329 ( .IN1(n25217), .IN2(n549), .IN3(n25225), .IN4(n592), .IN5(
        n3387), .Q(n3380) );
  OA22X1 U3330 ( .IN1(n25233), .IN2(n635), .IN3(n25241), .IN4(n678), .Q(n3387)
         );
  NAND4X0 U3331 ( .IN1(n3388), .IN2(n3389), .IN3(n3390), .IN4(n3391), .QN(
        n3359) );
  OA221X1 U3332 ( .IN1(n25185), .IN2(n33), .IN3(n25193), .IN4(n76), .IN5(n3392), .Q(n3391) );
  OA22X1 U3333 ( .IN1(n25201), .IN2(n119), .IN3(n25209), .IN4(n162), .Q(n3392)
         );
  OA221X1 U3334 ( .IN1(n25153), .IN2(n205), .IN3(n25161), .IN4(n248), .IN5(
        n3393), .Q(n3390) );
  OA22X1 U3335 ( .IN1(n25169), .IN2(n291), .IN3(n25177), .IN4(n334), .Q(n3393)
         );
  OA221X1 U3336 ( .IN1(n25121), .IN2(n377), .IN3(n25129), .IN4(n420), .IN5(
        n3394), .Q(n3389) );
  OA22X1 U3337 ( .IN1(n25137), .IN2(n463), .IN3(n25145), .IN4(n506), .Q(n3394)
         );
  OA221X1 U3338 ( .IN1(n25089), .IN2(n549), .IN3(n25097), .IN4(n592), .IN5(
        n3395), .Q(n3388) );
  OA22X1 U3339 ( .IN1(n25105), .IN2(n635), .IN3(n25113), .IN4(n678), .Q(n3395)
         );
  AO221X1 U3340 ( .IN1(n2328), .IN2(n3396), .IN3(n2330), .IN4(n3397), .IN5(
        n3398), .Q(n3281) );
  AO22X1 U3341 ( .IN1(n2333), .IN2(n3399), .IN3(n2335), .IN4(n3400), .Q(n3398)
         );
  NAND4X0 U3342 ( .IN1(n3401), .IN2(n3402), .IN3(n3403), .IN4(n3404), .QN(
        n3400) );
  OA221X1 U3343 ( .IN1(n25057), .IN2(n33), .IN3(n25065), .IN4(n76), .IN5(n3405), .Q(n3404) );
  OA22X1 U3344 ( .IN1(n25073), .IN2(n119), .IN3(n25081), .IN4(n162), .Q(n3405)
         );
  OA221X1 U3345 ( .IN1(n25025), .IN2(n205), .IN3(n25033), .IN4(n248), .IN5(
        n3406), .Q(n3403) );
  OA22X1 U3346 ( .IN1(n25041), .IN2(n291), .IN3(n25049), .IN4(n334), .Q(n3406)
         );
  OA221X1 U3347 ( .IN1(n24993), .IN2(n377), .IN3(n25001), .IN4(n420), .IN5(
        n3407), .Q(n3402) );
  OA22X1 U3348 ( .IN1(n25009), .IN2(n463), .IN3(n25017), .IN4(n506), .Q(n3407)
         );
  OA221X1 U3349 ( .IN1(n24961), .IN2(n549), .IN3(n24969), .IN4(n592), .IN5(
        n3408), .Q(n3401) );
  OA22X1 U3350 ( .IN1(n24977), .IN2(n635), .IN3(n24985), .IN4(n678), .Q(n3408)
         );
  NAND4X0 U3351 ( .IN1(n3409), .IN2(n3410), .IN3(n3411), .IN4(n3412), .QN(
        n3399) );
  OA221X1 U3352 ( .IN1(n24929), .IN2(n33), .IN3(n24937), .IN4(n76), .IN5(n3413), .Q(n3412) );
  OA22X1 U3353 ( .IN1(n24945), .IN2(n119), .IN3(n24953), .IN4(n162), .Q(n3413)
         );
  OA221X1 U3354 ( .IN1(n24897), .IN2(n205), .IN3(n24905), .IN4(n248), .IN5(
        n3414), .Q(n3411) );
  OA22X1 U3355 ( .IN1(n24913), .IN2(n291), .IN3(n24921), .IN4(n334), .Q(n3414)
         );
  OA221X1 U3356 ( .IN1(n24865), .IN2(n377), .IN3(n24873), .IN4(n420), .IN5(
        n3415), .Q(n3410) );
  OA22X1 U3357 ( .IN1(n24881), .IN2(n463), .IN3(n24889), .IN4(n506), .Q(n3415)
         );
  OA221X1 U3358 ( .IN1(n24833), .IN2(n549), .IN3(n24841), .IN4(n592), .IN5(
        n3416), .Q(n3409) );
  OA22X1 U3359 ( .IN1(n24849), .IN2(n635), .IN3(n24857), .IN4(n678), .Q(n3416)
         );
  NAND4X0 U3360 ( .IN1(n3417), .IN2(n3418), .IN3(n3419), .IN4(n3420), .QN(
        n3397) );
  OA221X1 U3361 ( .IN1(n24801), .IN2(n33), .IN3(n24809), .IN4(n76), .IN5(n3421), .Q(n3420) );
  OA22X1 U3362 ( .IN1(n24817), .IN2(n119), .IN3(n24825), .IN4(n162), .Q(n3421)
         );
  OA221X1 U3363 ( .IN1(n24769), .IN2(n205), .IN3(n24777), .IN4(n248), .IN5(
        n3422), .Q(n3419) );
  OA22X1 U3364 ( .IN1(n24785), .IN2(n291), .IN3(n24793), .IN4(n334), .Q(n3422)
         );
  OA221X1 U3365 ( .IN1(n24737), .IN2(n377), .IN3(n24745), .IN4(n420), .IN5(
        n3423), .Q(n3418) );
  OA22X1 U3366 ( .IN1(n24753), .IN2(n463), .IN3(n24761), .IN4(n506), .Q(n3423)
         );
  OA221X1 U3367 ( .IN1(n24705), .IN2(n549), .IN3(n24713), .IN4(n592), .IN5(
        n3424), .Q(n3417) );
  OA22X1 U3368 ( .IN1(n24721), .IN2(n635), .IN3(n24729), .IN4(n678), .Q(n3424)
         );
  NAND4X0 U3369 ( .IN1(n3425), .IN2(n3426), .IN3(n3427), .IN4(n3428), .QN(
        n3396) );
  OA221X1 U3370 ( .IN1(n24673), .IN2(n33), .IN3(n24681), .IN4(n76), .IN5(n3429), .Q(n3428) );
  OA22X1 U3371 ( .IN1(n24689), .IN2(n119), .IN3(n24697), .IN4(n162), .Q(n3429)
         );
  OA221X1 U3372 ( .IN1(n24641), .IN2(n205), .IN3(n24649), .IN4(n248), .IN5(
        n3430), .Q(n3427) );
  OA22X1 U3373 ( .IN1(n24657), .IN2(n291), .IN3(n24665), .IN4(n334), .Q(n3430)
         );
  OA221X1 U3374 ( .IN1(n24609), .IN2(n377), .IN3(n24617), .IN4(n420), .IN5(
        n3431), .Q(n3426) );
  OA22X1 U3375 ( .IN1(n24625), .IN2(n463), .IN3(n24633), .IN4(n506), .Q(n3431)
         );
  OA221X1 U3376 ( .IN1(n24577), .IN2(n549), .IN3(n24585), .IN4(n592), .IN5(
        n3432), .Q(n3425) );
  OA22X1 U3377 ( .IN1(n24593), .IN2(n635), .IN3(n24601), .IN4(n678), .Q(n3432)
         );
  OR4X1 U3378 ( .IN1(n3433), .IN2(n3434), .IN3(n3435), .IN4(n3436), .Q(n2195)
         );
  AO221X1 U3379 ( .IN1(n2157), .IN2(n3437), .IN3(n2159), .IN4(n3438), .IN5(
        n3439), .Q(n3436) );
  AO22X1 U3380 ( .IN1(n2162), .IN2(n3440), .IN3(n2164), .IN4(n3441), .Q(n3439)
         );
  NAND4X0 U3381 ( .IN1(n3442), .IN2(n3443), .IN3(n3444), .IN4(n3445), .QN(
        n3441) );
  OA221X1 U3382 ( .IN1(n26600), .IN2(n32), .IN3(n26608), .IN4(n75), .IN5(n3446), .Q(n3445) );
  OA22X1 U3383 ( .IN1(n26616), .IN2(n118), .IN3(n26624), .IN4(n161), .Q(n3446)
         );
  OA221X1 U3384 ( .IN1(n26568), .IN2(n204), .IN3(n26576), .IN4(n247), .IN5(
        n3447), .Q(n3444) );
  OA22X1 U3385 ( .IN1(n26584), .IN2(n290), .IN3(n26592), .IN4(n333), .Q(n3447)
         );
  OA221X1 U3386 ( .IN1(n26536), .IN2(n376), .IN3(n26544), .IN4(n419), .IN5(
        n3448), .Q(n3443) );
  OA22X1 U3387 ( .IN1(n26552), .IN2(n462), .IN3(n26560), .IN4(n505), .Q(n3448)
         );
  OA221X1 U3388 ( .IN1(n26504), .IN2(n548), .IN3(n26512), .IN4(n591), .IN5(
        n3449), .Q(n3442) );
  OA22X1 U3389 ( .IN1(n26520), .IN2(n634), .IN3(n26528), .IN4(n677), .Q(n3449)
         );
  NAND4X0 U3390 ( .IN1(n3450), .IN2(n3451), .IN3(n3452), .IN4(n3453), .QN(
        n3440) );
  OA221X1 U3391 ( .IN1(n26472), .IN2(n32), .IN3(n26480), .IN4(n75), .IN5(n3454), .Q(n3453) );
  OA22X1 U3392 ( .IN1(n26488), .IN2(n118), .IN3(n26496), .IN4(n161), .Q(n3454)
         );
  OA221X1 U3393 ( .IN1(n26440), .IN2(n204), .IN3(n26448), .IN4(n247), .IN5(
        n3455), .Q(n3452) );
  OA22X1 U3394 ( .IN1(n26456), .IN2(n290), .IN3(n26464), .IN4(n333), .Q(n3455)
         );
  OA221X1 U3395 ( .IN1(n26408), .IN2(n376), .IN3(n26416), .IN4(n419), .IN5(
        n3456), .Q(n3451) );
  OA22X1 U3396 ( .IN1(n26424), .IN2(n462), .IN3(n26432), .IN4(n505), .Q(n3456)
         );
  OA221X1 U3397 ( .IN1(n26376), .IN2(n548), .IN3(n26384), .IN4(n591), .IN5(
        n3457), .Q(n3450) );
  OA22X1 U3398 ( .IN1(n26392), .IN2(n634), .IN3(n26400), .IN4(n677), .Q(n3457)
         );
  NAND4X0 U3399 ( .IN1(n3458), .IN2(n3459), .IN3(n3460), .IN4(n3461), .QN(
        n3438) );
  OA221X1 U3400 ( .IN1(n26344), .IN2(n32), .IN3(n26352), .IN4(n75), .IN5(n3462), .Q(n3461) );
  OA22X1 U3401 ( .IN1(n26360), .IN2(n118), .IN3(n26368), .IN4(n161), .Q(n3462)
         );
  OA221X1 U3402 ( .IN1(n26312), .IN2(n204), .IN3(n26320), .IN4(n247), .IN5(
        n3463), .Q(n3460) );
  OA22X1 U3403 ( .IN1(n26328), .IN2(n290), .IN3(n26336), .IN4(n333), .Q(n3463)
         );
  OA221X1 U3404 ( .IN1(n26280), .IN2(n376), .IN3(n26288), .IN4(n419), .IN5(
        n3464), .Q(n3459) );
  OA22X1 U3405 ( .IN1(n26296), .IN2(n462), .IN3(n26304), .IN4(n505), .Q(n3464)
         );
  OA221X1 U3406 ( .IN1(n26248), .IN2(n548), .IN3(n26256), .IN4(n591), .IN5(
        n3465), .Q(n3458) );
  OA22X1 U3407 ( .IN1(n26264), .IN2(n634), .IN3(n26272), .IN4(n677), .Q(n3465)
         );
  NAND4X0 U3408 ( .IN1(n3466), .IN2(n3467), .IN3(n3468), .IN4(n3469), .QN(
        n3437) );
  OA221X1 U3409 ( .IN1(n26216), .IN2(n32), .IN3(n26224), .IN4(n75), .IN5(n3470), .Q(n3469) );
  OA22X1 U3410 ( .IN1(n26232), .IN2(n118), .IN3(n26240), .IN4(n161), .Q(n3470)
         );
  OA221X1 U3411 ( .IN1(n26184), .IN2(n204), .IN3(n26192), .IN4(n247), .IN5(
        n3471), .Q(n3468) );
  OA22X1 U3412 ( .IN1(n26200), .IN2(n290), .IN3(n26208), .IN4(n333), .Q(n3471)
         );
  OA221X1 U3413 ( .IN1(n26152), .IN2(n376), .IN3(n26160), .IN4(n419), .IN5(
        n3472), .Q(n3467) );
  OA22X1 U3414 ( .IN1(n26168), .IN2(n462), .IN3(n26176), .IN4(n505), .Q(n3472)
         );
  OA221X1 U3415 ( .IN1(n26120), .IN2(n548), .IN3(n26128), .IN4(n591), .IN5(
        n3473), .Q(n3466) );
  OA22X1 U3416 ( .IN1(n26136), .IN2(n634), .IN3(n26144), .IN4(n677), .Q(n3473)
         );
  AO221X1 U3417 ( .IN1(n2246), .IN2(n3474), .IN3(n2248), .IN4(n3475), .IN5(
        n3476), .Q(n3435) );
  AO22X1 U3418 ( .IN1(n2251), .IN2(n3477), .IN3(n2253), .IN4(n3478), .Q(n3476)
         );
  NAND4X0 U3419 ( .IN1(n3479), .IN2(n3480), .IN3(n3481), .IN4(n3482), .QN(
        n3478) );
  OA221X1 U3420 ( .IN1(n26088), .IN2(n32), .IN3(n26096), .IN4(n75), .IN5(n3483), .Q(n3482) );
  OA22X1 U3421 ( .IN1(n26104), .IN2(n118), .IN3(n26112), .IN4(n161), .Q(n3483)
         );
  OA221X1 U3422 ( .IN1(n26056), .IN2(n204), .IN3(n26064), .IN4(n247), .IN5(
        n3484), .Q(n3481) );
  OA22X1 U3423 ( .IN1(n26072), .IN2(n290), .IN3(n26080), .IN4(n333), .Q(n3484)
         );
  OA221X1 U3424 ( .IN1(n26024), .IN2(n376), .IN3(n26032), .IN4(n419), .IN5(
        n3485), .Q(n3480) );
  OA22X1 U3425 ( .IN1(n26040), .IN2(n462), .IN3(n26048), .IN4(n505), .Q(n3485)
         );
  OA221X1 U3426 ( .IN1(n25992), .IN2(n548), .IN3(n26000), .IN4(n591), .IN5(
        n3486), .Q(n3479) );
  OA22X1 U3427 ( .IN1(n26008), .IN2(n634), .IN3(n26016), .IN4(n677), .Q(n3486)
         );
  NAND4X0 U3428 ( .IN1(n3487), .IN2(n3488), .IN3(n3489), .IN4(n3490), .QN(
        n3477) );
  OA221X1 U3429 ( .IN1(n25960), .IN2(n32), .IN3(n25968), .IN4(n75), .IN5(n3491), .Q(n3490) );
  OA22X1 U3430 ( .IN1(n25976), .IN2(n118), .IN3(n25984), .IN4(n161), .Q(n3491)
         );
  OA221X1 U3431 ( .IN1(n25928), .IN2(n204), .IN3(n25936), .IN4(n247), .IN5(
        n3492), .Q(n3489) );
  OA22X1 U3432 ( .IN1(n25944), .IN2(n290), .IN3(n25952), .IN4(n333), .Q(n3492)
         );
  OA221X1 U3433 ( .IN1(n25896), .IN2(n376), .IN3(n25904), .IN4(n419), .IN5(
        n3493), .Q(n3488) );
  OA22X1 U3434 ( .IN1(n25912), .IN2(n462), .IN3(n25920), .IN4(n505), .Q(n3493)
         );
  OA221X1 U3435 ( .IN1(n25864), .IN2(n548), .IN3(n25872), .IN4(n591), .IN5(
        n3494), .Q(n3487) );
  OA22X1 U3436 ( .IN1(n25880), .IN2(n634), .IN3(n25888), .IN4(n677), .Q(n3494)
         );
  NAND4X0 U3437 ( .IN1(n3495), .IN2(n3496), .IN3(n3497), .IN4(n3498), .QN(
        n3475) );
  OA221X1 U3438 ( .IN1(n25832), .IN2(n32), .IN3(n25840), .IN4(n75), .IN5(n3499), .Q(n3498) );
  OA22X1 U3439 ( .IN1(n25848), .IN2(n118), .IN3(n25856), .IN4(n161), .Q(n3499)
         );
  OA221X1 U3440 ( .IN1(n25800), .IN2(n204), .IN3(n25808), .IN4(n247), .IN5(
        n3500), .Q(n3497) );
  OA22X1 U3441 ( .IN1(n25816), .IN2(n290), .IN3(n25824), .IN4(n333), .Q(n3500)
         );
  OA221X1 U3442 ( .IN1(n25768), .IN2(n376), .IN3(n25776), .IN4(n419), .IN5(
        n3501), .Q(n3496) );
  OA22X1 U3443 ( .IN1(n25784), .IN2(n462), .IN3(n25792), .IN4(n505), .Q(n3501)
         );
  OA221X1 U3444 ( .IN1(n25736), .IN2(n548), .IN3(n25744), .IN4(n591), .IN5(
        n3502), .Q(n3495) );
  OA22X1 U3445 ( .IN1(n25752), .IN2(n634), .IN3(n25760), .IN4(n677), .Q(n3502)
         );
  NAND4X0 U3446 ( .IN1(n3503), .IN2(n3504), .IN3(n3505), .IN4(n3506), .QN(
        n3474) );
  OA221X1 U3447 ( .IN1(n25704), .IN2(n32), .IN3(n25712), .IN4(n75), .IN5(n3507), .Q(n3506) );
  OA22X1 U3448 ( .IN1(n25720), .IN2(n118), .IN3(n25728), .IN4(n161), .Q(n3507)
         );
  OA221X1 U3449 ( .IN1(n25672), .IN2(n204), .IN3(n25680), .IN4(n247), .IN5(
        n3508), .Q(n3505) );
  OA22X1 U3450 ( .IN1(n25688), .IN2(n290), .IN3(n25696), .IN4(n333), .Q(n3508)
         );
  OA221X1 U3451 ( .IN1(n25640), .IN2(n376), .IN3(n25648), .IN4(n419), .IN5(
        n3509), .Q(n3504) );
  OA22X1 U3452 ( .IN1(n25656), .IN2(n462), .IN3(n25664), .IN4(n505), .Q(n3509)
         );
  OA221X1 U3453 ( .IN1(n25608), .IN2(n548), .IN3(n25616), .IN4(n591), .IN5(
        n3510), .Q(n3503) );
  OA22X1 U3454 ( .IN1(n25624), .IN2(n634), .IN3(n25632), .IN4(n677), .Q(n3510)
         );
  AO221X1 U3455 ( .IN1(n2287), .IN2(n3511), .IN3(n2289), .IN4(n3512), .IN5(
        n3513), .Q(n3434) );
  AO22X1 U3456 ( .IN1(n2292), .IN2(n3514), .IN3(n2294), .IN4(n3515), .Q(n3513)
         );
  NAND4X0 U3457 ( .IN1(n3516), .IN2(n3517), .IN3(n3518), .IN4(n3519), .QN(
        n3515) );
  OA221X1 U3458 ( .IN1(n27624), .IN2(n32), .IN3(n27632), .IN4(n75), .IN5(n3520), .Q(n3519) );
  OA22X1 U3459 ( .IN1(n27640), .IN2(n118), .IN3(n27648), .IN4(n161), .Q(n3520)
         );
  OA221X1 U3460 ( .IN1(n27592), .IN2(n204), .IN3(n27600), .IN4(n247), .IN5(
        n3521), .Q(n3518) );
  OA22X1 U3461 ( .IN1(n27608), .IN2(n290), .IN3(n27616), .IN4(n333), .Q(n3521)
         );
  OA221X1 U3462 ( .IN1(n27560), .IN2(n376), .IN3(n27568), .IN4(n419), .IN5(
        n3522), .Q(n3517) );
  OA22X1 U3463 ( .IN1(n27576), .IN2(n462), .IN3(n27584), .IN4(n505), .Q(n3522)
         );
  OA221X1 U3464 ( .IN1(n27528), .IN2(n548), .IN3(n27536), .IN4(n591), .IN5(
        n3523), .Q(n3516) );
  OA22X1 U3465 ( .IN1(n27544), .IN2(n634), .IN3(n27552), .IN4(n677), .Q(n3523)
         );
  NAND4X0 U3466 ( .IN1(n3524), .IN2(n3525), .IN3(n3526), .IN4(n3527), .QN(
        n3514) );
  OA221X1 U3467 ( .IN1(n27496), .IN2(n32), .IN3(n27504), .IN4(n75), .IN5(n3528), .Q(n3527) );
  OA22X1 U3468 ( .IN1(n27512), .IN2(n118), .IN3(n27520), .IN4(n161), .Q(n3528)
         );
  OA221X1 U3469 ( .IN1(n27464), .IN2(n204), .IN3(n27472), .IN4(n247), .IN5(
        n3529), .Q(n3526) );
  OA22X1 U3470 ( .IN1(n27480), .IN2(n290), .IN3(n27488), .IN4(n333), .Q(n3529)
         );
  OA221X1 U3471 ( .IN1(n27432), .IN2(n376), .IN3(n27440), .IN4(n419), .IN5(
        n3530), .Q(n3525) );
  OA22X1 U3472 ( .IN1(n27448), .IN2(n462), .IN3(n27456), .IN4(n505), .Q(n3530)
         );
  OA221X1 U3473 ( .IN1(n27400), .IN2(n548), .IN3(n27408), .IN4(n591), .IN5(
        n3531), .Q(n3524) );
  OA22X1 U3474 ( .IN1(n27416), .IN2(n634), .IN3(n27424), .IN4(n677), .Q(n3531)
         );
  NAND4X0 U3475 ( .IN1(n3532), .IN2(n3533), .IN3(n3534), .IN4(n3535), .QN(
        n3512) );
  OA221X1 U3476 ( .IN1(n27368), .IN2(n32), .IN3(n27376), .IN4(n75), .IN5(n3536), .Q(n3535) );
  OA22X1 U3477 ( .IN1(n27384), .IN2(n118), .IN3(n27392), .IN4(n161), .Q(n3536)
         );
  OA221X1 U3478 ( .IN1(n27336), .IN2(n204), .IN3(n27344), .IN4(n247), .IN5(
        n3537), .Q(n3534) );
  OA22X1 U3479 ( .IN1(n27352), .IN2(n290), .IN3(n27360), .IN4(n333), .Q(n3537)
         );
  OA221X1 U3480 ( .IN1(n27304), .IN2(n376), .IN3(n27312), .IN4(n419), .IN5(
        n3538), .Q(n3533) );
  OA22X1 U3481 ( .IN1(n27320), .IN2(n462), .IN3(n27328), .IN4(n505), .Q(n3538)
         );
  OA221X1 U3482 ( .IN1(n27272), .IN2(n548), .IN3(n27280), .IN4(n591), .IN5(
        n3539), .Q(n3532) );
  OA22X1 U3483 ( .IN1(n27288), .IN2(n634), .IN3(n27296), .IN4(n677), .Q(n3539)
         );
  NAND4X0 U3484 ( .IN1(n3540), .IN2(n3541), .IN3(n3542), .IN4(n3543), .QN(
        n3511) );
  OA221X1 U3485 ( .IN1(n27240), .IN2(n32), .IN3(n27248), .IN4(n75), .IN5(n3544), .Q(n3543) );
  OA22X1 U3486 ( .IN1(n27256), .IN2(n118), .IN3(n27264), .IN4(n161), .Q(n3544)
         );
  OA221X1 U3487 ( .IN1(n27208), .IN2(n204), .IN3(n27216), .IN4(n247), .IN5(
        n3545), .Q(n3542) );
  OA22X1 U3488 ( .IN1(n27224), .IN2(n290), .IN3(n27232), .IN4(n333), .Q(n3545)
         );
  OA221X1 U3489 ( .IN1(n27176), .IN2(n376), .IN3(n27184), .IN4(n419), .IN5(
        n3546), .Q(n3541) );
  OA22X1 U3490 ( .IN1(n27192), .IN2(n462), .IN3(n27200), .IN4(n505), .Q(n3546)
         );
  OA221X1 U3491 ( .IN1(n27144), .IN2(n548), .IN3(n27152), .IN4(n591), .IN5(
        n3547), .Q(n3540) );
  OA22X1 U3492 ( .IN1(n27160), .IN2(n634), .IN3(n27168), .IN4(n677), .Q(n3547)
         );
  AO221X1 U3493 ( .IN1(n2328), .IN2(n3548), .IN3(n2330), .IN4(n3549), .IN5(
        n3550), .Q(n3433) );
  AO22X1 U3494 ( .IN1(n2333), .IN2(n3551), .IN3(n2335), .IN4(n3552), .Q(n3550)
         );
  NAND4X0 U3495 ( .IN1(n3553), .IN2(n3554), .IN3(n3555), .IN4(n3556), .QN(
        n3552) );
  OA221X1 U3496 ( .IN1(n27112), .IN2(n31), .IN3(n27120), .IN4(n74), .IN5(n3557), .Q(n3556) );
  OA22X1 U3497 ( .IN1(n27128), .IN2(n117), .IN3(n27136), .IN4(n160), .Q(n3557)
         );
  OA221X1 U3498 ( .IN1(n27080), .IN2(n203), .IN3(n27088), .IN4(n246), .IN5(
        n3558), .Q(n3555) );
  OA22X1 U3499 ( .IN1(n27096), .IN2(n289), .IN3(n27104), .IN4(n332), .Q(n3558)
         );
  OA221X1 U3500 ( .IN1(n27048), .IN2(n375), .IN3(n27056), .IN4(n418), .IN5(
        n3559), .Q(n3554) );
  OA22X1 U3501 ( .IN1(n27064), .IN2(n461), .IN3(n27072), .IN4(n504), .Q(n3559)
         );
  OA221X1 U3502 ( .IN1(n27016), .IN2(n547), .IN3(n27024), .IN4(n590), .IN5(
        n3560), .Q(n3553) );
  OA22X1 U3503 ( .IN1(n27032), .IN2(n633), .IN3(n27040), .IN4(n676), .Q(n3560)
         );
  NAND4X0 U3504 ( .IN1(n3561), .IN2(n3562), .IN3(n3563), .IN4(n3564), .QN(
        n3551) );
  OA221X1 U3505 ( .IN1(n26984), .IN2(n31), .IN3(n26992), .IN4(n74), .IN5(n3565), .Q(n3564) );
  OA22X1 U3506 ( .IN1(n27000), .IN2(n117), .IN3(n27008), .IN4(n160), .Q(n3565)
         );
  OA221X1 U3507 ( .IN1(n26952), .IN2(n203), .IN3(n26960), .IN4(n246), .IN5(
        n3566), .Q(n3563) );
  OA22X1 U3508 ( .IN1(n26968), .IN2(n289), .IN3(n26976), .IN4(n332), .Q(n3566)
         );
  OA221X1 U3509 ( .IN1(n26920), .IN2(n375), .IN3(n26928), .IN4(n418), .IN5(
        n3567), .Q(n3562) );
  OA22X1 U3510 ( .IN1(n26936), .IN2(n461), .IN3(n26944), .IN4(n504), .Q(n3567)
         );
  OA221X1 U3511 ( .IN1(n26888), .IN2(n547), .IN3(n26896), .IN4(n590), .IN5(
        n3568), .Q(n3561) );
  OA22X1 U3512 ( .IN1(n26904), .IN2(n633), .IN3(n26912), .IN4(n676), .Q(n3568)
         );
  NAND4X0 U3513 ( .IN1(n3569), .IN2(n3570), .IN3(n3571), .IN4(n3572), .QN(
        n3549) );
  OA221X1 U3514 ( .IN1(n26856), .IN2(n31), .IN3(n26864), .IN4(n74), .IN5(n3573), .Q(n3572) );
  OA22X1 U3515 ( .IN1(n26872), .IN2(n117), .IN3(n26880), .IN4(n160), .Q(n3573)
         );
  OA221X1 U3516 ( .IN1(n26824), .IN2(n203), .IN3(n26832), .IN4(n246), .IN5(
        n3574), .Q(n3571) );
  OA22X1 U3517 ( .IN1(n26840), .IN2(n289), .IN3(n26848), .IN4(n332), .Q(n3574)
         );
  OA221X1 U3518 ( .IN1(n26792), .IN2(n375), .IN3(n26800), .IN4(n418), .IN5(
        n3575), .Q(n3570) );
  OA22X1 U3519 ( .IN1(n26808), .IN2(n461), .IN3(n26816), .IN4(n504), .Q(n3575)
         );
  OA221X1 U3520 ( .IN1(n26760), .IN2(n547), .IN3(n26768), .IN4(n590), .IN5(
        n3576), .Q(n3569) );
  OA22X1 U3521 ( .IN1(n26776), .IN2(n633), .IN3(n26784), .IN4(n676), .Q(n3576)
         );
  NAND4X0 U3522 ( .IN1(n3577), .IN2(n3578), .IN3(n3579), .IN4(n3580), .QN(
        n3548) );
  OA221X1 U3523 ( .IN1(n26728), .IN2(n31), .IN3(n26736), .IN4(n74), .IN5(n3581), .Q(n3580) );
  OA22X1 U3524 ( .IN1(n26744), .IN2(n117), .IN3(n26752), .IN4(n160), .Q(n3581)
         );
  OA221X1 U3525 ( .IN1(n26696), .IN2(n203), .IN3(n26704), .IN4(n246), .IN5(
        n3582), .Q(n3579) );
  OA22X1 U3526 ( .IN1(n26712), .IN2(n289), .IN3(n26720), .IN4(n332), .Q(n3582)
         );
  OA221X1 U3527 ( .IN1(n26664), .IN2(n375), .IN3(n26672), .IN4(n418), .IN5(
        n3583), .Q(n3578) );
  OA22X1 U3528 ( .IN1(n26680), .IN2(n461), .IN3(n26688), .IN4(n504), .Q(n3583)
         );
  OA221X1 U3529 ( .IN1(n26632), .IN2(n547), .IN3(n26640), .IN4(n590), .IN5(
        n3584), .Q(n3577) );
  OA22X1 U3530 ( .IN1(n26648), .IN2(n633), .IN3(n26656), .IN4(n676), .Q(n3584)
         );
  OR4X1 U3531 ( .IN1(n3585), .IN2(n3586), .IN3(n3587), .IN4(n3588), .Q(n2193)
         );
  AO221X1 U3532 ( .IN1(n2157), .IN2(n3589), .IN3(n2159), .IN4(n3590), .IN5(
        n3591), .Q(n3588) );
  AO22X1 U3533 ( .IN1(n2162), .IN2(n3592), .IN3(n2164), .IN4(n3593), .Q(n3591)
         );
  NAND4X0 U3534 ( .IN1(n3594), .IN2(n3595), .IN3(n3596), .IN4(n3597), .QN(
        n3593) );
  OA221X1 U3535 ( .IN1(n26599), .IN2(n31), .IN3(n26607), .IN4(n74), .IN5(n3598), .Q(n3597) );
  OA22X1 U3536 ( .IN1(n26615), .IN2(n117), .IN3(n26623), .IN4(n160), .Q(n3598)
         );
  OA221X1 U3537 ( .IN1(n26567), .IN2(n203), .IN3(n26575), .IN4(n246), .IN5(
        n3599), .Q(n3596) );
  OA22X1 U3538 ( .IN1(n26583), .IN2(n289), .IN3(n26591), .IN4(n332), .Q(n3599)
         );
  OA221X1 U3539 ( .IN1(n26535), .IN2(n375), .IN3(n26543), .IN4(n418), .IN5(
        n3600), .Q(n3595) );
  OA22X1 U3540 ( .IN1(n26551), .IN2(n461), .IN3(n26559), .IN4(n504), .Q(n3600)
         );
  OA221X1 U3541 ( .IN1(n26503), .IN2(n547), .IN3(n26511), .IN4(n590), .IN5(
        n3601), .Q(n3594) );
  OA22X1 U3542 ( .IN1(n26519), .IN2(n633), .IN3(n26527), .IN4(n676), .Q(n3601)
         );
  NAND4X0 U3543 ( .IN1(n3602), .IN2(n3603), .IN3(n3604), .IN4(n3605), .QN(
        n3592) );
  OA221X1 U3544 ( .IN1(n26471), .IN2(n31), .IN3(n26479), .IN4(n74), .IN5(n3606), .Q(n3605) );
  OA22X1 U3545 ( .IN1(n26487), .IN2(n117), .IN3(n26495), .IN4(n160), .Q(n3606)
         );
  OA221X1 U3546 ( .IN1(n26439), .IN2(n203), .IN3(n26447), .IN4(n246), .IN5(
        n3607), .Q(n3604) );
  OA22X1 U3547 ( .IN1(n26455), .IN2(n289), .IN3(n26463), .IN4(n332), .Q(n3607)
         );
  OA221X1 U3548 ( .IN1(n26407), .IN2(n375), .IN3(n26415), .IN4(n418), .IN5(
        n3608), .Q(n3603) );
  OA22X1 U3549 ( .IN1(n26423), .IN2(n461), .IN3(n26431), .IN4(n504), .Q(n3608)
         );
  OA221X1 U3550 ( .IN1(n26375), .IN2(n547), .IN3(n26383), .IN4(n590), .IN5(
        n3609), .Q(n3602) );
  OA22X1 U3551 ( .IN1(n26391), .IN2(n633), .IN3(n26399), .IN4(n676), .Q(n3609)
         );
  NAND4X0 U3552 ( .IN1(n3610), .IN2(n3611), .IN3(n3612), .IN4(n3613), .QN(
        n3590) );
  OA221X1 U3553 ( .IN1(n26343), .IN2(n31), .IN3(n26351), .IN4(n74), .IN5(n3614), .Q(n3613) );
  OA22X1 U3554 ( .IN1(n26359), .IN2(n117), .IN3(n26367), .IN4(n160), .Q(n3614)
         );
  OA221X1 U3555 ( .IN1(n26311), .IN2(n203), .IN3(n26319), .IN4(n246), .IN5(
        n3615), .Q(n3612) );
  OA22X1 U3556 ( .IN1(n26327), .IN2(n289), .IN3(n26335), .IN4(n332), .Q(n3615)
         );
  OA221X1 U3557 ( .IN1(n26279), .IN2(n375), .IN3(n26287), .IN4(n418), .IN5(
        n3616), .Q(n3611) );
  OA22X1 U3558 ( .IN1(n26295), .IN2(n461), .IN3(n26303), .IN4(n504), .Q(n3616)
         );
  OA221X1 U3559 ( .IN1(n26247), .IN2(n547), .IN3(n26255), .IN4(n590), .IN5(
        n3617), .Q(n3610) );
  OA22X1 U3560 ( .IN1(n26263), .IN2(n633), .IN3(n26271), .IN4(n676), .Q(n3617)
         );
  NAND4X0 U3561 ( .IN1(n3618), .IN2(n3619), .IN3(n3620), .IN4(n3621), .QN(
        n3589) );
  OA221X1 U3562 ( .IN1(n26215), .IN2(n31), .IN3(n26223), .IN4(n74), .IN5(n3622), .Q(n3621) );
  OA22X1 U3563 ( .IN1(n26231), .IN2(n117), .IN3(n26239), .IN4(n160), .Q(n3622)
         );
  OA221X1 U3564 ( .IN1(n26183), .IN2(n203), .IN3(n26191), .IN4(n246), .IN5(
        n3623), .Q(n3620) );
  OA22X1 U3565 ( .IN1(n26199), .IN2(n289), .IN3(n26207), .IN4(n332), .Q(n3623)
         );
  OA221X1 U3566 ( .IN1(n26151), .IN2(n375), .IN3(n26159), .IN4(n418), .IN5(
        n3624), .Q(n3619) );
  OA22X1 U3567 ( .IN1(n26167), .IN2(n461), .IN3(n26175), .IN4(n504), .Q(n3624)
         );
  OA221X1 U3568 ( .IN1(n26119), .IN2(n547), .IN3(n26127), .IN4(n590), .IN5(
        n3625), .Q(n3618) );
  OA22X1 U3569 ( .IN1(n26135), .IN2(n633), .IN3(n26143), .IN4(n676), .Q(n3625)
         );
  AO221X1 U3570 ( .IN1(n2246), .IN2(n3626), .IN3(n2248), .IN4(n3627), .IN5(
        n3628), .Q(n3587) );
  AO22X1 U3571 ( .IN1(n2251), .IN2(n3629), .IN3(n2253), .IN4(n3630), .Q(n3628)
         );
  NAND4X0 U3572 ( .IN1(n3631), .IN2(n3632), .IN3(n3633), .IN4(n3634), .QN(
        n3630) );
  OA221X1 U3573 ( .IN1(n26087), .IN2(n31), .IN3(n26095), .IN4(n74), .IN5(n3635), .Q(n3634) );
  OA22X1 U3574 ( .IN1(n26103), .IN2(n117), .IN3(n26111), .IN4(n160), .Q(n3635)
         );
  OA221X1 U3575 ( .IN1(n26055), .IN2(n203), .IN3(n26063), .IN4(n246), .IN5(
        n3636), .Q(n3633) );
  OA22X1 U3576 ( .IN1(n26071), .IN2(n289), .IN3(n26079), .IN4(n332), .Q(n3636)
         );
  OA221X1 U3577 ( .IN1(n26023), .IN2(n375), .IN3(n26031), .IN4(n418), .IN5(
        n3637), .Q(n3632) );
  OA22X1 U3578 ( .IN1(n26039), .IN2(n461), .IN3(n26047), .IN4(n504), .Q(n3637)
         );
  OA221X1 U3579 ( .IN1(n25991), .IN2(n547), .IN3(n25999), .IN4(n590), .IN5(
        n3638), .Q(n3631) );
  OA22X1 U3580 ( .IN1(n26007), .IN2(n633), .IN3(n26015), .IN4(n676), .Q(n3638)
         );
  NAND4X0 U3581 ( .IN1(n3639), .IN2(n3640), .IN3(n3641), .IN4(n3642), .QN(
        n3629) );
  OA221X1 U3582 ( .IN1(n25959), .IN2(n31), .IN3(n25967), .IN4(n74), .IN5(n3643), .Q(n3642) );
  OA22X1 U3583 ( .IN1(n25975), .IN2(n117), .IN3(n25983), .IN4(n160), .Q(n3643)
         );
  OA221X1 U3584 ( .IN1(n25927), .IN2(n203), .IN3(n25935), .IN4(n246), .IN5(
        n3644), .Q(n3641) );
  OA22X1 U3585 ( .IN1(n25943), .IN2(n289), .IN3(n25951), .IN4(n332), .Q(n3644)
         );
  OA221X1 U3586 ( .IN1(n25895), .IN2(n375), .IN3(n25903), .IN4(n418), .IN5(
        n3645), .Q(n3640) );
  OA22X1 U3587 ( .IN1(n25911), .IN2(n461), .IN3(n25919), .IN4(n504), .Q(n3645)
         );
  OA221X1 U3588 ( .IN1(n25863), .IN2(n547), .IN3(n25871), .IN4(n590), .IN5(
        n3646), .Q(n3639) );
  OA22X1 U3589 ( .IN1(n25879), .IN2(n633), .IN3(n25887), .IN4(n676), .Q(n3646)
         );
  NAND4X0 U3590 ( .IN1(n3647), .IN2(n3648), .IN3(n3649), .IN4(n3650), .QN(
        n3627) );
  OA221X1 U3591 ( .IN1(n25831), .IN2(n31), .IN3(n25839), .IN4(n74), .IN5(n3651), .Q(n3650) );
  OA22X1 U3592 ( .IN1(n25847), .IN2(n117), .IN3(n25855), .IN4(n160), .Q(n3651)
         );
  OA221X1 U3593 ( .IN1(n25799), .IN2(n203), .IN3(n25807), .IN4(n246), .IN5(
        n3652), .Q(n3649) );
  OA22X1 U3594 ( .IN1(n25815), .IN2(n289), .IN3(n25823), .IN4(n332), .Q(n3652)
         );
  OA221X1 U3595 ( .IN1(n25767), .IN2(n375), .IN3(n25775), .IN4(n418), .IN5(
        n3653), .Q(n3648) );
  OA22X1 U3596 ( .IN1(n25783), .IN2(n461), .IN3(n25791), .IN4(n504), .Q(n3653)
         );
  OA221X1 U3597 ( .IN1(n25735), .IN2(n547), .IN3(n25743), .IN4(n590), .IN5(
        n3654), .Q(n3647) );
  OA22X1 U3598 ( .IN1(n25751), .IN2(n633), .IN3(n25759), .IN4(n676), .Q(n3654)
         );
  NAND4X0 U3599 ( .IN1(n3655), .IN2(n3656), .IN3(n3657), .IN4(n3658), .QN(
        n3626) );
  OA221X1 U3600 ( .IN1(n25703), .IN2(n31), .IN3(n25711), .IN4(n74), .IN5(n3659), .Q(n3658) );
  OA22X1 U3601 ( .IN1(n25719), .IN2(n117), .IN3(n25727), .IN4(n160), .Q(n3659)
         );
  OA221X1 U3602 ( .IN1(n25671), .IN2(n203), .IN3(n25679), .IN4(n246), .IN5(
        n3660), .Q(n3657) );
  OA22X1 U3603 ( .IN1(n25687), .IN2(n289), .IN3(n25695), .IN4(n332), .Q(n3660)
         );
  OA221X1 U3604 ( .IN1(n25639), .IN2(n375), .IN3(n25647), .IN4(n418), .IN5(
        n3661), .Q(n3656) );
  OA22X1 U3605 ( .IN1(n25655), .IN2(n461), .IN3(n25663), .IN4(n504), .Q(n3661)
         );
  OA221X1 U3606 ( .IN1(n25607), .IN2(n547), .IN3(n25615), .IN4(n590), .IN5(
        n3662), .Q(n3655) );
  OA22X1 U3607 ( .IN1(n25623), .IN2(n633), .IN3(n25631), .IN4(n676), .Q(n3662)
         );
  AO221X1 U3608 ( .IN1(n2287), .IN2(n3663), .IN3(n2289), .IN4(n3664), .IN5(
        n3665), .Q(n3586) );
  AO22X1 U3609 ( .IN1(n2292), .IN2(n3666), .IN3(n2294), .IN4(n3667), .Q(n3665)
         );
  NAND4X0 U3610 ( .IN1(n3668), .IN2(n3669), .IN3(n3670), .IN4(n3671), .QN(
        n3667) );
  OA221X1 U3611 ( .IN1(n27623), .IN2(n30), .IN3(n27631), .IN4(n73), .IN5(n3672), .Q(n3671) );
  OA22X1 U3612 ( .IN1(n27639), .IN2(n116), .IN3(n27647), .IN4(n159), .Q(n3672)
         );
  OA221X1 U3613 ( .IN1(n27591), .IN2(n202), .IN3(n27599), .IN4(n245), .IN5(
        n3673), .Q(n3670) );
  OA22X1 U3614 ( .IN1(n27607), .IN2(n288), .IN3(n27615), .IN4(n331), .Q(n3673)
         );
  OA221X1 U3615 ( .IN1(n27559), .IN2(n374), .IN3(n27567), .IN4(n417), .IN5(
        n3674), .Q(n3669) );
  OA22X1 U3616 ( .IN1(n27575), .IN2(n460), .IN3(n27583), .IN4(n503), .Q(n3674)
         );
  OA221X1 U3617 ( .IN1(n27527), .IN2(n546), .IN3(n27535), .IN4(n589), .IN5(
        n3675), .Q(n3668) );
  OA22X1 U3618 ( .IN1(n27543), .IN2(n632), .IN3(n27551), .IN4(n675), .Q(n3675)
         );
  NAND4X0 U3619 ( .IN1(n3676), .IN2(n3677), .IN3(n3678), .IN4(n3679), .QN(
        n3666) );
  OA221X1 U3620 ( .IN1(n27495), .IN2(n30), .IN3(n27503), .IN4(n73), .IN5(n3680), .Q(n3679) );
  OA22X1 U3621 ( .IN1(n27511), .IN2(n116), .IN3(n27519), .IN4(n159), .Q(n3680)
         );
  OA221X1 U3622 ( .IN1(n27463), .IN2(n202), .IN3(n27471), .IN4(n245), .IN5(
        n3681), .Q(n3678) );
  OA22X1 U3623 ( .IN1(n27479), .IN2(n288), .IN3(n27487), .IN4(n331), .Q(n3681)
         );
  OA221X1 U3624 ( .IN1(n27431), .IN2(n374), .IN3(n27439), .IN4(n417), .IN5(
        n3682), .Q(n3677) );
  OA22X1 U3625 ( .IN1(n27447), .IN2(n460), .IN3(n27455), .IN4(n503), .Q(n3682)
         );
  OA221X1 U3626 ( .IN1(n27399), .IN2(n546), .IN3(n27407), .IN4(n589), .IN5(
        n3683), .Q(n3676) );
  OA22X1 U3627 ( .IN1(n27415), .IN2(n632), .IN3(n27423), .IN4(n675), .Q(n3683)
         );
  NAND4X0 U3628 ( .IN1(n3684), .IN2(n3685), .IN3(n3686), .IN4(n3687), .QN(
        n3664) );
  OA221X1 U3629 ( .IN1(n27367), .IN2(n30), .IN3(n27375), .IN4(n73), .IN5(n3688), .Q(n3687) );
  OA22X1 U3630 ( .IN1(n27383), .IN2(n116), .IN3(n27391), .IN4(n159), .Q(n3688)
         );
  OA221X1 U3631 ( .IN1(n27335), .IN2(n202), .IN3(n27343), .IN4(n245), .IN5(
        n3689), .Q(n3686) );
  OA22X1 U3632 ( .IN1(n27351), .IN2(n288), .IN3(n27359), .IN4(n331), .Q(n3689)
         );
  OA221X1 U3633 ( .IN1(n27303), .IN2(n374), .IN3(n27311), .IN4(n417), .IN5(
        n3690), .Q(n3685) );
  OA22X1 U3634 ( .IN1(n27319), .IN2(n460), .IN3(n27327), .IN4(n503), .Q(n3690)
         );
  OA221X1 U3635 ( .IN1(n27271), .IN2(n546), .IN3(n27279), .IN4(n589), .IN5(
        n3691), .Q(n3684) );
  OA22X1 U3636 ( .IN1(n27287), .IN2(n632), .IN3(n27295), .IN4(n675), .Q(n3691)
         );
  NAND4X0 U3637 ( .IN1(n3692), .IN2(n3693), .IN3(n3694), .IN4(n3695), .QN(
        n3663) );
  OA221X1 U3638 ( .IN1(n27239), .IN2(n30), .IN3(n27247), .IN4(n73), .IN5(n3696), .Q(n3695) );
  OA22X1 U3639 ( .IN1(n27255), .IN2(n116), .IN3(n27263), .IN4(n159), .Q(n3696)
         );
  OA221X1 U3640 ( .IN1(n27207), .IN2(n202), .IN3(n27215), .IN4(n245), .IN5(
        n3697), .Q(n3694) );
  OA22X1 U3641 ( .IN1(n27223), .IN2(n288), .IN3(n27231), .IN4(n331), .Q(n3697)
         );
  OA221X1 U3642 ( .IN1(n27175), .IN2(n374), .IN3(n27183), .IN4(n417), .IN5(
        n3698), .Q(n3693) );
  OA22X1 U3643 ( .IN1(n27191), .IN2(n460), .IN3(n27199), .IN4(n503), .Q(n3698)
         );
  OA221X1 U3644 ( .IN1(n27143), .IN2(n546), .IN3(n27151), .IN4(n589), .IN5(
        n3699), .Q(n3692) );
  OA22X1 U3645 ( .IN1(n27159), .IN2(n632), .IN3(n27167), .IN4(n675), .Q(n3699)
         );
  AO221X1 U3646 ( .IN1(n2328), .IN2(n3700), .IN3(n2330), .IN4(n3701), .IN5(
        n3702), .Q(n3585) );
  AO22X1 U3647 ( .IN1(n2333), .IN2(n3703), .IN3(n2335), .IN4(n3704), .Q(n3702)
         );
  NAND4X0 U3648 ( .IN1(n3705), .IN2(n3706), .IN3(n3707), .IN4(n3708), .QN(
        n3704) );
  OA221X1 U3649 ( .IN1(n27111), .IN2(n30), .IN3(n27119), .IN4(n73), .IN5(n3709), .Q(n3708) );
  OA22X1 U3650 ( .IN1(n27127), .IN2(n116), .IN3(n27135), .IN4(n159), .Q(n3709)
         );
  OA221X1 U3651 ( .IN1(n27079), .IN2(n202), .IN3(n27087), .IN4(n245), .IN5(
        n3710), .Q(n3707) );
  OA22X1 U3652 ( .IN1(n27095), .IN2(n288), .IN3(n27103), .IN4(n331), .Q(n3710)
         );
  OA221X1 U3653 ( .IN1(n27047), .IN2(n374), .IN3(n27055), .IN4(n417), .IN5(
        n3711), .Q(n3706) );
  OA22X1 U3654 ( .IN1(n27063), .IN2(n460), .IN3(n27071), .IN4(n503), .Q(n3711)
         );
  OA221X1 U3655 ( .IN1(n27015), .IN2(n546), .IN3(n27023), .IN4(n589), .IN5(
        n3712), .Q(n3705) );
  OA22X1 U3656 ( .IN1(n27031), .IN2(n632), .IN3(n27039), .IN4(n675), .Q(n3712)
         );
  NAND4X0 U3657 ( .IN1(n3713), .IN2(n3714), .IN3(n3715), .IN4(n3716), .QN(
        n3703) );
  OA221X1 U3658 ( .IN1(n26983), .IN2(n30), .IN3(n26991), .IN4(n73), .IN5(n3717), .Q(n3716) );
  OA22X1 U3659 ( .IN1(n26999), .IN2(n116), .IN3(n27007), .IN4(n159), .Q(n3717)
         );
  OA221X1 U3660 ( .IN1(n26951), .IN2(n202), .IN3(n26959), .IN4(n245), .IN5(
        n3718), .Q(n3715) );
  OA22X1 U3661 ( .IN1(n26967), .IN2(n288), .IN3(n26975), .IN4(n331), .Q(n3718)
         );
  OA221X1 U3662 ( .IN1(n26919), .IN2(n374), .IN3(n26927), .IN4(n417), .IN5(
        n3719), .Q(n3714) );
  OA22X1 U3663 ( .IN1(n26935), .IN2(n460), .IN3(n26943), .IN4(n503), .Q(n3719)
         );
  OA221X1 U3664 ( .IN1(n26887), .IN2(n546), .IN3(n26895), .IN4(n589), .IN5(
        n3720), .Q(n3713) );
  OA22X1 U3665 ( .IN1(n26903), .IN2(n632), .IN3(n26911), .IN4(n675), .Q(n3720)
         );
  NAND4X0 U3666 ( .IN1(n3721), .IN2(n3722), .IN3(n3723), .IN4(n3724), .QN(
        n3701) );
  OA221X1 U3667 ( .IN1(n26855), .IN2(n30), .IN3(n26863), .IN4(n73), .IN5(n3725), .Q(n3724) );
  OA22X1 U3668 ( .IN1(n26871), .IN2(n116), .IN3(n26879), .IN4(n159), .Q(n3725)
         );
  OA221X1 U3669 ( .IN1(n26823), .IN2(n202), .IN3(n26831), .IN4(n245), .IN5(
        n3726), .Q(n3723) );
  OA22X1 U3670 ( .IN1(n26839), .IN2(n288), .IN3(n26847), .IN4(n331), .Q(n3726)
         );
  OA221X1 U3671 ( .IN1(n26791), .IN2(n374), .IN3(n26799), .IN4(n417), .IN5(
        n3727), .Q(n3722) );
  OA22X1 U3672 ( .IN1(n26807), .IN2(n460), .IN3(n26815), .IN4(n503), .Q(n3727)
         );
  OA221X1 U3673 ( .IN1(n26759), .IN2(n546), .IN3(n26767), .IN4(n589), .IN5(
        n3728), .Q(n3721) );
  OA22X1 U3674 ( .IN1(n26775), .IN2(n632), .IN3(n26783), .IN4(n675), .Q(n3728)
         );
  NAND4X0 U3675 ( .IN1(n3729), .IN2(n3730), .IN3(n3731), .IN4(n3732), .QN(
        n3700) );
  OA221X1 U3676 ( .IN1(n26727), .IN2(n30), .IN3(n26735), .IN4(n73), .IN5(n3733), .Q(n3732) );
  OA22X1 U3677 ( .IN1(n26743), .IN2(n116), .IN3(n26751), .IN4(n159), .Q(n3733)
         );
  OA221X1 U3678 ( .IN1(n26695), .IN2(n202), .IN3(n26703), .IN4(n245), .IN5(
        n3734), .Q(n3731) );
  OA22X1 U3679 ( .IN1(n26711), .IN2(n288), .IN3(n26719), .IN4(n331), .Q(n3734)
         );
  OA221X1 U3680 ( .IN1(n26663), .IN2(n374), .IN3(n26671), .IN4(n417), .IN5(
        n3735), .Q(n3730) );
  OA22X1 U3681 ( .IN1(n26679), .IN2(n460), .IN3(n26687), .IN4(n503), .Q(n3735)
         );
  OA221X1 U3682 ( .IN1(n26631), .IN2(n546), .IN3(n26639), .IN4(n589), .IN5(
        n3736), .Q(n3729) );
  OA22X1 U3683 ( .IN1(n26647), .IN2(n632), .IN3(n26655), .IN4(n675), .Q(n3736)
         );
  OR4X1 U3684 ( .IN1(n3737), .IN2(n3738), .IN3(n3739), .IN4(n3740), .Q(n2192)
         );
  AO221X1 U3685 ( .IN1(n2157), .IN2(n3741), .IN3(n2159), .IN4(n3742), .IN5(
        n3743), .Q(n3740) );
  AO22X1 U3686 ( .IN1(n2162), .IN2(n3744), .IN3(n2164), .IN4(n3745), .Q(n3743)
         );
  NAND4X0 U3687 ( .IN1(n3746), .IN2(n3747), .IN3(n3748), .IN4(n3749), .QN(
        n3745) );
  OA221X1 U3688 ( .IN1(n26598), .IN2(n30), .IN3(n26606), .IN4(n73), .IN5(n3750), .Q(n3749) );
  OA22X1 U3689 ( .IN1(n26614), .IN2(n116), .IN3(n26622), .IN4(n159), .Q(n3750)
         );
  OA221X1 U3690 ( .IN1(n26566), .IN2(n202), .IN3(n26574), .IN4(n245), .IN5(
        n3751), .Q(n3748) );
  OA22X1 U3691 ( .IN1(n26582), .IN2(n288), .IN3(n26590), .IN4(n331), .Q(n3751)
         );
  OA221X1 U3692 ( .IN1(n26534), .IN2(n374), .IN3(n26542), .IN4(n417), .IN5(
        n3752), .Q(n3747) );
  OA22X1 U3693 ( .IN1(n26550), .IN2(n460), .IN3(n26558), .IN4(n503), .Q(n3752)
         );
  OA221X1 U3694 ( .IN1(n26502), .IN2(n546), .IN3(n26510), .IN4(n589), .IN5(
        n3753), .Q(n3746) );
  OA22X1 U3695 ( .IN1(n26518), .IN2(n632), .IN3(n26526), .IN4(n675), .Q(n3753)
         );
  NAND4X0 U3696 ( .IN1(n3754), .IN2(n3755), .IN3(n3756), .IN4(n3757), .QN(
        n3744) );
  OA221X1 U3697 ( .IN1(n26470), .IN2(n30), .IN3(n26478), .IN4(n73), .IN5(n3758), .Q(n3757) );
  OA22X1 U3698 ( .IN1(n26486), .IN2(n116), .IN3(n26494), .IN4(n159), .Q(n3758)
         );
  OA221X1 U3699 ( .IN1(n26438), .IN2(n202), .IN3(n26446), .IN4(n245), .IN5(
        n3759), .Q(n3756) );
  OA22X1 U3700 ( .IN1(n26454), .IN2(n288), .IN3(n26462), .IN4(n331), .Q(n3759)
         );
  OA221X1 U3701 ( .IN1(n26406), .IN2(n374), .IN3(n26414), .IN4(n417), .IN5(
        n3760), .Q(n3755) );
  OA22X1 U3702 ( .IN1(n26422), .IN2(n460), .IN3(n26430), .IN4(n503), .Q(n3760)
         );
  OA221X1 U3703 ( .IN1(n26374), .IN2(n546), .IN3(n26382), .IN4(n589), .IN5(
        n3761), .Q(n3754) );
  OA22X1 U3704 ( .IN1(n26390), .IN2(n632), .IN3(n26398), .IN4(n675), .Q(n3761)
         );
  NAND4X0 U3705 ( .IN1(n3762), .IN2(n3763), .IN3(n3764), .IN4(n3765), .QN(
        n3742) );
  OA221X1 U3706 ( .IN1(n26342), .IN2(n30), .IN3(n26350), .IN4(n73), .IN5(n3766), .Q(n3765) );
  OA22X1 U3707 ( .IN1(n26358), .IN2(n116), .IN3(n26366), .IN4(n159), .Q(n3766)
         );
  OA221X1 U3708 ( .IN1(n26310), .IN2(n202), .IN3(n26318), .IN4(n245), .IN5(
        n3767), .Q(n3764) );
  OA22X1 U3709 ( .IN1(n26326), .IN2(n288), .IN3(n26334), .IN4(n331), .Q(n3767)
         );
  OA221X1 U3710 ( .IN1(n26278), .IN2(n374), .IN3(n26286), .IN4(n417), .IN5(
        n3768), .Q(n3763) );
  OA22X1 U3711 ( .IN1(n26294), .IN2(n460), .IN3(n26302), .IN4(n503), .Q(n3768)
         );
  OA221X1 U3712 ( .IN1(n26246), .IN2(n546), .IN3(n26254), .IN4(n589), .IN5(
        n3769), .Q(n3762) );
  OA22X1 U3713 ( .IN1(n26262), .IN2(n632), .IN3(n26270), .IN4(n675), .Q(n3769)
         );
  NAND4X0 U3714 ( .IN1(n3770), .IN2(n3771), .IN3(n3772), .IN4(n3773), .QN(
        n3741) );
  OA221X1 U3715 ( .IN1(n26214), .IN2(n30), .IN3(n26222), .IN4(n73), .IN5(n3774), .Q(n3773) );
  OA22X1 U3716 ( .IN1(n26230), .IN2(n116), .IN3(n26238), .IN4(n159), .Q(n3774)
         );
  OA221X1 U3717 ( .IN1(n26182), .IN2(n202), .IN3(n26190), .IN4(n245), .IN5(
        n3775), .Q(n3772) );
  OA22X1 U3718 ( .IN1(n26198), .IN2(n288), .IN3(n26206), .IN4(n331), .Q(n3775)
         );
  OA221X1 U3719 ( .IN1(n26150), .IN2(n374), .IN3(n26158), .IN4(n417), .IN5(
        n3776), .Q(n3771) );
  OA22X1 U3720 ( .IN1(n26166), .IN2(n460), .IN3(n26174), .IN4(n503), .Q(n3776)
         );
  OA221X1 U3721 ( .IN1(n26118), .IN2(n546), .IN3(n26126), .IN4(n589), .IN5(
        n3777), .Q(n3770) );
  OA22X1 U3722 ( .IN1(n26134), .IN2(n632), .IN3(n26142), .IN4(n675), .Q(n3777)
         );
  AO221X1 U3723 ( .IN1(n2246), .IN2(n3778), .IN3(n2248), .IN4(n3779), .IN5(
        n3780), .Q(n3739) );
  AO22X1 U3724 ( .IN1(n2251), .IN2(n3781), .IN3(n2253), .IN4(n3782), .Q(n3780)
         );
  NAND4X0 U3725 ( .IN1(n3783), .IN2(n3784), .IN3(n3785), .IN4(n3786), .QN(
        n3782) );
  OA221X1 U3726 ( .IN1(n26086), .IN2(n29), .IN3(n26094), .IN4(n72), .IN5(n3787), .Q(n3786) );
  OA22X1 U3727 ( .IN1(n26102), .IN2(n115), .IN3(n26110), .IN4(n158), .Q(n3787)
         );
  OA221X1 U3728 ( .IN1(n26054), .IN2(n201), .IN3(n26062), .IN4(n244), .IN5(
        n3788), .Q(n3785) );
  OA22X1 U3729 ( .IN1(n26070), .IN2(n287), .IN3(n26078), .IN4(n330), .Q(n3788)
         );
  OA221X1 U3730 ( .IN1(n26022), .IN2(n373), .IN3(n26030), .IN4(n416), .IN5(
        n3789), .Q(n3784) );
  OA22X1 U3731 ( .IN1(n26038), .IN2(n459), .IN3(n26046), .IN4(n502), .Q(n3789)
         );
  OA221X1 U3732 ( .IN1(n25990), .IN2(n545), .IN3(n25998), .IN4(n588), .IN5(
        n3790), .Q(n3783) );
  OA22X1 U3733 ( .IN1(n26006), .IN2(n631), .IN3(n26014), .IN4(n674), .Q(n3790)
         );
  NAND4X0 U3734 ( .IN1(n3791), .IN2(n3792), .IN3(n3793), .IN4(n3794), .QN(
        n3781) );
  OA221X1 U3735 ( .IN1(n25958), .IN2(n29), .IN3(n25966), .IN4(n72), .IN5(n3795), .Q(n3794) );
  OA22X1 U3736 ( .IN1(n25974), .IN2(n115), .IN3(n25982), .IN4(n158), .Q(n3795)
         );
  OA221X1 U3737 ( .IN1(n25926), .IN2(n201), .IN3(n25934), .IN4(n244), .IN5(
        n3796), .Q(n3793) );
  OA22X1 U3738 ( .IN1(n25942), .IN2(n287), .IN3(n25950), .IN4(n330), .Q(n3796)
         );
  OA221X1 U3739 ( .IN1(n25894), .IN2(n373), .IN3(n25902), .IN4(n416), .IN5(
        n3797), .Q(n3792) );
  OA22X1 U3740 ( .IN1(n25910), .IN2(n459), .IN3(n25918), .IN4(n502), .Q(n3797)
         );
  OA221X1 U3741 ( .IN1(n25862), .IN2(n545), .IN3(n25870), .IN4(n588), .IN5(
        n3798), .Q(n3791) );
  OA22X1 U3742 ( .IN1(n25878), .IN2(n631), .IN3(n25886), .IN4(n674), .Q(n3798)
         );
  NAND4X0 U3743 ( .IN1(n3799), .IN2(n3800), .IN3(n3801), .IN4(n3802), .QN(
        n3779) );
  OA221X1 U3744 ( .IN1(n25830), .IN2(n29), .IN3(n25838), .IN4(n72), .IN5(n3803), .Q(n3802) );
  OA22X1 U3745 ( .IN1(n25846), .IN2(n115), .IN3(n25854), .IN4(n158), .Q(n3803)
         );
  OA221X1 U3746 ( .IN1(n25798), .IN2(n201), .IN3(n25806), .IN4(n244), .IN5(
        n3804), .Q(n3801) );
  OA22X1 U3747 ( .IN1(n25814), .IN2(n287), .IN3(n25822), .IN4(n330), .Q(n3804)
         );
  OA221X1 U3748 ( .IN1(n25766), .IN2(n373), .IN3(n25774), .IN4(n416), .IN5(
        n3805), .Q(n3800) );
  OA22X1 U3749 ( .IN1(n25782), .IN2(n459), .IN3(n25790), .IN4(n502), .Q(n3805)
         );
  OA221X1 U3750 ( .IN1(n25734), .IN2(n545), .IN3(n25742), .IN4(n588), .IN5(
        n3806), .Q(n3799) );
  OA22X1 U3751 ( .IN1(n25750), .IN2(n631), .IN3(n25758), .IN4(n674), .Q(n3806)
         );
  NAND4X0 U3752 ( .IN1(n3807), .IN2(n3808), .IN3(n3809), .IN4(n3810), .QN(
        n3778) );
  OA221X1 U3753 ( .IN1(n25702), .IN2(n29), .IN3(n25710), .IN4(n72), .IN5(n3811), .Q(n3810) );
  OA22X1 U3754 ( .IN1(n25718), .IN2(n115), .IN3(n25726), .IN4(n158), .Q(n3811)
         );
  OA221X1 U3755 ( .IN1(n25670), .IN2(n201), .IN3(n25678), .IN4(n244), .IN5(
        n3812), .Q(n3809) );
  OA22X1 U3756 ( .IN1(n25686), .IN2(n287), .IN3(n25694), .IN4(n330), .Q(n3812)
         );
  OA221X1 U3757 ( .IN1(n25638), .IN2(n373), .IN3(n25646), .IN4(n416), .IN5(
        n3813), .Q(n3808) );
  OA22X1 U3758 ( .IN1(n25654), .IN2(n459), .IN3(n25662), .IN4(n502), .Q(n3813)
         );
  OA221X1 U3759 ( .IN1(n25606), .IN2(n545), .IN3(n25614), .IN4(n588), .IN5(
        n3814), .Q(n3807) );
  OA22X1 U3760 ( .IN1(n25622), .IN2(n631), .IN3(n25630), .IN4(n674), .Q(n3814)
         );
  AO221X1 U3761 ( .IN1(n2287), .IN2(n3815), .IN3(n2289), .IN4(n3816), .IN5(
        n3817), .Q(n3738) );
  AO22X1 U3762 ( .IN1(n2292), .IN2(n3818), .IN3(n2294), .IN4(n3819), .Q(n3817)
         );
  NAND4X0 U3763 ( .IN1(n3820), .IN2(n3821), .IN3(n3822), .IN4(n3823), .QN(
        n3819) );
  OA221X1 U3764 ( .IN1(n27622), .IN2(n29), .IN3(n27630), .IN4(n72), .IN5(n3824), .Q(n3823) );
  OA22X1 U3765 ( .IN1(n27638), .IN2(n115), .IN3(n27646), .IN4(n158), .Q(n3824)
         );
  OA221X1 U3766 ( .IN1(n27590), .IN2(n201), .IN3(n27598), .IN4(n244), .IN5(
        n3825), .Q(n3822) );
  OA22X1 U3767 ( .IN1(n27606), .IN2(n287), .IN3(n27614), .IN4(n330), .Q(n3825)
         );
  OA221X1 U3768 ( .IN1(n27558), .IN2(n373), .IN3(n27566), .IN4(n416), .IN5(
        n3826), .Q(n3821) );
  OA22X1 U3769 ( .IN1(n27574), .IN2(n459), .IN3(n27582), .IN4(n502), .Q(n3826)
         );
  OA221X1 U3770 ( .IN1(n27526), .IN2(n545), .IN3(n27534), .IN4(n588), .IN5(
        n3827), .Q(n3820) );
  OA22X1 U3771 ( .IN1(n27542), .IN2(n631), .IN3(n27550), .IN4(n674), .Q(n3827)
         );
  NAND4X0 U3772 ( .IN1(n3828), .IN2(n3829), .IN3(n3830), .IN4(n3831), .QN(
        n3818) );
  OA221X1 U3773 ( .IN1(n27494), .IN2(n29), .IN3(n27502), .IN4(n72), .IN5(n3832), .Q(n3831) );
  OA22X1 U3774 ( .IN1(n27510), .IN2(n115), .IN3(n27518), .IN4(n158), .Q(n3832)
         );
  OA221X1 U3775 ( .IN1(n27462), .IN2(n201), .IN3(n27470), .IN4(n244), .IN5(
        n3833), .Q(n3830) );
  OA22X1 U3776 ( .IN1(n27478), .IN2(n287), .IN3(n27486), .IN4(n330), .Q(n3833)
         );
  OA221X1 U3777 ( .IN1(n27430), .IN2(n373), .IN3(n27438), .IN4(n416), .IN5(
        n3834), .Q(n3829) );
  OA22X1 U3778 ( .IN1(n27446), .IN2(n459), .IN3(n27454), .IN4(n502), .Q(n3834)
         );
  OA221X1 U3779 ( .IN1(n27398), .IN2(n545), .IN3(n27406), .IN4(n588), .IN5(
        n3835), .Q(n3828) );
  OA22X1 U3780 ( .IN1(n27414), .IN2(n631), .IN3(n27422), .IN4(n674), .Q(n3835)
         );
  NAND4X0 U3781 ( .IN1(n3836), .IN2(n3837), .IN3(n3838), .IN4(n3839), .QN(
        n3816) );
  OA221X1 U3782 ( .IN1(n27366), .IN2(n29), .IN3(n27374), .IN4(n72), .IN5(n3840), .Q(n3839) );
  OA22X1 U3783 ( .IN1(n27382), .IN2(n115), .IN3(n27390), .IN4(n158), .Q(n3840)
         );
  OA221X1 U3784 ( .IN1(n27334), .IN2(n201), .IN3(n27342), .IN4(n244), .IN5(
        n3841), .Q(n3838) );
  OA22X1 U3785 ( .IN1(n27350), .IN2(n287), .IN3(n27358), .IN4(n330), .Q(n3841)
         );
  OA221X1 U3786 ( .IN1(n27302), .IN2(n373), .IN3(n27310), .IN4(n416), .IN5(
        n3842), .Q(n3837) );
  OA22X1 U3787 ( .IN1(n27318), .IN2(n459), .IN3(n27326), .IN4(n502), .Q(n3842)
         );
  OA221X1 U3788 ( .IN1(n27270), .IN2(n545), .IN3(n27278), .IN4(n588), .IN5(
        n3843), .Q(n3836) );
  OA22X1 U3789 ( .IN1(n27286), .IN2(n631), .IN3(n27294), .IN4(n674), .Q(n3843)
         );
  NAND4X0 U3790 ( .IN1(n3844), .IN2(n3845), .IN3(n3846), .IN4(n3847), .QN(
        n3815) );
  OA221X1 U3791 ( .IN1(n27238), .IN2(n29), .IN3(n27246), .IN4(n72), .IN5(n3848), .Q(n3847) );
  OA22X1 U3792 ( .IN1(n27254), .IN2(n115), .IN3(n27262), .IN4(n158), .Q(n3848)
         );
  OA221X1 U3793 ( .IN1(n27206), .IN2(n201), .IN3(n27214), .IN4(n244), .IN5(
        n3849), .Q(n3846) );
  OA22X1 U3794 ( .IN1(n27222), .IN2(n287), .IN3(n27230), .IN4(n330), .Q(n3849)
         );
  OA221X1 U3795 ( .IN1(n27174), .IN2(n373), .IN3(n27182), .IN4(n416), .IN5(
        n3850), .Q(n3845) );
  OA22X1 U3796 ( .IN1(n27190), .IN2(n459), .IN3(n27198), .IN4(n502), .Q(n3850)
         );
  OA221X1 U3797 ( .IN1(n27142), .IN2(n545), .IN3(n27150), .IN4(n588), .IN5(
        n3851), .Q(n3844) );
  OA22X1 U3798 ( .IN1(n27158), .IN2(n631), .IN3(n27166), .IN4(n674), .Q(n3851)
         );
  AO221X1 U3799 ( .IN1(n2328), .IN2(n3852), .IN3(n2330), .IN4(n3853), .IN5(
        n3854), .Q(n3737) );
  AO22X1 U3800 ( .IN1(n2333), .IN2(n3855), .IN3(n2335), .IN4(n3856), .Q(n3854)
         );
  NAND4X0 U3801 ( .IN1(n3857), .IN2(n3858), .IN3(n3859), .IN4(n3860), .QN(
        n3856) );
  OA221X1 U3802 ( .IN1(n27110), .IN2(n29), .IN3(n27118), .IN4(n72), .IN5(n3861), .Q(n3860) );
  OA22X1 U3803 ( .IN1(n27126), .IN2(n115), .IN3(n27134), .IN4(n158), .Q(n3861)
         );
  OA221X1 U3804 ( .IN1(n27078), .IN2(n201), .IN3(n27086), .IN4(n244), .IN5(
        n3862), .Q(n3859) );
  OA22X1 U3805 ( .IN1(n27094), .IN2(n287), .IN3(n27102), .IN4(n330), .Q(n3862)
         );
  OA221X1 U3806 ( .IN1(n27046), .IN2(n373), .IN3(n27054), .IN4(n416), .IN5(
        n3863), .Q(n3858) );
  OA22X1 U3807 ( .IN1(n27062), .IN2(n459), .IN3(n27070), .IN4(n502), .Q(n3863)
         );
  OA221X1 U3808 ( .IN1(n27014), .IN2(n545), .IN3(n27022), .IN4(n588), .IN5(
        n3864), .Q(n3857) );
  OA22X1 U3809 ( .IN1(n27030), .IN2(n631), .IN3(n27038), .IN4(n674), .Q(n3864)
         );
  NAND4X0 U3810 ( .IN1(n3865), .IN2(n3866), .IN3(n3867), .IN4(n3868), .QN(
        n3855) );
  OA221X1 U3811 ( .IN1(n26982), .IN2(n29), .IN3(n26990), .IN4(n72), .IN5(n3869), .Q(n3868) );
  OA22X1 U3812 ( .IN1(n26998), .IN2(n115), .IN3(n27006), .IN4(n158), .Q(n3869)
         );
  OA221X1 U3813 ( .IN1(n26950), .IN2(n201), .IN3(n26958), .IN4(n244), .IN5(
        n3870), .Q(n3867) );
  OA22X1 U3814 ( .IN1(n26966), .IN2(n287), .IN3(n26974), .IN4(n330), .Q(n3870)
         );
  OA221X1 U3815 ( .IN1(n26918), .IN2(n373), .IN3(n26926), .IN4(n416), .IN5(
        n3871), .Q(n3866) );
  OA22X1 U3816 ( .IN1(n26934), .IN2(n459), .IN3(n26942), .IN4(n502), .Q(n3871)
         );
  OA221X1 U3817 ( .IN1(n26886), .IN2(n545), .IN3(n26894), .IN4(n588), .IN5(
        n3872), .Q(n3865) );
  OA22X1 U3818 ( .IN1(n26902), .IN2(n631), .IN3(n26910), .IN4(n674), .Q(n3872)
         );
  NAND4X0 U3819 ( .IN1(n3873), .IN2(n3874), .IN3(n3875), .IN4(n3876), .QN(
        n3853) );
  OA221X1 U3820 ( .IN1(n26854), .IN2(n29), .IN3(n26862), .IN4(n72), .IN5(n3877), .Q(n3876) );
  OA22X1 U3821 ( .IN1(n26870), .IN2(n115), .IN3(n26878), .IN4(n158), .Q(n3877)
         );
  OA221X1 U3822 ( .IN1(n26822), .IN2(n201), .IN3(n26830), .IN4(n244), .IN5(
        n3878), .Q(n3875) );
  OA22X1 U3823 ( .IN1(n26838), .IN2(n287), .IN3(n26846), .IN4(n330), .Q(n3878)
         );
  OA221X1 U3824 ( .IN1(n26790), .IN2(n373), .IN3(n26798), .IN4(n416), .IN5(
        n3879), .Q(n3874) );
  OA22X1 U3825 ( .IN1(n26806), .IN2(n459), .IN3(n26814), .IN4(n502), .Q(n3879)
         );
  OA221X1 U3826 ( .IN1(n26758), .IN2(n545), .IN3(n26766), .IN4(n588), .IN5(
        n3880), .Q(n3873) );
  OA22X1 U3827 ( .IN1(n26774), .IN2(n631), .IN3(n26782), .IN4(n674), .Q(n3880)
         );
  NAND4X0 U3828 ( .IN1(n3881), .IN2(n3882), .IN3(n3883), .IN4(n3884), .QN(
        n3852) );
  OA221X1 U3829 ( .IN1(n26726), .IN2(n29), .IN3(n26734), .IN4(n72), .IN5(n3885), .Q(n3884) );
  OA22X1 U3830 ( .IN1(n26742), .IN2(n115), .IN3(n26750), .IN4(n158), .Q(n3885)
         );
  OA221X1 U3831 ( .IN1(n26694), .IN2(n201), .IN3(n26702), .IN4(n244), .IN5(
        n3886), .Q(n3883) );
  OA22X1 U3832 ( .IN1(n26710), .IN2(n287), .IN3(n26718), .IN4(n330), .Q(n3886)
         );
  OA221X1 U3833 ( .IN1(n26662), .IN2(n373), .IN3(n26670), .IN4(n416), .IN5(
        n3887), .Q(n3882) );
  OA22X1 U3834 ( .IN1(n26678), .IN2(n459), .IN3(n26686), .IN4(n502), .Q(n3887)
         );
  OA221X1 U3835 ( .IN1(n26630), .IN2(n545), .IN3(n26638), .IN4(n588), .IN5(
        n3888), .Q(n3881) );
  OA22X1 U3836 ( .IN1(n26646), .IN2(n631), .IN3(n26654), .IN4(n674), .Q(n3888)
         );
  OR4X1 U3837 ( .IN1(n3889), .IN2(n3890), .IN3(n3891), .IN4(n3892), .Q(n2191)
         );
  AO221X1 U3838 ( .IN1(n2157), .IN2(n3893), .IN3(n2159), .IN4(n3894), .IN5(
        n3895), .Q(n3892) );
  AO22X1 U3839 ( .IN1(n2162), .IN2(n3896), .IN3(n2164), .IN4(n3897), .Q(n3895)
         );
  NAND4X0 U3840 ( .IN1(n3898), .IN2(n3899), .IN3(n3900), .IN4(n3901), .QN(
        n3897) );
  OA221X1 U3841 ( .IN1(n26597), .IN2(n28), .IN3(n26605), .IN4(n71), .IN5(n3902), .Q(n3901) );
  OA22X1 U3842 ( .IN1(n26613), .IN2(n114), .IN3(n26621), .IN4(n157), .Q(n3902)
         );
  OA221X1 U3843 ( .IN1(n26565), .IN2(n200), .IN3(n26573), .IN4(n243), .IN5(
        n3903), .Q(n3900) );
  OA22X1 U3844 ( .IN1(n26581), .IN2(n286), .IN3(n26589), .IN4(n329), .Q(n3903)
         );
  OA221X1 U3845 ( .IN1(n26533), .IN2(n372), .IN3(n26541), .IN4(n415), .IN5(
        n3904), .Q(n3899) );
  OA22X1 U3846 ( .IN1(n26549), .IN2(n458), .IN3(n26557), .IN4(n501), .Q(n3904)
         );
  OA221X1 U3847 ( .IN1(n26501), .IN2(n544), .IN3(n26509), .IN4(n587), .IN5(
        n3905), .Q(n3898) );
  OA22X1 U3848 ( .IN1(n26517), .IN2(n630), .IN3(n26525), .IN4(n673), .Q(n3905)
         );
  NAND4X0 U3849 ( .IN1(n3906), .IN2(n3907), .IN3(n3908), .IN4(n3909), .QN(
        n3896) );
  OA221X1 U3850 ( .IN1(n26469), .IN2(n28), .IN3(n26477), .IN4(n71), .IN5(n3910), .Q(n3909) );
  OA22X1 U3851 ( .IN1(n26485), .IN2(n114), .IN3(n26493), .IN4(n157), .Q(n3910)
         );
  OA221X1 U3852 ( .IN1(n26437), .IN2(n200), .IN3(n26445), .IN4(n243), .IN5(
        n3911), .Q(n3908) );
  OA22X1 U3853 ( .IN1(n26453), .IN2(n286), .IN3(n26461), .IN4(n329), .Q(n3911)
         );
  OA221X1 U3854 ( .IN1(n26405), .IN2(n372), .IN3(n26413), .IN4(n415), .IN5(
        n3912), .Q(n3907) );
  OA22X1 U3855 ( .IN1(n26421), .IN2(n458), .IN3(n26429), .IN4(n501), .Q(n3912)
         );
  OA221X1 U3856 ( .IN1(n26373), .IN2(n544), .IN3(n26381), .IN4(n587), .IN5(
        n3913), .Q(n3906) );
  OA22X1 U3857 ( .IN1(n26389), .IN2(n630), .IN3(n26397), .IN4(n673), .Q(n3913)
         );
  NAND4X0 U3858 ( .IN1(n3914), .IN2(n3915), .IN3(n3916), .IN4(n3917), .QN(
        n3894) );
  OA221X1 U3859 ( .IN1(n26341), .IN2(n28), .IN3(n26349), .IN4(n71), .IN5(n3918), .Q(n3917) );
  OA22X1 U3860 ( .IN1(n26357), .IN2(n114), .IN3(n26365), .IN4(n157), .Q(n3918)
         );
  OA221X1 U3861 ( .IN1(n26309), .IN2(n200), .IN3(n26317), .IN4(n243), .IN5(
        n3919), .Q(n3916) );
  OA22X1 U3862 ( .IN1(n26325), .IN2(n286), .IN3(n26333), .IN4(n329), .Q(n3919)
         );
  OA221X1 U3863 ( .IN1(n26277), .IN2(n372), .IN3(n26285), .IN4(n415), .IN5(
        n3920), .Q(n3915) );
  OA22X1 U3864 ( .IN1(n26293), .IN2(n458), .IN3(n26301), .IN4(n501), .Q(n3920)
         );
  OA221X1 U3865 ( .IN1(n26245), .IN2(n544), .IN3(n26253), .IN4(n587), .IN5(
        n3921), .Q(n3914) );
  OA22X1 U3866 ( .IN1(n26261), .IN2(n630), .IN3(n26269), .IN4(n673), .Q(n3921)
         );
  NAND4X0 U3867 ( .IN1(n3922), .IN2(n3923), .IN3(n3924), .IN4(n3925), .QN(
        n3893) );
  OA221X1 U3868 ( .IN1(n26213), .IN2(n28), .IN3(n26221), .IN4(n71), .IN5(n3926), .Q(n3925) );
  OA22X1 U3869 ( .IN1(n26229), .IN2(n114), .IN3(n26237), .IN4(n157), .Q(n3926)
         );
  OA221X1 U3870 ( .IN1(n26181), .IN2(n200), .IN3(n26189), .IN4(n243), .IN5(
        n3927), .Q(n3924) );
  OA22X1 U3871 ( .IN1(n26197), .IN2(n286), .IN3(n26205), .IN4(n329), .Q(n3927)
         );
  OA221X1 U3872 ( .IN1(n26149), .IN2(n372), .IN3(n26157), .IN4(n415), .IN5(
        n3928), .Q(n3923) );
  OA22X1 U3873 ( .IN1(n26165), .IN2(n458), .IN3(n26173), .IN4(n501), .Q(n3928)
         );
  OA221X1 U3874 ( .IN1(n26117), .IN2(n544), .IN3(n26125), .IN4(n587), .IN5(
        n3929), .Q(n3922) );
  OA22X1 U3875 ( .IN1(n26133), .IN2(n630), .IN3(n26141), .IN4(n673), .Q(n3929)
         );
  AO221X1 U3876 ( .IN1(n2246), .IN2(n3930), .IN3(n2248), .IN4(n3931), .IN5(
        n3932), .Q(n3891) );
  AO22X1 U3877 ( .IN1(n2251), .IN2(n3933), .IN3(n2253), .IN4(n3934), .Q(n3932)
         );
  NAND4X0 U3878 ( .IN1(n3935), .IN2(n3936), .IN3(n3937), .IN4(n3938), .QN(
        n3934) );
  OA221X1 U3879 ( .IN1(n26085), .IN2(n28), .IN3(n26093), .IN4(n71), .IN5(n3939), .Q(n3938) );
  OA22X1 U3880 ( .IN1(n26101), .IN2(n114), .IN3(n26109), .IN4(n157), .Q(n3939)
         );
  OA221X1 U3881 ( .IN1(n26053), .IN2(n200), .IN3(n26061), .IN4(n243), .IN5(
        n3940), .Q(n3937) );
  OA22X1 U3882 ( .IN1(n26069), .IN2(n286), .IN3(n26077), .IN4(n329), .Q(n3940)
         );
  OA221X1 U3883 ( .IN1(n26021), .IN2(n372), .IN3(n26029), .IN4(n415), .IN5(
        n3941), .Q(n3936) );
  OA22X1 U3884 ( .IN1(n26037), .IN2(n458), .IN3(n26045), .IN4(n501), .Q(n3941)
         );
  OA221X1 U3885 ( .IN1(n25989), .IN2(n544), .IN3(n25997), .IN4(n587), .IN5(
        n3942), .Q(n3935) );
  OA22X1 U3886 ( .IN1(n26005), .IN2(n630), .IN3(n26013), .IN4(n673), .Q(n3942)
         );
  NAND4X0 U3887 ( .IN1(n3943), .IN2(n3944), .IN3(n3945), .IN4(n3946), .QN(
        n3933) );
  OA221X1 U3888 ( .IN1(n25957), .IN2(n28), .IN3(n25965), .IN4(n71), .IN5(n3947), .Q(n3946) );
  OA22X1 U3889 ( .IN1(n25973), .IN2(n114), .IN3(n25981), .IN4(n157), .Q(n3947)
         );
  OA221X1 U3890 ( .IN1(n25925), .IN2(n200), .IN3(n25933), .IN4(n243), .IN5(
        n3948), .Q(n3945) );
  OA22X1 U3891 ( .IN1(n25941), .IN2(n286), .IN3(n25949), .IN4(n329), .Q(n3948)
         );
  OA221X1 U3892 ( .IN1(n25893), .IN2(n372), .IN3(n25901), .IN4(n415), .IN5(
        n3949), .Q(n3944) );
  OA22X1 U3893 ( .IN1(n25909), .IN2(n458), .IN3(n25917), .IN4(n501), .Q(n3949)
         );
  OA221X1 U3894 ( .IN1(n25861), .IN2(n544), .IN3(n25869), .IN4(n587), .IN5(
        n3950), .Q(n3943) );
  OA22X1 U3895 ( .IN1(n25877), .IN2(n630), .IN3(n25885), .IN4(n673), .Q(n3950)
         );
  NAND4X0 U3896 ( .IN1(n3951), .IN2(n3952), .IN3(n3953), .IN4(n3954), .QN(
        n3931) );
  OA221X1 U3897 ( .IN1(n25829), .IN2(n28), .IN3(n25837), .IN4(n71), .IN5(n3955), .Q(n3954) );
  OA22X1 U3898 ( .IN1(n25845), .IN2(n114), .IN3(n25853), .IN4(n157), .Q(n3955)
         );
  OA221X1 U3899 ( .IN1(n25797), .IN2(n200), .IN3(n25805), .IN4(n243), .IN5(
        n3956), .Q(n3953) );
  OA22X1 U3900 ( .IN1(n25813), .IN2(n286), .IN3(n25821), .IN4(n329), .Q(n3956)
         );
  OA221X1 U3901 ( .IN1(n25765), .IN2(n372), .IN3(n25773), .IN4(n415), .IN5(
        n3957), .Q(n3952) );
  OA22X1 U3902 ( .IN1(n25781), .IN2(n458), .IN3(n25789), .IN4(n501), .Q(n3957)
         );
  OA221X1 U3903 ( .IN1(n25733), .IN2(n544), .IN3(n25741), .IN4(n587), .IN5(
        n3958), .Q(n3951) );
  OA22X1 U3904 ( .IN1(n25749), .IN2(n630), .IN3(n25757), .IN4(n673), .Q(n3958)
         );
  NAND4X0 U3905 ( .IN1(n3959), .IN2(n3960), .IN3(n3961), .IN4(n3962), .QN(
        n3930) );
  OA221X1 U3906 ( .IN1(n25701), .IN2(n28), .IN3(n25709), .IN4(n71), .IN5(n3963), .Q(n3962) );
  OA22X1 U3907 ( .IN1(n25717), .IN2(n114), .IN3(n25725), .IN4(n157), .Q(n3963)
         );
  OA221X1 U3908 ( .IN1(n25669), .IN2(n200), .IN3(n25677), .IN4(n243), .IN5(
        n3964), .Q(n3961) );
  OA22X1 U3909 ( .IN1(n25685), .IN2(n286), .IN3(n25693), .IN4(n329), .Q(n3964)
         );
  OA221X1 U3910 ( .IN1(n25637), .IN2(n372), .IN3(n25645), .IN4(n415), .IN5(
        n3965), .Q(n3960) );
  OA22X1 U3911 ( .IN1(n25653), .IN2(n458), .IN3(n25661), .IN4(n501), .Q(n3965)
         );
  OA221X1 U3912 ( .IN1(n25605), .IN2(n544), .IN3(n25613), .IN4(n587), .IN5(
        n3966), .Q(n3959) );
  OA22X1 U3913 ( .IN1(n25621), .IN2(n630), .IN3(n25629), .IN4(n673), .Q(n3966)
         );
  AO221X1 U3914 ( .IN1(n2287), .IN2(n3967), .IN3(n2289), .IN4(n3968), .IN5(
        n3969), .Q(n3890) );
  AO22X1 U3915 ( .IN1(n2292), .IN2(n3970), .IN3(n2294), .IN4(n3971), .Q(n3969)
         );
  NAND4X0 U3916 ( .IN1(n3972), .IN2(n3973), .IN3(n3974), .IN4(n3975), .QN(
        n3971) );
  OA221X1 U3917 ( .IN1(n27621), .IN2(n28), .IN3(n27629), .IN4(n71), .IN5(n3976), .Q(n3975) );
  OA22X1 U3918 ( .IN1(n27637), .IN2(n114), .IN3(n27645), .IN4(n157), .Q(n3976)
         );
  OA221X1 U3919 ( .IN1(n27589), .IN2(n200), .IN3(n27597), .IN4(n243), .IN5(
        n3977), .Q(n3974) );
  OA22X1 U3920 ( .IN1(n27605), .IN2(n286), .IN3(n27613), .IN4(n329), .Q(n3977)
         );
  OA221X1 U3921 ( .IN1(n27557), .IN2(n372), .IN3(n27565), .IN4(n415), .IN5(
        n3978), .Q(n3973) );
  OA22X1 U3922 ( .IN1(n27573), .IN2(n458), .IN3(n27581), .IN4(n501), .Q(n3978)
         );
  OA221X1 U3923 ( .IN1(n27525), .IN2(n544), .IN3(n27533), .IN4(n587), .IN5(
        n3979), .Q(n3972) );
  OA22X1 U3924 ( .IN1(n27541), .IN2(n630), .IN3(n27549), .IN4(n673), .Q(n3979)
         );
  NAND4X0 U3925 ( .IN1(n3980), .IN2(n3981), .IN3(n3982), .IN4(n3983), .QN(
        n3970) );
  OA221X1 U3926 ( .IN1(n27493), .IN2(n28), .IN3(n27501), .IN4(n71), .IN5(n3984), .Q(n3983) );
  OA22X1 U3927 ( .IN1(n27509), .IN2(n114), .IN3(n27517), .IN4(n157), .Q(n3984)
         );
  OA221X1 U3928 ( .IN1(n27461), .IN2(n200), .IN3(n27469), .IN4(n243), .IN5(
        n3985), .Q(n3982) );
  OA22X1 U3929 ( .IN1(n27477), .IN2(n286), .IN3(n27485), .IN4(n329), .Q(n3985)
         );
  OA221X1 U3930 ( .IN1(n27429), .IN2(n372), .IN3(n27437), .IN4(n415), .IN5(
        n3986), .Q(n3981) );
  OA22X1 U3931 ( .IN1(n27445), .IN2(n458), .IN3(n27453), .IN4(n501), .Q(n3986)
         );
  OA221X1 U3932 ( .IN1(n27397), .IN2(n544), .IN3(n27405), .IN4(n587), .IN5(
        n3987), .Q(n3980) );
  OA22X1 U3933 ( .IN1(n27413), .IN2(n630), .IN3(n27421), .IN4(n673), .Q(n3987)
         );
  NAND4X0 U3934 ( .IN1(n3988), .IN2(n3989), .IN3(n3990), .IN4(n3991), .QN(
        n3968) );
  OA221X1 U3935 ( .IN1(n27365), .IN2(n28), .IN3(n27373), .IN4(n71), .IN5(n3992), .Q(n3991) );
  OA22X1 U3936 ( .IN1(n27381), .IN2(n114), .IN3(n27389), .IN4(n157), .Q(n3992)
         );
  OA221X1 U3937 ( .IN1(n27333), .IN2(n200), .IN3(n27341), .IN4(n243), .IN5(
        n3993), .Q(n3990) );
  OA22X1 U3938 ( .IN1(n27349), .IN2(n286), .IN3(n27357), .IN4(n329), .Q(n3993)
         );
  OA221X1 U3939 ( .IN1(n27301), .IN2(n372), .IN3(n27309), .IN4(n415), .IN5(
        n3994), .Q(n3989) );
  OA22X1 U3940 ( .IN1(n27317), .IN2(n458), .IN3(n27325), .IN4(n501), .Q(n3994)
         );
  OA221X1 U3941 ( .IN1(n27269), .IN2(n544), .IN3(n27277), .IN4(n587), .IN5(
        n3995), .Q(n3988) );
  OA22X1 U3942 ( .IN1(n27285), .IN2(n630), .IN3(n27293), .IN4(n673), .Q(n3995)
         );
  NAND4X0 U3943 ( .IN1(n3996), .IN2(n3997), .IN3(n3998), .IN4(n3999), .QN(
        n3967) );
  OA221X1 U3944 ( .IN1(n27237), .IN2(n28), .IN3(n27245), .IN4(n71), .IN5(n4000), .Q(n3999) );
  OA22X1 U3945 ( .IN1(n27253), .IN2(n114), .IN3(n27261), .IN4(n157), .Q(n4000)
         );
  OA221X1 U3946 ( .IN1(n27205), .IN2(n200), .IN3(n27213), .IN4(n243), .IN5(
        n4001), .Q(n3998) );
  OA22X1 U3947 ( .IN1(n27221), .IN2(n286), .IN3(n27229), .IN4(n329), .Q(n4001)
         );
  OA221X1 U3948 ( .IN1(n27173), .IN2(n372), .IN3(n27181), .IN4(n415), .IN5(
        n4002), .Q(n3997) );
  OA22X1 U3949 ( .IN1(n27189), .IN2(n458), .IN3(n27197), .IN4(n501), .Q(n4002)
         );
  OA221X1 U3950 ( .IN1(n27141), .IN2(n544), .IN3(n27149), .IN4(n587), .IN5(
        n4003), .Q(n3996) );
  OA22X1 U3951 ( .IN1(n27157), .IN2(n630), .IN3(n27165), .IN4(n673), .Q(n4003)
         );
  AO221X1 U3952 ( .IN1(n2328), .IN2(n4004), .IN3(n2330), .IN4(n4005), .IN5(
        n4006), .Q(n3889) );
  AO22X1 U3953 ( .IN1(n2333), .IN2(n4007), .IN3(n2335), .IN4(n4008), .Q(n4006)
         );
  NAND4X0 U3954 ( .IN1(n4009), .IN2(n4010), .IN3(n4011), .IN4(n4012), .QN(
        n4008) );
  OA221X1 U3955 ( .IN1(n27109), .IN2(n27), .IN3(n27117), .IN4(n70), .IN5(n4013), .Q(n4012) );
  OA22X1 U3956 ( .IN1(n27125), .IN2(n113), .IN3(n27133), .IN4(n156), .Q(n4013)
         );
  OA221X1 U3957 ( .IN1(n27077), .IN2(n199), .IN3(n27085), .IN4(n242), .IN5(
        n4014), .Q(n4011) );
  OA22X1 U3958 ( .IN1(n27093), .IN2(n285), .IN3(n27101), .IN4(n328), .Q(n4014)
         );
  OA221X1 U3959 ( .IN1(n27045), .IN2(n371), .IN3(n27053), .IN4(n414), .IN5(
        n4015), .Q(n4010) );
  OA22X1 U3960 ( .IN1(n27061), .IN2(n457), .IN3(n27069), .IN4(n500), .Q(n4015)
         );
  OA221X1 U3961 ( .IN1(n27013), .IN2(n543), .IN3(n27021), .IN4(n586), .IN5(
        n4016), .Q(n4009) );
  OA22X1 U3962 ( .IN1(n27029), .IN2(n629), .IN3(n27037), .IN4(n672), .Q(n4016)
         );
  NAND4X0 U3963 ( .IN1(n4017), .IN2(n4018), .IN3(n4019), .IN4(n4020), .QN(
        n4007) );
  OA221X1 U3964 ( .IN1(n26981), .IN2(n27), .IN3(n26989), .IN4(n70), .IN5(n4021), .Q(n4020) );
  OA22X1 U3965 ( .IN1(n26997), .IN2(n113), .IN3(n27005), .IN4(n156), .Q(n4021)
         );
  OA221X1 U3966 ( .IN1(n26949), .IN2(n199), .IN3(n26957), .IN4(n242), .IN5(
        n4022), .Q(n4019) );
  OA22X1 U3967 ( .IN1(n26965), .IN2(n285), .IN3(n26973), .IN4(n328), .Q(n4022)
         );
  OA221X1 U3968 ( .IN1(n26917), .IN2(n371), .IN3(n26925), .IN4(n414), .IN5(
        n4023), .Q(n4018) );
  OA22X1 U3969 ( .IN1(n26933), .IN2(n457), .IN3(n26941), .IN4(n500), .Q(n4023)
         );
  OA221X1 U3970 ( .IN1(n26885), .IN2(n543), .IN3(n26893), .IN4(n586), .IN5(
        n4024), .Q(n4017) );
  OA22X1 U3971 ( .IN1(n26901), .IN2(n629), .IN3(n26909), .IN4(n672), .Q(n4024)
         );
  NAND4X0 U3972 ( .IN1(n4025), .IN2(n4026), .IN3(n4027), .IN4(n4028), .QN(
        n4005) );
  OA221X1 U3973 ( .IN1(n26853), .IN2(n27), .IN3(n26861), .IN4(n70), .IN5(n4029), .Q(n4028) );
  OA22X1 U3974 ( .IN1(n26869), .IN2(n113), .IN3(n26877), .IN4(n156), .Q(n4029)
         );
  OA221X1 U3975 ( .IN1(n26821), .IN2(n199), .IN3(n26829), .IN4(n242), .IN5(
        n4030), .Q(n4027) );
  OA22X1 U3976 ( .IN1(n26837), .IN2(n285), .IN3(n26845), .IN4(n328), .Q(n4030)
         );
  OA221X1 U3977 ( .IN1(n26789), .IN2(n371), .IN3(n26797), .IN4(n414), .IN5(
        n4031), .Q(n4026) );
  OA22X1 U3978 ( .IN1(n26805), .IN2(n457), .IN3(n26813), .IN4(n500), .Q(n4031)
         );
  OA221X1 U3979 ( .IN1(n26757), .IN2(n543), .IN3(n26765), .IN4(n586), .IN5(
        n4032), .Q(n4025) );
  OA22X1 U3980 ( .IN1(n26773), .IN2(n629), .IN3(n26781), .IN4(n672), .Q(n4032)
         );
  NAND4X0 U3981 ( .IN1(n4033), .IN2(n4034), .IN3(n4035), .IN4(n4036), .QN(
        n4004) );
  OA221X1 U3982 ( .IN1(n26725), .IN2(n27), .IN3(n26733), .IN4(n70), .IN5(n4037), .Q(n4036) );
  OA22X1 U3983 ( .IN1(n26741), .IN2(n113), .IN3(n26749), .IN4(n156), .Q(n4037)
         );
  OA221X1 U3984 ( .IN1(n26693), .IN2(n199), .IN3(n26701), .IN4(n242), .IN5(
        n4038), .Q(n4035) );
  OA22X1 U3985 ( .IN1(n26709), .IN2(n285), .IN3(n26717), .IN4(n328), .Q(n4038)
         );
  OA221X1 U3986 ( .IN1(n26661), .IN2(n371), .IN3(n26669), .IN4(n414), .IN5(
        n4039), .Q(n4034) );
  OA22X1 U3987 ( .IN1(n26677), .IN2(n457), .IN3(n26685), .IN4(n500), .Q(n4039)
         );
  OA221X1 U3988 ( .IN1(n26629), .IN2(n543), .IN3(n26637), .IN4(n586), .IN5(
        n4040), .Q(n4033) );
  OA22X1 U3989 ( .IN1(n26645), .IN2(n629), .IN3(n26653), .IN4(n672), .Q(n4040)
         );
  OR4X1 U3990 ( .IN1(n4041), .IN2(n4042), .IN3(n4043), .IN4(n4044), .Q(n2190)
         );
  AO221X1 U3991 ( .IN1(n2157), .IN2(n4045), .IN3(n2159), .IN4(n4046), .IN5(
        n4047), .Q(n4044) );
  AO22X1 U3992 ( .IN1(n2162), .IN2(n4048), .IN3(n2164), .IN4(n4049), .Q(n4047)
         );
  NAND4X0 U3993 ( .IN1(n4050), .IN2(n4051), .IN3(n4052), .IN4(n4053), .QN(
        n4049) );
  OA221X1 U3994 ( .IN1(n26596), .IN2(n27), .IN3(n26604), .IN4(n70), .IN5(n4054), .Q(n4053) );
  OA22X1 U3995 ( .IN1(n26612), .IN2(n113), .IN3(n26620), .IN4(n156), .Q(n4054)
         );
  OA221X1 U3996 ( .IN1(n26564), .IN2(n199), .IN3(n26572), .IN4(n242), .IN5(
        n4055), .Q(n4052) );
  OA22X1 U3997 ( .IN1(n26580), .IN2(n285), .IN3(n26588), .IN4(n328), .Q(n4055)
         );
  OA221X1 U3998 ( .IN1(n26532), .IN2(n371), .IN3(n26540), .IN4(n414), .IN5(
        n4056), .Q(n4051) );
  OA22X1 U3999 ( .IN1(n26548), .IN2(n457), .IN3(n26556), .IN4(n500), .Q(n4056)
         );
  OA221X1 U4000 ( .IN1(n26500), .IN2(n543), .IN3(n26508), .IN4(n586), .IN5(
        n4057), .Q(n4050) );
  OA22X1 U4001 ( .IN1(n26516), .IN2(n629), .IN3(n26524), .IN4(n672), .Q(n4057)
         );
  NAND4X0 U4002 ( .IN1(n4058), .IN2(n4059), .IN3(n4060), .IN4(n4061), .QN(
        n4048) );
  OA221X1 U4003 ( .IN1(n26468), .IN2(n27), .IN3(n26476), .IN4(n70), .IN5(n4062), .Q(n4061) );
  OA22X1 U4004 ( .IN1(n26484), .IN2(n113), .IN3(n26492), .IN4(n156), .Q(n4062)
         );
  OA221X1 U4005 ( .IN1(n26436), .IN2(n199), .IN3(n26444), .IN4(n242), .IN5(
        n4063), .Q(n4060) );
  OA22X1 U4006 ( .IN1(n26452), .IN2(n285), .IN3(n26460), .IN4(n328), .Q(n4063)
         );
  OA221X1 U4007 ( .IN1(n26404), .IN2(n371), .IN3(n26412), .IN4(n414), .IN5(
        n4064), .Q(n4059) );
  OA22X1 U4008 ( .IN1(n26420), .IN2(n457), .IN3(n26428), .IN4(n500), .Q(n4064)
         );
  OA221X1 U4009 ( .IN1(n26372), .IN2(n543), .IN3(n26380), .IN4(n586), .IN5(
        n4065), .Q(n4058) );
  OA22X1 U4010 ( .IN1(n26388), .IN2(n629), .IN3(n26396), .IN4(n672), .Q(n4065)
         );
  NAND4X0 U4011 ( .IN1(n4066), .IN2(n4067), .IN3(n4068), .IN4(n4069), .QN(
        n4046) );
  OA221X1 U4012 ( .IN1(n26340), .IN2(n27), .IN3(n26348), .IN4(n70), .IN5(n4070), .Q(n4069) );
  OA22X1 U4013 ( .IN1(n26356), .IN2(n113), .IN3(n26364), .IN4(n156), .Q(n4070)
         );
  OA221X1 U4014 ( .IN1(n26308), .IN2(n199), .IN3(n26316), .IN4(n242), .IN5(
        n4071), .Q(n4068) );
  OA22X1 U4015 ( .IN1(n26324), .IN2(n285), .IN3(n26332), .IN4(n328), .Q(n4071)
         );
  OA221X1 U4016 ( .IN1(n26276), .IN2(n371), .IN3(n26284), .IN4(n414), .IN5(
        n4072), .Q(n4067) );
  OA22X1 U4017 ( .IN1(n26292), .IN2(n457), .IN3(n26300), .IN4(n500), .Q(n4072)
         );
  OA221X1 U4018 ( .IN1(n26244), .IN2(n543), .IN3(n26252), .IN4(n586), .IN5(
        n4073), .Q(n4066) );
  OA22X1 U4019 ( .IN1(n26260), .IN2(n629), .IN3(n26268), .IN4(n672), .Q(n4073)
         );
  NAND4X0 U4020 ( .IN1(n4074), .IN2(n4075), .IN3(n4076), .IN4(n4077), .QN(
        n4045) );
  OA221X1 U4021 ( .IN1(n26212), .IN2(n27), .IN3(n26220), .IN4(n70), .IN5(n4078), .Q(n4077) );
  OA22X1 U4022 ( .IN1(n26228), .IN2(n113), .IN3(n26236), .IN4(n156), .Q(n4078)
         );
  OA221X1 U4023 ( .IN1(n26180), .IN2(n199), .IN3(n26188), .IN4(n242), .IN5(
        n4079), .Q(n4076) );
  OA22X1 U4024 ( .IN1(n26196), .IN2(n285), .IN3(n26204), .IN4(n328), .Q(n4079)
         );
  OA221X1 U4025 ( .IN1(n26148), .IN2(n371), .IN3(n26156), .IN4(n414), .IN5(
        n4080), .Q(n4075) );
  OA22X1 U4026 ( .IN1(n26164), .IN2(n457), .IN3(n26172), .IN4(n500), .Q(n4080)
         );
  OA221X1 U4027 ( .IN1(n26116), .IN2(n543), .IN3(n26124), .IN4(n586), .IN5(
        n4081), .Q(n4074) );
  OA22X1 U4028 ( .IN1(n26132), .IN2(n629), .IN3(n26140), .IN4(n672), .Q(n4081)
         );
  AO221X1 U4029 ( .IN1(n2246), .IN2(n4082), .IN3(n2248), .IN4(n4083), .IN5(
        n4084), .Q(n4043) );
  AO22X1 U4030 ( .IN1(n2251), .IN2(n4085), .IN3(n2253), .IN4(n4086), .Q(n4084)
         );
  NAND4X0 U4031 ( .IN1(n4087), .IN2(n4088), .IN3(n4089), .IN4(n4090), .QN(
        n4086) );
  OA221X1 U4032 ( .IN1(n26084), .IN2(n27), .IN3(n26092), .IN4(n70), .IN5(n4091), .Q(n4090) );
  OA22X1 U4033 ( .IN1(n26100), .IN2(n113), .IN3(n26108), .IN4(n156), .Q(n4091)
         );
  OA221X1 U4034 ( .IN1(n26052), .IN2(n199), .IN3(n26060), .IN4(n242), .IN5(
        n4092), .Q(n4089) );
  OA22X1 U4035 ( .IN1(n26068), .IN2(n285), .IN3(n26076), .IN4(n328), .Q(n4092)
         );
  OA221X1 U4036 ( .IN1(n26020), .IN2(n371), .IN3(n26028), .IN4(n414), .IN5(
        n4093), .Q(n4088) );
  OA22X1 U4037 ( .IN1(n26036), .IN2(n457), .IN3(n26044), .IN4(n500), .Q(n4093)
         );
  OA221X1 U4038 ( .IN1(n25988), .IN2(n543), .IN3(n25996), .IN4(n586), .IN5(
        n4094), .Q(n4087) );
  OA22X1 U4039 ( .IN1(n26004), .IN2(n629), .IN3(n26012), .IN4(n672), .Q(n4094)
         );
  NAND4X0 U4040 ( .IN1(n4095), .IN2(n4096), .IN3(n4097), .IN4(n4098), .QN(
        n4085) );
  OA221X1 U4041 ( .IN1(n25956), .IN2(n27), .IN3(n25964), .IN4(n70), .IN5(n4099), .Q(n4098) );
  OA22X1 U4042 ( .IN1(n25972), .IN2(n113), .IN3(n25980), .IN4(n156), .Q(n4099)
         );
  OA221X1 U4043 ( .IN1(n25924), .IN2(n199), .IN3(n25932), .IN4(n242), .IN5(
        n4100), .Q(n4097) );
  OA22X1 U4044 ( .IN1(n25940), .IN2(n285), .IN3(n25948), .IN4(n328), .Q(n4100)
         );
  OA221X1 U4045 ( .IN1(n25892), .IN2(n371), .IN3(n25900), .IN4(n414), .IN5(
        n4101), .Q(n4096) );
  OA22X1 U4046 ( .IN1(n25908), .IN2(n457), .IN3(n25916), .IN4(n500), .Q(n4101)
         );
  OA221X1 U4047 ( .IN1(n25860), .IN2(n543), .IN3(n25868), .IN4(n586), .IN5(
        n4102), .Q(n4095) );
  OA22X1 U4048 ( .IN1(n25876), .IN2(n629), .IN3(n25884), .IN4(n672), .Q(n4102)
         );
  NAND4X0 U4049 ( .IN1(n4103), .IN2(n4104), .IN3(n4105), .IN4(n4106), .QN(
        n4083) );
  OA221X1 U4050 ( .IN1(n25828), .IN2(n27), .IN3(n25836), .IN4(n70), .IN5(n4107), .Q(n4106) );
  OA22X1 U4051 ( .IN1(n25844), .IN2(n113), .IN3(n25852), .IN4(n156), .Q(n4107)
         );
  OA221X1 U4052 ( .IN1(n25796), .IN2(n199), .IN3(n25804), .IN4(n242), .IN5(
        n4108), .Q(n4105) );
  OA22X1 U4053 ( .IN1(n25812), .IN2(n285), .IN3(n25820), .IN4(n328), .Q(n4108)
         );
  OA221X1 U4054 ( .IN1(n25764), .IN2(n371), .IN3(n25772), .IN4(n414), .IN5(
        n4109), .Q(n4104) );
  OA22X1 U4055 ( .IN1(n25780), .IN2(n457), .IN3(n25788), .IN4(n500), .Q(n4109)
         );
  OA221X1 U4056 ( .IN1(n25732), .IN2(n543), .IN3(n25740), .IN4(n586), .IN5(
        n4110), .Q(n4103) );
  OA22X1 U4057 ( .IN1(n25748), .IN2(n629), .IN3(n25756), .IN4(n672), .Q(n4110)
         );
  NAND4X0 U4058 ( .IN1(n4111), .IN2(n4112), .IN3(n4113), .IN4(n4114), .QN(
        n4082) );
  OA221X1 U4059 ( .IN1(n25700), .IN2(n27), .IN3(n25708), .IN4(n70), .IN5(n4115), .Q(n4114) );
  OA22X1 U4060 ( .IN1(n25716), .IN2(n113), .IN3(n25724), .IN4(n156), .Q(n4115)
         );
  OA221X1 U4061 ( .IN1(n25668), .IN2(n199), .IN3(n25676), .IN4(n242), .IN5(
        n4116), .Q(n4113) );
  OA22X1 U4062 ( .IN1(n25684), .IN2(n285), .IN3(n25692), .IN4(n328), .Q(n4116)
         );
  OA221X1 U4063 ( .IN1(n25636), .IN2(n371), .IN3(n25644), .IN4(n414), .IN5(
        n4117), .Q(n4112) );
  OA22X1 U4064 ( .IN1(n25652), .IN2(n457), .IN3(n25660), .IN4(n500), .Q(n4117)
         );
  OA221X1 U4065 ( .IN1(n25604), .IN2(n543), .IN3(n25612), .IN4(n586), .IN5(
        n4118), .Q(n4111) );
  OA22X1 U4066 ( .IN1(n25620), .IN2(n629), .IN3(n25628), .IN4(n672), .Q(n4118)
         );
  AO221X1 U4067 ( .IN1(n2287), .IN2(n4119), .IN3(n2289), .IN4(n4120), .IN5(
        n4121), .Q(n4042) );
  AO22X1 U4068 ( .IN1(n2292), .IN2(n4122), .IN3(n2294), .IN4(n4123), .Q(n4121)
         );
  NAND4X0 U4069 ( .IN1(n4124), .IN2(n4125), .IN3(n4126), .IN4(n4127), .QN(
        n4123) );
  OA221X1 U4070 ( .IN1(n27620), .IN2(n26), .IN3(n27628), .IN4(n69), .IN5(n4128), .Q(n4127) );
  OA22X1 U4071 ( .IN1(n27636), .IN2(n112), .IN3(n27644), .IN4(n155), .Q(n4128)
         );
  OA221X1 U4072 ( .IN1(n27588), .IN2(n198), .IN3(n27596), .IN4(n241), .IN5(
        n4129), .Q(n4126) );
  OA22X1 U4073 ( .IN1(n27604), .IN2(n284), .IN3(n27612), .IN4(n327), .Q(n4129)
         );
  OA221X1 U4074 ( .IN1(n27556), .IN2(n370), .IN3(n27564), .IN4(n413), .IN5(
        n4130), .Q(n4125) );
  OA22X1 U4075 ( .IN1(n27572), .IN2(n456), .IN3(n27580), .IN4(n499), .Q(n4130)
         );
  OA221X1 U4076 ( .IN1(n27524), .IN2(n542), .IN3(n27532), .IN4(n585), .IN5(
        n4131), .Q(n4124) );
  OA22X1 U4077 ( .IN1(n27540), .IN2(n628), .IN3(n27548), .IN4(n671), .Q(n4131)
         );
  NAND4X0 U4078 ( .IN1(n4132), .IN2(n4133), .IN3(n4134), .IN4(n4135), .QN(
        n4122) );
  OA221X1 U4079 ( .IN1(n27492), .IN2(n26), .IN3(n27500), .IN4(n69), .IN5(n4136), .Q(n4135) );
  OA22X1 U4080 ( .IN1(n27508), .IN2(n112), .IN3(n27516), .IN4(n155), .Q(n4136)
         );
  OA221X1 U4081 ( .IN1(n27460), .IN2(n198), .IN3(n27468), .IN4(n241), .IN5(
        n4137), .Q(n4134) );
  OA22X1 U4082 ( .IN1(n27476), .IN2(n284), .IN3(n27484), .IN4(n327), .Q(n4137)
         );
  OA221X1 U4083 ( .IN1(n27428), .IN2(n370), .IN3(n27436), .IN4(n413), .IN5(
        n4138), .Q(n4133) );
  OA22X1 U4084 ( .IN1(n27444), .IN2(n456), .IN3(n27452), .IN4(n499), .Q(n4138)
         );
  OA221X1 U4085 ( .IN1(n27396), .IN2(n542), .IN3(n27404), .IN4(n585), .IN5(
        n4139), .Q(n4132) );
  OA22X1 U4086 ( .IN1(n27412), .IN2(n628), .IN3(n27420), .IN4(n671), .Q(n4139)
         );
  NAND4X0 U4087 ( .IN1(n4140), .IN2(n4141), .IN3(n4142), .IN4(n4143), .QN(
        n4120) );
  OA221X1 U4088 ( .IN1(n27364), .IN2(n26), .IN3(n27372), .IN4(n69), .IN5(n4144), .Q(n4143) );
  OA22X1 U4089 ( .IN1(n27380), .IN2(n112), .IN3(n27388), .IN4(n155), .Q(n4144)
         );
  OA221X1 U4090 ( .IN1(n27332), .IN2(n198), .IN3(n27340), .IN4(n241), .IN5(
        n4145), .Q(n4142) );
  OA22X1 U4091 ( .IN1(n27348), .IN2(n284), .IN3(n27356), .IN4(n327), .Q(n4145)
         );
  OA221X1 U4092 ( .IN1(n27300), .IN2(n370), .IN3(n27308), .IN4(n413), .IN5(
        n4146), .Q(n4141) );
  OA22X1 U4093 ( .IN1(n27316), .IN2(n456), .IN3(n27324), .IN4(n499), .Q(n4146)
         );
  OA221X1 U4094 ( .IN1(n27268), .IN2(n542), .IN3(n27276), .IN4(n585), .IN5(
        n4147), .Q(n4140) );
  OA22X1 U4095 ( .IN1(n27284), .IN2(n628), .IN3(n27292), .IN4(n671), .Q(n4147)
         );
  NAND4X0 U4096 ( .IN1(n4148), .IN2(n4149), .IN3(n4150), .IN4(n4151), .QN(
        n4119) );
  OA221X1 U4097 ( .IN1(n27236), .IN2(n26), .IN3(n27244), .IN4(n69), .IN5(n4152), .Q(n4151) );
  OA22X1 U4098 ( .IN1(n27252), .IN2(n112), .IN3(n27260), .IN4(n155), .Q(n4152)
         );
  OA221X1 U4099 ( .IN1(n27204), .IN2(n198), .IN3(n27212), .IN4(n241), .IN5(
        n4153), .Q(n4150) );
  OA22X1 U4100 ( .IN1(n27220), .IN2(n284), .IN3(n27228), .IN4(n327), .Q(n4153)
         );
  OA221X1 U4101 ( .IN1(n27172), .IN2(n370), .IN3(n27180), .IN4(n413), .IN5(
        n4154), .Q(n4149) );
  OA22X1 U4102 ( .IN1(n27188), .IN2(n456), .IN3(n27196), .IN4(n499), .Q(n4154)
         );
  OA221X1 U4103 ( .IN1(n27140), .IN2(n542), .IN3(n27148), .IN4(n585), .IN5(
        n4155), .Q(n4148) );
  OA22X1 U4104 ( .IN1(n27156), .IN2(n628), .IN3(n27164), .IN4(n671), .Q(n4155)
         );
  AO221X1 U4105 ( .IN1(n2328), .IN2(n4156), .IN3(n2330), .IN4(n4157), .IN5(
        n4158), .Q(n4041) );
  AO22X1 U4106 ( .IN1(n2333), .IN2(n4159), .IN3(n2335), .IN4(n4160), .Q(n4158)
         );
  NAND4X0 U4107 ( .IN1(n4161), .IN2(n4162), .IN3(n4163), .IN4(n4164), .QN(
        n4160) );
  OA221X1 U4108 ( .IN1(n27108), .IN2(n26), .IN3(n27116), .IN4(n69), .IN5(n4165), .Q(n4164) );
  OA22X1 U4109 ( .IN1(n27124), .IN2(n112), .IN3(n27132), .IN4(n155), .Q(n4165)
         );
  OA221X1 U4110 ( .IN1(n27076), .IN2(n198), .IN3(n27084), .IN4(n241), .IN5(
        n4166), .Q(n4163) );
  OA22X1 U4111 ( .IN1(n27092), .IN2(n284), .IN3(n27100), .IN4(n327), .Q(n4166)
         );
  OA221X1 U4112 ( .IN1(n27044), .IN2(n370), .IN3(n27052), .IN4(n413), .IN5(
        n4167), .Q(n4162) );
  OA22X1 U4113 ( .IN1(n27060), .IN2(n456), .IN3(n27068), .IN4(n499), .Q(n4167)
         );
  OA221X1 U4114 ( .IN1(n27012), .IN2(n542), .IN3(n27020), .IN4(n585), .IN5(
        n4168), .Q(n4161) );
  OA22X1 U4115 ( .IN1(n27028), .IN2(n628), .IN3(n27036), .IN4(n671), .Q(n4168)
         );
  NAND4X0 U4116 ( .IN1(n4169), .IN2(n4170), .IN3(n4171), .IN4(n4172), .QN(
        n4159) );
  OA221X1 U4117 ( .IN1(n26980), .IN2(n26), .IN3(n26988), .IN4(n69), .IN5(n4173), .Q(n4172) );
  OA22X1 U4118 ( .IN1(n26996), .IN2(n112), .IN3(n27004), .IN4(n155), .Q(n4173)
         );
  OA221X1 U4119 ( .IN1(n26948), .IN2(n198), .IN3(n26956), .IN4(n241), .IN5(
        n4174), .Q(n4171) );
  OA22X1 U4120 ( .IN1(n26964), .IN2(n284), .IN3(n26972), .IN4(n327), .Q(n4174)
         );
  OA221X1 U4121 ( .IN1(n26916), .IN2(n370), .IN3(n26924), .IN4(n413), .IN5(
        n4175), .Q(n4170) );
  OA22X1 U4122 ( .IN1(n26932), .IN2(n456), .IN3(n26940), .IN4(n499), .Q(n4175)
         );
  OA221X1 U4123 ( .IN1(n26884), .IN2(n542), .IN3(n26892), .IN4(n585), .IN5(
        n4176), .Q(n4169) );
  OA22X1 U4124 ( .IN1(n26900), .IN2(n628), .IN3(n26908), .IN4(n671), .Q(n4176)
         );
  NAND4X0 U4125 ( .IN1(n4177), .IN2(n4178), .IN3(n4179), .IN4(n4180), .QN(
        n4157) );
  OA221X1 U4126 ( .IN1(n26852), .IN2(n26), .IN3(n26860), .IN4(n69), .IN5(n4181), .Q(n4180) );
  OA22X1 U4127 ( .IN1(n26868), .IN2(n112), .IN3(n26876), .IN4(n155), .Q(n4181)
         );
  OA221X1 U4128 ( .IN1(n26820), .IN2(n198), .IN3(n26828), .IN4(n241), .IN5(
        n4182), .Q(n4179) );
  OA22X1 U4129 ( .IN1(n26836), .IN2(n284), .IN3(n26844), .IN4(n327), .Q(n4182)
         );
  OA221X1 U4130 ( .IN1(n26788), .IN2(n370), .IN3(n26796), .IN4(n413), .IN5(
        n4183), .Q(n4178) );
  OA22X1 U4131 ( .IN1(n26804), .IN2(n456), .IN3(n26812), .IN4(n499), .Q(n4183)
         );
  OA221X1 U4132 ( .IN1(n26756), .IN2(n542), .IN3(n26764), .IN4(n585), .IN5(
        n4184), .Q(n4177) );
  OA22X1 U4133 ( .IN1(n26772), .IN2(n628), .IN3(n26780), .IN4(n671), .Q(n4184)
         );
  NAND4X0 U4134 ( .IN1(n4185), .IN2(n4186), .IN3(n4187), .IN4(n4188), .QN(
        n4156) );
  OA221X1 U4135 ( .IN1(n26724), .IN2(n26), .IN3(n26732), .IN4(n69), .IN5(n4189), .Q(n4188) );
  OA22X1 U4136 ( .IN1(n26740), .IN2(n112), .IN3(n26748), .IN4(n155), .Q(n4189)
         );
  OA221X1 U4137 ( .IN1(n26692), .IN2(n198), .IN3(n26700), .IN4(n241), .IN5(
        n4190), .Q(n4187) );
  OA22X1 U4138 ( .IN1(n26708), .IN2(n284), .IN3(n26716), .IN4(n327), .Q(n4190)
         );
  OA221X1 U4139 ( .IN1(n26660), .IN2(n370), .IN3(n26668), .IN4(n413), .IN5(
        n4191), .Q(n4186) );
  OA22X1 U4140 ( .IN1(n26676), .IN2(n456), .IN3(n26684), .IN4(n499), .Q(n4191)
         );
  OA221X1 U4141 ( .IN1(n26628), .IN2(n542), .IN3(n26636), .IN4(n585), .IN5(
        n4192), .Q(n4185) );
  OA22X1 U4142 ( .IN1(n26644), .IN2(n628), .IN3(n26652), .IN4(n671), .Q(n4192)
         );
  OR4X1 U4143 ( .IN1(n4193), .IN2(n4194), .IN3(n4195), .IN4(n4196), .Q(n2189)
         );
  AO221X1 U4144 ( .IN1(n2157), .IN2(n4197), .IN3(n2159), .IN4(n4198), .IN5(
        n4199), .Q(n4196) );
  AO22X1 U4145 ( .IN1(n2162), .IN2(n4200), .IN3(n2164), .IN4(n4201), .Q(n4199)
         );
  NAND4X0 U4146 ( .IN1(n4202), .IN2(n4203), .IN3(n4204), .IN4(n4205), .QN(
        n4201) );
  OA221X1 U4147 ( .IN1(n26595), .IN2(n26), .IN3(n26603), .IN4(n69), .IN5(n4206), .Q(n4205) );
  OA22X1 U4148 ( .IN1(n26611), .IN2(n112), .IN3(n26619), .IN4(n155), .Q(n4206)
         );
  OA221X1 U4149 ( .IN1(n26563), .IN2(n198), .IN3(n26571), .IN4(n241), .IN5(
        n4207), .Q(n4204) );
  OA22X1 U4150 ( .IN1(n26579), .IN2(n284), .IN3(n26587), .IN4(n327), .Q(n4207)
         );
  OA221X1 U4151 ( .IN1(n26531), .IN2(n370), .IN3(n26539), .IN4(n413), .IN5(
        n4208), .Q(n4203) );
  OA22X1 U4152 ( .IN1(n26547), .IN2(n456), .IN3(n26555), .IN4(n499), .Q(n4208)
         );
  OA221X1 U4153 ( .IN1(n26499), .IN2(n542), .IN3(n26507), .IN4(n585), .IN5(
        n4209), .Q(n4202) );
  OA22X1 U4154 ( .IN1(n26515), .IN2(n628), .IN3(n26523), .IN4(n671), .Q(n4209)
         );
  NAND4X0 U4155 ( .IN1(n4210), .IN2(n4211), .IN3(n4212), .IN4(n4213), .QN(
        n4200) );
  OA221X1 U4156 ( .IN1(n26467), .IN2(n26), .IN3(n26475), .IN4(n69), .IN5(n4214), .Q(n4213) );
  OA22X1 U4157 ( .IN1(n26483), .IN2(n112), .IN3(n26491), .IN4(n155), .Q(n4214)
         );
  OA221X1 U4158 ( .IN1(n26435), .IN2(n198), .IN3(n26443), .IN4(n241), .IN5(
        n4215), .Q(n4212) );
  OA22X1 U4159 ( .IN1(n26451), .IN2(n284), .IN3(n26459), .IN4(n327), .Q(n4215)
         );
  OA221X1 U4160 ( .IN1(n26403), .IN2(n370), .IN3(n26411), .IN4(n413), .IN5(
        n4216), .Q(n4211) );
  OA22X1 U4161 ( .IN1(n26419), .IN2(n456), .IN3(n26427), .IN4(n499), .Q(n4216)
         );
  OA221X1 U4162 ( .IN1(n26371), .IN2(n542), .IN3(n26379), .IN4(n585), .IN5(
        n4217), .Q(n4210) );
  OA22X1 U4163 ( .IN1(n26387), .IN2(n628), .IN3(n26395), .IN4(n671), .Q(n4217)
         );
  NAND4X0 U4164 ( .IN1(n4218), .IN2(n4219), .IN3(n4220), .IN4(n4221), .QN(
        n4198) );
  OA221X1 U4165 ( .IN1(n26339), .IN2(n26), .IN3(n26347), .IN4(n69), .IN5(n4222), .Q(n4221) );
  OA22X1 U4166 ( .IN1(n26355), .IN2(n112), .IN3(n26363), .IN4(n155), .Q(n4222)
         );
  OA221X1 U4167 ( .IN1(n26307), .IN2(n198), .IN3(n26315), .IN4(n241), .IN5(
        n4223), .Q(n4220) );
  OA22X1 U4168 ( .IN1(n26323), .IN2(n284), .IN3(n26331), .IN4(n327), .Q(n4223)
         );
  OA221X1 U4169 ( .IN1(n26275), .IN2(n370), .IN3(n26283), .IN4(n413), .IN5(
        n4224), .Q(n4219) );
  OA22X1 U4170 ( .IN1(n26291), .IN2(n456), .IN3(n26299), .IN4(n499), .Q(n4224)
         );
  OA221X1 U4171 ( .IN1(n26243), .IN2(n542), .IN3(n26251), .IN4(n585), .IN5(
        n4225), .Q(n4218) );
  OA22X1 U4172 ( .IN1(n26259), .IN2(n628), .IN3(n26267), .IN4(n671), .Q(n4225)
         );
  NAND4X0 U4173 ( .IN1(n4226), .IN2(n4227), .IN3(n4228), .IN4(n4229), .QN(
        n4197) );
  OA221X1 U4174 ( .IN1(n26211), .IN2(n26), .IN3(n26219), .IN4(n69), .IN5(n4230), .Q(n4229) );
  OA22X1 U4175 ( .IN1(n26227), .IN2(n112), .IN3(n26235), .IN4(n155), .Q(n4230)
         );
  OA221X1 U4176 ( .IN1(n26179), .IN2(n198), .IN3(n26187), .IN4(n241), .IN5(
        n4231), .Q(n4228) );
  OA22X1 U4177 ( .IN1(n26195), .IN2(n284), .IN3(n26203), .IN4(n327), .Q(n4231)
         );
  OA221X1 U4178 ( .IN1(n26147), .IN2(n370), .IN3(n26155), .IN4(n413), .IN5(
        n4232), .Q(n4227) );
  OA22X1 U4179 ( .IN1(n26163), .IN2(n456), .IN3(n26171), .IN4(n499), .Q(n4232)
         );
  OA221X1 U4180 ( .IN1(n26115), .IN2(n542), .IN3(n26123), .IN4(n585), .IN5(
        n4233), .Q(n4226) );
  OA22X1 U4181 ( .IN1(n26131), .IN2(n628), .IN3(n26139), .IN4(n671), .Q(n4233)
         );
  AO221X1 U4182 ( .IN1(n2246), .IN2(n4234), .IN3(n2248), .IN4(n4235), .IN5(
        n4236), .Q(n4195) );
  AO22X1 U4183 ( .IN1(n2251), .IN2(n4237), .IN3(n2253), .IN4(n4238), .Q(n4236)
         );
  NAND4X0 U4184 ( .IN1(n4239), .IN2(n4240), .IN3(n4241), .IN4(n4242), .QN(
        n4238) );
  OA221X1 U4185 ( .IN1(n26083), .IN2(n25), .IN3(n26091), .IN4(n68), .IN5(n4243), .Q(n4242) );
  OA22X1 U4186 ( .IN1(n26099), .IN2(n111), .IN3(n26107), .IN4(n154), .Q(n4243)
         );
  OA221X1 U4187 ( .IN1(n26051), .IN2(n197), .IN3(n26059), .IN4(n240), .IN5(
        n4244), .Q(n4241) );
  OA22X1 U4188 ( .IN1(n26067), .IN2(n283), .IN3(n26075), .IN4(n326), .Q(n4244)
         );
  OA221X1 U4189 ( .IN1(n26019), .IN2(n369), .IN3(n26027), .IN4(n412), .IN5(
        n4245), .Q(n4240) );
  OA22X1 U4190 ( .IN1(n26035), .IN2(n455), .IN3(n26043), .IN4(n498), .Q(n4245)
         );
  OA221X1 U4191 ( .IN1(n25987), .IN2(n541), .IN3(n25995), .IN4(n584), .IN5(
        n4246), .Q(n4239) );
  OA22X1 U4192 ( .IN1(n26003), .IN2(n627), .IN3(n26011), .IN4(n670), .Q(n4246)
         );
  NAND4X0 U4193 ( .IN1(n4247), .IN2(n4248), .IN3(n4249), .IN4(n4250), .QN(
        n4237) );
  OA221X1 U4194 ( .IN1(n25955), .IN2(n25), .IN3(n25963), .IN4(n68), .IN5(n4251), .Q(n4250) );
  OA22X1 U4195 ( .IN1(n25971), .IN2(n111), .IN3(n25979), .IN4(n154), .Q(n4251)
         );
  OA221X1 U4196 ( .IN1(n25923), .IN2(n197), .IN3(n25931), .IN4(n240), .IN5(
        n4252), .Q(n4249) );
  OA22X1 U4197 ( .IN1(n25939), .IN2(n283), .IN3(n25947), .IN4(n326), .Q(n4252)
         );
  OA221X1 U4198 ( .IN1(n25891), .IN2(n369), .IN3(n25899), .IN4(n412), .IN5(
        n4253), .Q(n4248) );
  OA22X1 U4199 ( .IN1(n25907), .IN2(n455), .IN3(n25915), .IN4(n498), .Q(n4253)
         );
  OA221X1 U4200 ( .IN1(n25859), .IN2(n541), .IN3(n25867), .IN4(n584), .IN5(
        n4254), .Q(n4247) );
  OA22X1 U4201 ( .IN1(n25875), .IN2(n627), .IN3(n25883), .IN4(n670), .Q(n4254)
         );
  NAND4X0 U4202 ( .IN1(n4255), .IN2(n4256), .IN3(n4257), .IN4(n4258), .QN(
        n4235) );
  OA221X1 U4203 ( .IN1(n25827), .IN2(n25), .IN3(n25835), .IN4(n68), .IN5(n4259), .Q(n4258) );
  OA22X1 U4204 ( .IN1(n25843), .IN2(n111), .IN3(n25851), .IN4(n154), .Q(n4259)
         );
  OA221X1 U4205 ( .IN1(n25795), .IN2(n197), .IN3(n25803), .IN4(n240), .IN5(
        n4260), .Q(n4257) );
  OA22X1 U4206 ( .IN1(n25811), .IN2(n283), .IN3(n25819), .IN4(n326), .Q(n4260)
         );
  OA221X1 U4207 ( .IN1(n25763), .IN2(n369), .IN3(n25771), .IN4(n412), .IN5(
        n4261), .Q(n4256) );
  OA22X1 U4208 ( .IN1(n25779), .IN2(n455), .IN3(n25787), .IN4(n498), .Q(n4261)
         );
  OA221X1 U4209 ( .IN1(n25731), .IN2(n541), .IN3(n25739), .IN4(n584), .IN5(
        n4262), .Q(n4255) );
  OA22X1 U4210 ( .IN1(n25747), .IN2(n627), .IN3(n25755), .IN4(n670), .Q(n4262)
         );
  NAND4X0 U4211 ( .IN1(n4263), .IN2(n4264), .IN3(n4265), .IN4(n4266), .QN(
        n4234) );
  OA221X1 U4212 ( .IN1(n25699), .IN2(n25), .IN3(n25707), .IN4(n68), .IN5(n4267), .Q(n4266) );
  OA22X1 U4213 ( .IN1(n25715), .IN2(n111), .IN3(n25723), .IN4(n154), .Q(n4267)
         );
  OA221X1 U4214 ( .IN1(n25667), .IN2(n197), .IN3(n25675), .IN4(n240), .IN5(
        n4268), .Q(n4265) );
  OA22X1 U4215 ( .IN1(n25683), .IN2(n283), .IN3(n25691), .IN4(n326), .Q(n4268)
         );
  OA221X1 U4216 ( .IN1(n25635), .IN2(n369), .IN3(n25643), .IN4(n412), .IN5(
        n4269), .Q(n4264) );
  OA22X1 U4217 ( .IN1(n25651), .IN2(n455), .IN3(n25659), .IN4(n498), .Q(n4269)
         );
  OA221X1 U4218 ( .IN1(n25603), .IN2(n541), .IN3(n25611), .IN4(n584), .IN5(
        n4270), .Q(n4263) );
  OA22X1 U4219 ( .IN1(n25619), .IN2(n627), .IN3(n25627), .IN4(n670), .Q(n4270)
         );
  AO221X1 U4220 ( .IN1(n2287), .IN2(n4271), .IN3(n2289), .IN4(n4272), .IN5(
        n4273), .Q(n4194) );
  AO22X1 U4221 ( .IN1(n2292), .IN2(n4274), .IN3(n2294), .IN4(n4275), .Q(n4273)
         );
  NAND4X0 U4222 ( .IN1(n4276), .IN2(n4277), .IN3(n4278), .IN4(n4279), .QN(
        n4275) );
  OA221X1 U4223 ( .IN1(n27619), .IN2(n25), .IN3(n27627), .IN4(n68), .IN5(n4280), .Q(n4279) );
  OA22X1 U4224 ( .IN1(n27635), .IN2(n111), .IN3(n27643), .IN4(n154), .Q(n4280)
         );
  OA221X1 U4225 ( .IN1(n27587), .IN2(n197), .IN3(n27595), .IN4(n240), .IN5(
        n4281), .Q(n4278) );
  OA22X1 U4226 ( .IN1(n27603), .IN2(n283), .IN3(n27611), .IN4(n326), .Q(n4281)
         );
  OA221X1 U4227 ( .IN1(n27555), .IN2(n369), .IN3(n27563), .IN4(n412), .IN5(
        n4282), .Q(n4277) );
  OA22X1 U4228 ( .IN1(n27571), .IN2(n455), .IN3(n27579), .IN4(n498), .Q(n4282)
         );
  OA221X1 U4229 ( .IN1(n27523), .IN2(n541), .IN3(n27531), .IN4(n584), .IN5(
        n4283), .Q(n4276) );
  OA22X1 U4230 ( .IN1(n27539), .IN2(n627), .IN3(n27547), .IN4(n670), .Q(n4283)
         );
  NAND4X0 U4231 ( .IN1(n4284), .IN2(n4285), .IN3(n4286), .IN4(n4287), .QN(
        n4274) );
  OA221X1 U4232 ( .IN1(n27491), .IN2(n25), .IN3(n27499), .IN4(n68), .IN5(n4288), .Q(n4287) );
  OA22X1 U4233 ( .IN1(n27507), .IN2(n111), .IN3(n27515), .IN4(n154), .Q(n4288)
         );
  OA221X1 U4234 ( .IN1(n27459), .IN2(n197), .IN3(n27467), .IN4(n240), .IN5(
        n4289), .Q(n4286) );
  OA22X1 U4235 ( .IN1(n27475), .IN2(n283), .IN3(n27483), .IN4(n326), .Q(n4289)
         );
  OA221X1 U4236 ( .IN1(n27427), .IN2(n369), .IN3(n27435), .IN4(n412), .IN5(
        n4290), .Q(n4285) );
  OA22X1 U4237 ( .IN1(n27443), .IN2(n455), .IN3(n27451), .IN4(n498), .Q(n4290)
         );
  OA221X1 U4238 ( .IN1(n27395), .IN2(n541), .IN3(n27403), .IN4(n584), .IN5(
        n4291), .Q(n4284) );
  OA22X1 U4239 ( .IN1(n27411), .IN2(n627), .IN3(n27419), .IN4(n670), .Q(n4291)
         );
  NAND4X0 U4240 ( .IN1(n4292), .IN2(n4293), .IN3(n4294), .IN4(n4295), .QN(
        n4272) );
  OA221X1 U4241 ( .IN1(n27363), .IN2(n25), .IN3(n27371), .IN4(n68), .IN5(n4296), .Q(n4295) );
  OA22X1 U4242 ( .IN1(n27379), .IN2(n111), .IN3(n27387), .IN4(n154), .Q(n4296)
         );
  OA221X1 U4243 ( .IN1(n27331), .IN2(n197), .IN3(n27339), .IN4(n240), .IN5(
        n4297), .Q(n4294) );
  OA22X1 U4244 ( .IN1(n27347), .IN2(n283), .IN3(n27355), .IN4(n326), .Q(n4297)
         );
  OA221X1 U4245 ( .IN1(n27299), .IN2(n369), .IN3(n27307), .IN4(n412), .IN5(
        n4298), .Q(n4293) );
  OA22X1 U4246 ( .IN1(n27315), .IN2(n455), .IN3(n27323), .IN4(n498), .Q(n4298)
         );
  OA221X1 U4247 ( .IN1(n27267), .IN2(n541), .IN3(n27275), .IN4(n584), .IN5(
        n4299), .Q(n4292) );
  OA22X1 U4248 ( .IN1(n27283), .IN2(n627), .IN3(n27291), .IN4(n670), .Q(n4299)
         );
  NAND4X0 U4249 ( .IN1(n4300), .IN2(n4301), .IN3(n4302), .IN4(n4303), .QN(
        n4271) );
  OA221X1 U4250 ( .IN1(n27235), .IN2(n25), .IN3(n27243), .IN4(n68), .IN5(n4304), .Q(n4303) );
  OA22X1 U4251 ( .IN1(n27251), .IN2(n111), .IN3(n27259), .IN4(n154), .Q(n4304)
         );
  OA221X1 U4252 ( .IN1(n27203), .IN2(n197), .IN3(n27211), .IN4(n240), .IN5(
        n4305), .Q(n4302) );
  OA22X1 U4253 ( .IN1(n27219), .IN2(n283), .IN3(n27227), .IN4(n326), .Q(n4305)
         );
  OA221X1 U4254 ( .IN1(n27171), .IN2(n369), .IN3(n27179), .IN4(n412), .IN5(
        n4306), .Q(n4301) );
  OA22X1 U4255 ( .IN1(n27187), .IN2(n455), .IN3(n27195), .IN4(n498), .Q(n4306)
         );
  OA221X1 U4256 ( .IN1(n27139), .IN2(n541), .IN3(n27147), .IN4(n584), .IN5(
        n4307), .Q(n4300) );
  OA22X1 U4257 ( .IN1(n27155), .IN2(n627), .IN3(n27163), .IN4(n670), .Q(n4307)
         );
  AO221X1 U4258 ( .IN1(n2328), .IN2(n4308), .IN3(n2330), .IN4(n4309), .IN5(
        n4310), .Q(n4193) );
  AO22X1 U4259 ( .IN1(n2333), .IN2(n4311), .IN3(n2335), .IN4(n4312), .Q(n4310)
         );
  NAND4X0 U4260 ( .IN1(n4313), .IN2(n4314), .IN3(n4315), .IN4(n4316), .QN(
        n4312) );
  OA221X1 U4261 ( .IN1(n27107), .IN2(n25), .IN3(n27115), .IN4(n68), .IN5(n4317), .Q(n4316) );
  OA22X1 U4262 ( .IN1(n27123), .IN2(n111), .IN3(n27131), .IN4(n154), .Q(n4317)
         );
  OA221X1 U4263 ( .IN1(n27075), .IN2(n197), .IN3(n27083), .IN4(n240), .IN5(
        n4318), .Q(n4315) );
  OA22X1 U4264 ( .IN1(n27091), .IN2(n283), .IN3(n27099), .IN4(n326), .Q(n4318)
         );
  OA221X1 U4265 ( .IN1(n27043), .IN2(n369), .IN3(n27051), .IN4(n412), .IN5(
        n4319), .Q(n4314) );
  OA22X1 U4266 ( .IN1(n27059), .IN2(n455), .IN3(n27067), .IN4(n498), .Q(n4319)
         );
  OA221X1 U4267 ( .IN1(n27011), .IN2(n541), .IN3(n27019), .IN4(n584), .IN5(
        n4320), .Q(n4313) );
  OA22X1 U4268 ( .IN1(n27027), .IN2(n627), .IN3(n27035), .IN4(n670), .Q(n4320)
         );
  NAND4X0 U4269 ( .IN1(n4321), .IN2(n4322), .IN3(n4323), .IN4(n4324), .QN(
        n4311) );
  OA221X1 U4270 ( .IN1(n26979), .IN2(n25), .IN3(n26987), .IN4(n68), .IN5(n4325), .Q(n4324) );
  OA22X1 U4271 ( .IN1(n26995), .IN2(n111), .IN3(n27003), .IN4(n154), .Q(n4325)
         );
  OA221X1 U4272 ( .IN1(n26947), .IN2(n197), .IN3(n26955), .IN4(n240), .IN5(
        n4326), .Q(n4323) );
  OA22X1 U4273 ( .IN1(n26963), .IN2(n283), .IN3(n26971), .IN4(n326), .Q(n4326)
         );
  OA221X1 U4274 ( .IN1(n26915), .IN2(n369), .IN3(n26923), .IN4(n412), .IN5(
        n4327), .Q(n4322) );
  OA22X1 U4275 ( .IN1(n26931), .IN2(n455), .IN3(n26939), .IN4(n498), .Q(n4327)
         );
  OA221X1 U4276 ( .IN1(n26883), .IN2(n541), .IN3(n26891), .IN4(n584), .IN5(
        n4328), .Q(n4321) );
  OA22X1 U4277 ( .IN1(n26899), .IN2(n627), .IN3(n26907), .IN4(n670), .Q(n4328)
         );
  NAND4X0 U4278 ( .IN1(n4329), .IN2(n4330), .IN3(n4331), .IN4(n4332), .QN(
        n4309) );
  OA221X1 U4279 ( .IN1(n26851), .IN2(n25), .IN3(n26859), .IN4(n68), .IN5(n4333), .Q(n4332) );
  OA22X1 U4280 ( .IN1(n26867), .IN2(n111), .IN3(n26875), .IN4(n154), .Q(n4333)
         );
  OA221X1 U4281 ( .IN1(n26819), .IN2(n197), .IN3(n26827), .IN4(n240), .IN5(
        n4334), .Q(n4331) );
  OA22X1 U4282 ( .IN1(n26835), .IN2(n283), .IN3(n26843), .IN4(n326), .Q(n4334)
         );
  OA221X1 U4283 ( .IN1(n26787), .IN2(n369), .IN3(n26795), .IN4(n412), .IN5(
        n4335), .Q(n4330) );
  OA22X1 U4284 ( .IN1(n26803), .IN2(n455), .IN3(n26811), .IN4(n498), .Q(n4335)
         );
  OA221X1 U4285 ( .IN1(n26755), .IN2(n541), .IN3(n26763), .IN4(n584), .IN5(
        n4336), .Q(n4329) );
  OA22X1 U4286 ( .IN1(n26771), .IN2(n627), .IN3(n26779), .IN4(n670), .Q(n4336)
         );
  NAND4X0 U4287 ( .IN1(n4337), .IN2(n4338), .IN3(n4339), .IN4(n4340), .QN(
        n4308) );
  OA221X1 U4288 ( .IN1(n26723), .IN2(n25), .IN3(n26731), .IN4(n68), .IN5(n4341), .Q(n4340) );
  OA22X1 U4289 ( .IN1(n26739), .IN2(n111), .IN3(n26747), .IN4(n154), .Q(n4341)
         );
  OA221X1 U4290 ( .IN1(n26691), .IN2(n197), .IN3(n26699), .IN4(n240), .IN5(
        n4342), .Q(n4339) );
  OA22X1 U4291 ( .IN1(n26707), .IN2(n283), .IN3(n26715), .IN4(n326), .Q(n4342)
         );
  OA221X1 U4292 ( .IN1(n26659), .IN2(n369), .IN3(n26667), .IN4(n412), .IN5(
        n4343), .Q(n4338) );
  OA22X1 U4293 ( .IN1(n26675), .IN2(n455), .IN3(n26683), .IN4(n498), .Q(n4343)
         );
  OA221X1 U4294 ( .IN1(n26627), .IN2(n541), .IN3(n26635), .IN4(n584), .IN5(
        n4344), .Q(n4337) );
  OA22X1 U4295 ( .IN1(n26643), .IN2(n627), .IN3(n26651), .IN4(n670), .Q(n4344)
         );
  OR4X1 U4296 ( .IN1(n4345), .IN2(n4346), .IN3(n4347), .IN4(n4348), .Q(n2188)
         );
  AO221X1 U4297 ( .IN1(n2157), .IN2(n4349), .IN3(n2159), .IN4(n4350), .IN5(
        n4351), .Q(n4348) );
  AO22X1 U4298 ( .IN1(n2162), .IN2(n4352), .IN3(n2164), .IN4(n4353), .Q(n4351)
         );
  NAND4X0 U4299 ( .IN1(n4354), .IN2(n4355), .IN3(n4356), .IN4(n4357), .QN(
        n4353) );
  OA221X1 U4300 ( .IN1(n26594), .IN2(n24), .IN3(n26602), .IN4(n67), .IN5(n4358), .Q(n4357) );
  OA22X1 U4301 ( .IN1(n26610), .IN2(n110), .IN3(n26618), .IN4(n153), .Q(n4358)
         );
  OA221X1 U4302 ( .IN1(n26562), .IN2(n196), .IN3(n26570), .IN4(n239), .IN5(
        n4359), .Q(n4356) );
  OA22X1 U4303 ( .IN1(n26578), .IN2(n282), .IN3(n26586), .IN4(n325), .Q(n4359)
         );
  OA221X1 U4304 ( .IN1(n26530), .IN2(n368), .IN3(n26538), .IN4(n411), .IN5(
        n4360), .Q(n4355) );
  OA22X1 U4305 ( .IN1(n26546), .IN2(n454), .IN3(n26554), .IN4(n497), .Q(n4360)
         );
  OA221X1 U4306 ( .IN1(n26498), .IN2(n540), .IN3(n26506), .IN4(n583), .IN5(
        n4361), .Q(n4354) );
  OA22X1 U4307 ( .IN1(n26514), .IN2(n626), .IN3(n26522), .IN4(n669), .Q(n4361)
         );
  NAND4X0 U4308 ( .IN1(n4362), .IN2(n4363), .IN3(n4364), .IN4(n4365), .QN(
        n4352) );
  OA221X1 U4309 ( .IN1(n26466), .IN2(n24), .IN3(n26474), .IN4(n67), .IN5(n4366), .Q(n4365) );
  OA22X1 U4310 ( .IN1(n26482), .IN2(n110), .IN3(n26490), .IN4(n153), .Q(n4366)
         );
  OA221X1 U4311 ( .IN1(n26434), .IN2(n196), .IN3(n26442), .IN4(n239), .IN5(
        n4367), .Q(n4364) );
  OA22X1 U4312 ( .IN1(n26450), .IN2(n282), .IN3(n26458), .IN4(n325), .Q(n4367)
         );
  OA221X1 U4313 ( .IN1(n26402), .IN2(n368), .IN3(n26410), .IN4(n411), .IN5(
        n4368), .Q(n4363) );
  OA22X1 U4314 ( .IN1(n26418), .IN2(n454), .IN3(n26426), .IN4(n497), .Q(n4368)
         );
  OA221X1 U4315 ( .IN1(n26370), .IN2(n540), .IN3(n26378), .IN4(n583), .IN5(
        n4369), .Q(n4362) );
  OA22X1 U4316 ( .IN1(n26386), .IN2(n626), .IN3(n26394), .IN4(n669), .Q(n4369)
         );
  NAND4X0 U4317 ( .IN1(n4370), .IN2(n4371), .IN3(n4372), .IN4(n4373), .QN(
        n4350) );
  OA221X1 U4318 ( .IN1(n26338), .IN2(n24), .IN3(n26346), .IN4(n67), .IN5(n4374), .Q(n4373) );
  OA22X1 U4319 ( .IN1(n26354), .IN2(n110), .IN3(n26362), .IN4(n153), .Q(n4374)
         );
  OA221X1 U4320 ( .IN1(n26306), .IN2(n196), .IN3(n26314), .IN4(n239), .IN5(
        n4375), .Q(n4372) );
  OA22X1 U4321 ( .IN1(n26322), .IN2(n282), .IN3(n26330), .IN4(n325), .Q(n4375)
         );
  OA221X1 U4322 ( .IN1(n26274), .IN2(n368), .IN3(n26282), .IN4(n411), .IN5(
        n4376), .Q(n4371) );
  OA22X1 U4323 ( .IN1(n26290), .IN2(n454), .IN3(n26298), .IN4(n497), .Q(n4376)
         );
  OA221X1 U4324 ( .IN1(n26242), .IN2(n540), .IN3(n26250), .IN4(n583), .IN5(
        n4377), .Q(n4370) );
  OA22X1 U4325 ( .IN1(n26258), .IN2(n626), .IN3(n26266), .IN4(n669), .Q(n4377)
         );
  NAND4X0 U4326 ( .IN1(n4378), .IN2(n4379), .IN3(n4380), .IN4(n4381), .QN(
        n4349) );
  OA221X1 U4327 ( .IN1(n26210), .IN2(n24), .IN3(n26218), .IN4(n67), .IN5(n4382), .Q(n4381) );
  OA22X1 U4328 ( .IN1(n26226), .IN2(n110), .IN3(n26234), .IN4(n153), .Q(n4382)
         );
  OA221X1 U4329 ( .IN1(n26178), .IN2(n196), .IN3(n26186), .IN4(n239), .IN5(
        n4383), .Q(n4380) );
  OA22X1 U4330 ( .IN1(n26194), .IN2(n282), .IN3(n26202), .IN4(n325), .Q(n4383)
         );
  OA221X1 U4331 ( .IN1(n26146), .IN2(n368), .IN3(n26154), .IN4(n411), .IN5(
        n4384), .Q(n4379) );
  OA22X1 U4332 ( .IN1(n26162), .IN2(n454), .IN3(n26170), .IN4(n497), .Q(n4384)
         );
  OA221X1 U4333 ( .IN1(n26114), .IN2(n540), .IN3(n26122), .IN4(n583), .IN5(
        n4385), .Q(n4378) );
  OA22X1 U4334 ( .IN1(n26130), .IN2(n626), .IN3(n26138), .IN4(n669), .Q(n4385)
         );
  AO221X1 U4335 ( .IN1(n2246), .IN2(n4386), .IN3(n2248), .IN4(n4387), .IN5(
        n4388), .Q(n4347) );
  AO22X1 U4336 ( .IN1(n2251), .IN2(n4389), .IN3(n2253), .IN4(n4390), .Q(n4388)
         );
  NAND4X0 U4337 ( .IN1(n4391), .IN2(n4392), .IN3(n4393), .IN4(n4394), .QN(
        n4390) );
  OA221X1 U4338 ( .IN1(n26082), .IN2(n24), .IN3(n26090), .IN4(n67), .IN5(n4395), .Q(n4394) );
  OA22X1 U4339 ( .IN1(n26098), .IN2(n110), .IN3(n26106), .IN4(n153), .Q(n4395)
         );
  OA221X1 U4340 ( .IN1(n26050), .IN2(n196), .IN3(n26058), .IN4(n239), .IN5(
        n4396), .Q(n4393) );
  OA22X1 U4341 ( .IN1(n26066), .IN2(n282), .IN3(n26074), .IN4(n325), .Q(n4396)
         );
  OA221X1 U4342 ( .IN1(n26018), .IN2(n368), .IN3(n26026), .IN4(n411), .IN5(
        n4397), .Q(n4392) );
  OA22X1 U4343 ( .IN1(n26034), .IN2(n454), .IN3(n26042), .IN4(n497), .Q(n4397)
         );
  OA221X1 U4344 ( .IN1(n25986), .IN2(n540), .IN3(n25994), .IN4(n583), .IN5(
        n4398), .Q(n4391) );
  OA22X1 U4345 ( .IN1(n26002), .IN2(n626), .IN3(n26010), .IN4(n669), .Q(n4398)
         );
  NAND4X0 U4346 ( .IN1(n4399), .IN2(n4400), .IN3(n4401), .IN4(n4402), .QN(
        n4389) );
  OA221X1 U4347 ( .IN1(n25954), .IN2(n24), .IN3(n25962), .IN4(n67), .IN5(n4403), .Q(n4402) );
  OA22X1 U4348 ( .IN1(n25970), .IN2(n110), .IN3(n25978), .IN4(n153), .Q(n4403)
         );
  OA221X1 U4349 ( .IN1(n25922), .IN2(n196), .IN3(n25930), .IN4(n239), .IN5(
        n4404), .Q(n4401) );
  OA22X1 U4350 ( .IN1(n25938), .IN2(n282), .IN3(n25946), .IN4(n325), .Q(n4404)
         );
  OA221X1 U4351 ( .IN1(n25890), .IN2(n368), .IN3(n25898), .IN4(n411), .IN5(
        n4405), .Q(n4400) );
  OA22X1 U4352 ( .IN1(n25906), .IN2(n454), .IN3(n25914), .IN4(n497), .Q(n4405)
         );
  OA221X1 U4353 ( .IN1(n25858), .IN2(n540), .IN3(n25866), .IN4(n583), .IN5(
        n4406), .Q(n4399) );
  OA22X1 U4354 ( .IN1(n25874), .IN2(n626), .IN3(n25882), .IN4(n669), .Q(n4406)
         );
  NAND4X0 U4355 ( .IN1(n4407), .IN2(n4408), .IN3(n4409), .IN4(n4410), .QN(
        n4387) );
  OA221X1 U4356 ( .IN1(n25826), .IN2(n24), .IN3(n25834), .IN4(n67), .IN5(n4411), .Q(n4410) );
  OA22X1 U4357 ( .IN1(n25842), .IN2(n110), .IN3(n25850), .IN4(n153), .Q(n4411)
         );
  OA221X1 U4358 ( .IN1(n25794), .IN2(n196), .IN3(n25802), .IN4(n239), .IN5(
        n4412), .Q(n4409) );
  OA22X1 U4359 ( .IN1(n25810), .IN2(n282), .IN3(n25818), .IN4(n325), .Q(n4412)
         );
  OA221X1 U4360 ( .IN1(n25762), .IN2(n368), .IN3(n25770), .IN4(n411), .IN5(
        n4413), .Q(n4408) );
  OA22X1 U4361 ( .IN1(n25778), .IN2(n454), .IN3(n25786), .IN4(n497), .Q(n4413)
         );
  OA221X1 U4362 ( .IN1(n25730), .IN2(n540), .IN3(n25738), .IN4(n583), .IN5(
        n4414), .Q(n4407) );
  OA22X1 U4363 ( .IN1(n25746), .IN2(n626), .IN3(n25754), .IN4(n669), .Q(n4414)
         );
  NAND4X0 U4364 ( .IN1(n4415), .IN2(n4416), .IN3(n4417), .IN4(n4418), .QN(
        n4386) );
  OA221X1 U4365 ( .IN1(n25698), .IN2(n24), .IN3(n25706), .IN4(n67), .IN5(n4419), .Q(n4418) );
  OA22X1 U4366 ( .IN1(n25714), .IN2(n110), .IN3(n25722), .IN4(n153), .Q(n4419)
         );
  OA221X1 U4367 ( .IN1(n25666), .IN2(n196), .IN3(n25674), .IN4(n239), .IN5(
        n4420), .Q(n4417) );
  OA22X1 U4368 ( .IN1(n25682), .IN2(n282), .IN3(n25690), .IN4(n325), .Q(n4420)
         );
  OA221X1 U4369 ( .IN1(n25634), .IN2(n368), .IN3(n25642), .IN4(n411), .IN5(
        n4421), .Q(n4416) );
  OA22X1 U4370 ( .IN1(n25650), .IN2(n454), .IN3(n25658), .IN4(n497), .Q(n4421)
         );
  OA221X1 U4371 ( .IN1(n25602), .IN2(n540), .IN3(n25610), .IN4(n583), .IN5(
        n4422), .Q(n4415) );
  OA22X1 U4372 ( .IN1(n25618), .IN2(n626), .IN3(n25626), .IN4(n669), .Q(n4422)
         );
  AO221X1 U4373 ( .IN1(n2287), .IN2(n4423), .IN3(n2289), .IN4(n4424), .IN5(
        n4425), .Q(n4346) );
  AO22X1 U4374 ( .IN1(n2292), .IN2(n4426), .IN3(n2294), .IN4(n4427), .Q(n4425)
         );
  NAND4X0 U4375 ( .IN1(n4428), .IN2(n4429), .IN3(n4430), .IN4(n4431), .QN(
        n4427) );
  OA221X1 U4376 ( .IN1(n27618), .IN2(n24), .IN3(n27626), .IN4(n67), .IN5(n4432), .Q(n4431) );
  OA22X1 U4377 ( .IN1(n27634), .IN2(n110), .IN3(n27642), .IN4(n153), .Q(n4432)
         );
  OA221X1 U4378 ( .IN1(n27586), .IN2(n196), .IN3(n27594), .IN4(n239), .IN5(
        n4433), .Q(n4430) );
  OA22X1 U4379 ( .IN1(n27602), .IN2(n282), .IN3(n27610), .IN4(n325), .Q(n4433)
         );
  OA221X1 U4380 ( .IN1(n27554), .IN2(n368), .IN3(n27562), .IN4(n411), .IN5(
        n4434), .Q(n4429) );
  OA22X1 U4381 ( .IN1(n27570), .IN2(n454), .IN3(n27578), .IN4(n497), .Q(n4434)
         );
  OA221X1 U4382 ( .IN1(n27522), .IN2(n540), .IN3(n27530), .IN4(n583), .IN5(
        n4435), .Q(n4428) );
  OA22X1 U4383 ( .IN1(n27538), .IN2(n626), .IN3(n27546), .IN4(n669), .Q(n4435)
         );
  NAND4X0 U4384 ( .IN1(n4436), .IN2(n4437), .IN3(n4438), .IN4(n4439), .QN(
        n4426) );
  OA221X1 U4385 ( .IN1(n27490), .IN2(n24), .IN3(n27498), .IN4(n67), .IN5(n4440), .Q(n4439) );
  OA22X1 U4386 ( .IN1(n27506), .IN2(n110), .IN3(n27514), .IN4(n153), .Q(n4440)
         );
  OA221X1 U4387 ( .IN1(n27458), .IN2(n196), .IN3(n27466), .IN4(n239), .IN5(
        n4441), .Q(n4438) );
  OA22X1 U4388 ( .IN1(n27474), .IN2(n282), .IN3(n27482), .IN4(n325), .Q(n4441)
         );
  OA221X1 U4389 ( .IN1(n27426), .IN2(n368), .IN3(n27434), .IN4(n411), .IN5(
        n4442), .Q(n4437) );
  OA22X1 U4390 ( .IN1(n27442), .IN2(n454), .IN3(n27450), .IN4(n497), .Q(n4442)
         );
  OA221X1 U4391 ( .IN1(n27394), .IN2(n540), .IN3(n27402), .IN4(n583), .IN5(
        n4443), .Q(n4436) );
  OA22X1 U4392 ( .IN1(n27410), .IN2(n626), .IN3(n27418), .IN4(n669), .Q(n4443)
         );
  NAND4X0 U4393 ( .IN1(n4444), .IN2(n4445), .IN3(n4446), .IN4(n4447), .QN(
        n4424) );
  OA221X1 U4394 ( .IN1(n27362), .IN2(n24), .IN3(n27370), .IN4(n67), .IN5(n4448), .Q(n4447) );
  OA22X1 U4395 ( .IN1(n27378), .IN2(n110), .IN3(n27386), .IN4(n153), .Q(n4448)
         );
  OA221X1 U4396 ( .IN1(n27330), .IN2(n196), .IN3(n27338), .IN4(n239), .IN5(
        n4449), .Q(n4446) );
  OA22X1 U4397 ( .IN1(n27346), .IN2(n282), .IN3(n27354), .IN4(n325), .Q(n4449)
         );
  OA221X1 U4398 ( .IN1(n27298), .IN2(n368), .IN3(n27306), .IN4(n411), .IN5(
        n4450), .Q(n4445) );
  OA22X1 U4399 ( .IN1(n27314), .IN2(n454), .IN3(n27322), .IN4(n497), .Q(n4450)
         );
  OA221X1 U4400 ( .IN1(n27266), .IN2(n540), .IN3(n27274), .IN4(n583), .IN5(
        n4451), .Q(n4444) );
  OA22X1 U4401 ( .IN1(n27282), .IN2(n626), .IN3(n27290), .IN4(n669), .Q(n4451)
         );
  NAND4X0 U4402 ( .IN1(n4452), .IN2(n4453), .IN3(n4454), .IN4(n4455), .QN(
        n4423) );
  OA221X1 U4403 ( .IN1(n27234), .IN2(n24), .IN3(n27242), .IN4(n67), .IN5(n4456), .Q(n4455) );
  OA22X1 U4404 ( .IN1(n27250), .IN2(n110), .IN3(n27258), .IN4(n153), .Q(n4456)
         );
  OA221X1 U4405 ( .IN1(n27202), .IN2(n196), .IN3(n27210), .IN4(n239), .IN5(
        n4457), .Q(n4454) );
  OA22X1 U4406 ( .IN1(n27218), .IN2(n282), .IN3(n27226), .IN4(n325), .Q(n4457)
         );
  OA221X1 U4407 ( .IN1(n27170), .IN2(n368), .IN3(n27178), .IN4(n411), .IN5(
        n4458), .Q(n4453) );
  OA22X1 U4408 ( .IN1(n27186), .IN2(n454), .IN3(n27194), .IN4(n497), .Q(n4458)
         );
  OA221X1 U4409 ( .IN1(n27138), .IN2(n540), .IN3(n27146), .IN4(n583), .IN5(
        n4459), .Q(n4452) );
  OA22X1 U4410 ( .IN1(n27154), .IN2(n626), .IN3(n27162), .IN4(n669), .Q(n4459)
         );
  AO221X1 U4411 ( .IN1(n2328), .IN2(n4460), .IN3(n2330), .IN4(n4461), .IN5(
        n4462), .Q(n4345) );
  AO22X1 U4412 ( .IN1(n2333), .IN2(n4463), .IN3(n2335), .IN4(n4464), .Q(n4462)
         );
  NAND4X0 U4413 ( .IN1(n4465), .IN2(n4466), .IN3(n4467), .IN4(n4468), .QN(
        n4464) );
  OA221X1 U4414 ( .IN1(n27106), .IN2(n23), .IN3(n27114), .IN4(n66), .IN5(n4469), .Q(n4468) );
  OA22X1 U4415 ( .IN1(n27122), .IN2(n109), .IN3(n27130), .IN4(n152), .Q(n4469)
         );
  OA221X1 U4416 ( .IN1(n27074), .IN2(n195), .IN3(n27082), .IN4(n238), .IN5(
        n4470), .Q(n4467) );
  OA22X1 U4417 ( .IN1(n27090), .IN2(n281), .IN3(n27098), .IN4(n324), .Q(n4470)
         );
  OA221X1 U4418 ( .IN1(n27042), .IN2(n367), .IN3(n27050), .IN4(n410), .IN5(
        n4471), .Q(n4466) );
  OA22X1 U4419 ( .IN1(n27058), .IN2(n453), .IN3(n27066), .IN4(n496), .Q(n4471)
         );
  OA221X1 U4420 ( .IN1(n27010), .IN2(n539), .IN3(n27018), .IN4(n582), .IN5(
        n4472), .Q(n4465) );
  OA22X1 U4421 ( .IN1(n27026), .IN2(n625), .IN3(n27034), .IN4(n668), .Q(n4472)
         );
  NAND4X0 U4422 ( .IN1(n4473), .IN2(n4474), .IN3(n4475), .IN4(n4476), .QN(
        n4463) );
  OA221X1 U4423 ( .IN1(n26978), .IN2(n23), .IN3(n26986), .IN4(n66), .IN5(n4477), .Q(n4476) );
  OA22X1 U4424 ( .IN1(n26994), .IN2(n109), .IN3(n27002), .IN4(n152), .Q(n4477)
         );
  OA221X1 U4425 ( .IN1(n26946), .IN2(n195), .IN3(n26954), .IN4(n238), .IN5(
        n4478), .Q(n4475) );
  OA22X1 U4426 ( .IN1(n26962), .IN2(n281), .IN3(n26970), .IN4(n324), .Q(n4478)
         );
  OA221X1 U4427 ( .IN1(n26914), .IN2(n367), .IN3(n26922), .IN4(n410), .IN5(
        n4479), .Q(n4474) );
  OA22X1 U4428 ( .IN1(n26930), .IN2(n453), .IN3(n26938), .IN4(n496), .Q(n4479)
         );
  OA221X1 U4429 ( .IN1(n26882), .IN2(n539), .IN3(n26890), .IN4(n582), .IN5(
        n4480), .Q(n4473) );
  OA22X1 U4430 ( .IN1(n26898), .IN2(n625), .IN3(n26906), .IN4(n668), .Q(n4480)
         );
  NAND4X0 U4431 ( .IN1(n4481), .IN2(n4482), .IN3(n4483), .IN4(n4484), .QN(
        n4461) );
  OA221X1 U4432 ( .IN1(n26850), .IN2(n23), .IN3(n26858), .IN4(n66), .IN5(n4485), .Q(n4484) );
  OA22X1 U4433 ( .IN1(n26866), .IN2(n109), .IN3(n26874), .IN4(n152), .Q(n4485)
         );
  OA221X1 U4434 ( .IN1(n26818), .IN2(n195), .IN3(n26826), .IN4(n238), .IN5(
        n4486), .Q(n4483) );
  OA22X1 U4435 ( .IN1(n26834), .IN2(n281), .IN3(n26842), .IN4(n324), .Q(n4486)
         );
  OA221X1 U4436 ( .IN1(n26786), .IN2(n367), .IN3(n26794), .IN4(n410), .IN5(
        n4487), .Q(n4482) );
  OA22X1 U4437 ( .IN1(n26802), .IN2(n453), .IN3(n26810), .IN4(n496), .Q(n4487)
         );
  OA221X1 U4438 ( .IN1(n26754), .IN2(n539), .IN3(n26762), .IN4(n582), .IN5(
        n4488), .Q(n4481) );
  OA22X1 U4439 ( .IN1(n26770), .IN2(n625), .IN3(n26778), .IN4(n668), .Q(n4488)
         );
  NAND4X0 U4440 ( .IN1(n4489), .IN2(n4490), .IN3(n4491), .IN4(n4492), .QN(
        n4460) );
  OA221X1 U4441 ( .IN1(n26722), .IN2(n23), .IN3(n26730), .IN4(n66), .IN5(n4493), .Q(n4492) );
  OA22X1 U4442 ( .IN1(n26738), .IN2(n109), .IN3(n26746), .IN4(n152), .Q(n4493)
         );
  OA221X1 U4443 ( .IN1(n26690), .IN2(n195), .IN3(n26698), .IN4(n238), .IN5(
        n4494), .Q(n4491) );
  OA22X1 U4444 ( .IN1(n26706), .IN2(n281), .IN3(n26714), .IN4(n324), .Q(n4494)
         );
  OA221X1 U4445 ( .IN1(n26658), .IN2(n367), .IN3(n26666), .IN4(n410), .IN5(
        n4495), .Q(n4490) );
  OA22X1 U4446 ( .IN1(n26674), .IN2(n453), .IN3(n26682), .IN4(n496), .Q(n4495)
         );
  OA221X1 U4447 ( .IN1(n26626), .IN2(n539), .IN3(n26634), .IN4(n582), .IN5(
        n4496), .Q(n4489) );
  OA22X1 U4448 ( .IN1(n26642), .IN2(n625), .IN3(n26650), .IN4(n668), .Q(n4496)
         );
  OR4X1 U4449 ( .IN1(n4497), .IN2(n4498), .IN3(n4499), .IN4(n4500), .Q(n2187)
         );
  AO221X1 U4450 ( .IN1(n2157), .IN2(n4501), .IN3(n2159), .IN4(n4502), .IN5(
        n4503), .Q(n4500) );
  AO22X1 U4451 ( .IN1(n2162), .IN2(n4504), .IN3(n2164), .IN4(n4505), .Q(n4503)
         );
  NAND4X0 U4452 ( .IN1(n4506), .IN2(n4507), .IN3(n4508), .IN4(n4509), .QN(
        n4505) );
  OA221X1 U4453 ( .IN1(n26593), .IN2(n23), .IN3(n26601), .IN4(n66), .IN5(n4510), .Q(n4509) );
  OA22X1 U4454 ( .IN1(n26609), .IN2(n109), .IN3(n26617), .IN4(n152), .Q(n4510)
         );
  OA221X1 U4455 ( .IN1(n26561), .IN2(n195), .IN3(n26569), .IN4(n238), .IN5(
        n4511), .Q(n4508) );
  OA22X1 U4456 ( .IN1(n26577), .IN2(n281), .IN3(n26585), .IN4(n324), .Q(n4511)
         );
  OA221X1 U4457 ( .IN1(n26529), .IN2(n367), .IN3(n26537), .IN4(n410), .IN5(
        n4512), .Q(n4507) );
  OA22X1 U4458 ( .IN1(n26545), .IN2(n453), .IN3(n26553), .IN4(n496), .Q(n4512)
         );
  OA221X1 U4459 ( .IN1(n26497), .IN2(n539), .IN3(n26505), .IN4(n582), .IN5(
        n4513), .Q(n4506) );
  OA22X1 U4460 ( .IN1(n26513), .IN2(n625), .IN3(n26521), .IN4(n668), .Q(n4513)
         );
  NAND4X0 U4461 ( .IN1(n4514), .IN2(n4515), .IN3(n4516), .IN4(n4517), .QN(
        n4504) );
  OA221X1 U4462 ( .IN1(n26465), .IN2(n23), .IN3(n26473), .IN4(n66), .IN5(n4518), .Q(n4517) );
  OA22X1 U4463 ( .IN1(n26481), .IN2(n109), .IN3(n26489), .IN4(n152), .Q(n4518)
         );
  OA221X1 U4464 ( .IN1(n26433), .IN2(n195), .IN3(n26441), .IN4(n238), .IN5(
        n4519), .Q(n4516) );
  OA22X1 U4465 ( .IN1(n26449), .IN2(n281), .IN3(n26457), .IN4(n324), .Q(n4519)
         );
  OA221X1 U4466 ( .IN1(n26401), .IN2(n367), .IN3(n26409), .IN4(n410), .IN5(
        n4520), .Q(n4515) );
  OA22X1 U4467 ( .IN1(n26417), .IN2(n453), .IN3(n26425), .IN4(n496), .Q(n4520)
         );
  OA221X1 U4468 ( .IN1(n26369), .IN2(n539), .IN3(n26377), .IN4(n582), .IN5(
        n4521), .Q(n4514) );
  OA22X1 U4469 ( .IN1(n26385), .IN2(n625), .IN3(n26393), .IN4(n668), .Q(n4521)
         );
  NAND4X0 U4470 ( .IN1(n4522), .IN2(n4523), .IN3(n4524), .IN4(n4525), .QN(
        n4502) );
  OA221X1 U4471 ( .IN1(n26337), .IN2(n23), .IN3(n26345), .IN4(n66), .IN5(n4526), .Q(n4525) );
  OA22X1 U4472 ( .IN1(n26353), .IN2(n109), .IN3(n26361), .IN4(n152), .Q(n4526)
         );
  OA221X1 U4473 ( .IN1(n26305), .IN2(n195), .IN3(n26313), .IN4(n238), .IN5(
        n4527), .Q(n4524) );
  OA22X1 U4474 ( .IN1(n26321), .IN2(n281), .IN3(n26329), .IN4(n324), .Q(n4527)
         );
  OA221X1 U4475 ( .IN1(n26273), .IN2(n367), .IN3(n26281), .IN4(n410), .IN5(
        n4528), .Q(n4523) );
  OA22X1 U4476 ( .IN1(n26289), .IN2(n453), .IN3(n26297), .IN4(n496), .Q(n4528)
         );
  OA221X1 U4477 ( .IN1(n26241), .IN2(n539), .IN3(n26249), .IN4(n582), .IN5(
        n4529), .Q(n4522) );
  OA22X1 U4478 ( .IN1(n26257), .IN2(n625), .IN3(n26265), .IN4(n668), .Q(n4529)
         );
  NAND4X0 U4479 ( .IN1(n4530), .IN2(n4531), .IN3(n4532), .IN4(n4533), .QN(
        n4501) );
  OA221X1 U4480 ( .IN1(n26209), .IN2(n23), .IN3(n26217), .IN4(n66), .IN5(n4534), .Q(n4533) );
  OA22X1 U4481 ( .IN1(n26225), .IN2(n109), .IN3(n26233), .IN4(n152), .Q(n4534)
         );
  OA221X1 U4482 ( .IN1(n26177), .IN2(n195), .IN3(n26185), .IN4(n238), .IN5(
        n4535), .Q(n4532) );
  OA22X1 U4483 ( .IN1(n26193), .IN2(n281), .IN3(n26201), .IN4(n324), .Q(n4535)
         );
  OA221X1 U4484 ( .IN1(n26145), .IN2(n367), .IN3(n26153), .IN4(n410), .IN5(
        n4536), .Q(n4531) );
  OA22X1 U4485 ( .IN1(n26161), .IN2(n453), .IN3(n26169), .IN4(n496), .Q(n4536)
         );
  OA221X1 U4486 ( .IN1(n26113), .IN2(n539), .IN3(n26121), .IN4(n582), .IN5(
        n4537), .Q(n4530) );
  OA22X1 U4487 ( .IN1(n26129), .IN2(n625), .IN3(n26137), .IN4(n668), .Q(n4537)
         );
  AO221X1 U4488 ( .IN1(n2246), .IN2(n4538), .IN3(n2248), .IN4(n4539), .IN5(
        n4540), .Q(n4499) );
  AO22X1 U4489 ( .IN1(n2251), .IN2(n4541), .IN3(n2253), .IN4(n4542), .Q(n4540)
         );
  NAND4X0 U4490 ( .IN1(n4543), .IN2(n4544), .IN3(n4545), .IN4(n4546), .QN(
        n4542) );
  OA221X1 U4491 ( .IN1(n26081), .IN2(n23), .IN3(n26089), .IN4(n66), .IN5(n4547), .Q(n4546) );
  OA22X1 U4492 ( .IN1(n26097), .IN2(n109), .IN3(n26105), .IN4(n152), .Q(n4547)
         );
  OA221X1 U4493 ( .IN1(n26049), .IN2(n195), .IN3(n26057), .IN4(n238), .IN5(
        n4548), .Q(n4545) );
  OA22X1 U4494 ( .IN1(n26065), .IN2(n281), .IN3(n26073), .IN4(n324), .Q(n4548)
         );
  OA221X1 U4495 ( .IN1(n26017), .IN2(n367), .IN3(n26025), .IN4(n410), .IN5(
        n4549), .Q(n4544) );
  OA22X1 U4496 ( .IN1(n26033), .IN2(n453), .IN3(n26041), .IN4(n496), .Q(n4549)
         );
  OA221X1 U4497 ( .IN1(n25985), .IN2(n539), .IN3(n25993), .IN4(n582), .IN5(
        n4550), .Q(n4543) );
  OA22X1 U4498 ( .IN1(n26001), .IN2(n625), .IN3(n26009), .IN4(n668), .Q(n4550)
         );
  NAND4X0 U4499 ( .IN1(n4551), .IN2(n4552), .IN3(n4553), .IN4(n4554), .QN(
        n4541) );
  OA221X1 U4500 ( .IN1(n25953), .IN2(n23), .IN3(n25961), .IN4(n66), .IN5(n4555), .Q(n4554) );
  OA22X1 U4501 ( .IN1(n25969), .IN2(n109), .IN3(n25977), .IN4(n152), .Q(n4555)
         );
  OA221X1 U4502 ( .IN1(n25921), .IN2(n195), .IN3(n25929), .IN4(n238), .IN5(
        n4556), .Q(n4553) );
  OA22X1 U4503 ( .IN1(n25937), .IN2(n281), .IN3(n25945), .IN4(n324), .Q(n4556)
         );
  OA221X1 U4504 ( .IN1(n25889), .IN2(n367), .IN3(n25897), .IN4(n410), .IN5(
        n4557), .Q(n4552) );
  OA22X1 U4505 ( .IN1(n25905), .IN2(n453), .IN3(n25913), .IN4(n496), .Q(n4557)
         );
  OA221X1 U4506 ( .IN1(n25857), .IN2(n539), .IN3(n25865), .IN4(n582), .IN5(
        n4558), .Q(n4551) );
  OA22X1 U4507 ( .IN1(n25873), .IN2(n625), .IN3(n25881), .IN4(n668), .Q(n4558)
         );
  NAND4X0 U4508 ( .IN1(n4559), .IN2(n4560), .IN3(n4561), .IN4(n4562), .QN(
        n4539) );
  OA221X1 U4509 ( .IN1(n25825), .IN2(n23), .IN3(n25833), .IN4(n66), .IN5(n4563), .Q(n4562) );
  OA22X1 U4510 ( .IN1(n25841), .IN2(n109), .IN3(n25849), .IN4(n152), .Q(n4563)
         );
  OA221X1 U4511 ( .IN1(n25793), .IN2(n195), .IN3(n25801), .IN4(n238), .IN5(
        n4564), .Q(n4561) );
  OA22X1 U4512 ( .IN1(n25809), .IN2(n281), .IN3(n25817), .IN4(n324), .Q(n4564)
         );
  OA221X1 U4513 ( .IN1(n25761), .IN2(n367), .IN3(n25769), .IN4(n410), .IN5(
        n4565), .Q(n4560) );
  OA22X1 U4514 ( .IN1(n25777), .IN2(n453), .IN3(n25785), .IN4(n496), .Q(n4565)
         );
  OA221X1 U4515 ( .IN1(n25729), .IN2(n539), .IN3(n25737), .IN4(n582), .IN5(
        n4566), .Q(n4559) );
  OA22X1 U4516 ( .IN1(n25745), .IN2(n625), .IN3(n25753), .IN4(n668), .Q(n4566)
         );
  NAND4X0 U4517 ( .IN1(n4567), .IN2(n4568), .IN3(n4569), .IN4(n4570), .QN(
        n4538) );
  OA221X1 U4518 ( .IN1(n25697), .IN2(n23), .IN3(n25705), .IN4(n66), .IN5(n4571), .Q(n4570) );
  OA22X1 U4519 ( .IN1(n25713), .IN2(n109), .IN3(n25721), .IN4(n152), .Q(n4571)
         );
  OA221X1 U4520 ( .IN1(n25665), .IN2(n195), .IN3(n25673), .IN4(n238), .IN5(
        n4572), .Q(n4569) );
  OA22X1 U4521 ( .IN1(n25681), .IN2(n281), .IN3(n25689), .IN4(n324), .Q(n4572)
         );
  OA221X1 U4522 ( .IN1(n25633), .IN2(n367), .IN3(n25641), .IN4(n410), .IN5(
        n4573), .Q(n4568) );
  OA22X1 U4523 ( .IN1(n25649), .IN2(n453), .IN3(n25657), .IN4(n496), .Q(n4573)
         );
  OA221X1 U4524 ( .IN1(n25601), .IN2(n539), .IN3(n25609), .IN4(n582), .IN5(
        n4574), .Q(n4567) );
  OA22X1 U4525 ( .IN1(n25617), .IN2(n625), .IN3(n25625), .IN4(n668), .Q(n4574)
         );
  AO221X1 U4526 ( .IN1(n2287), .IN2(n4575), .IN3(n2289), .IN4(n4576), .IN5(
        n4577), .Q(n4498) );
  AO22X1 U4527 ( .IN1(n2292), .IN2(n4578), .IN3(n2294), .IN4(n4579), .Q(n4577)
         );
  NAND4X0 U4528 ( .IN1(n4580), .IN2(n4581), .IN3(n4582), .IN4(n4583), .QN(
        n4579) );
  OA221X1 U4529 ( .IN1(n27617), .IN2(n22), .IN3(n27625), .IN4(n65), .IN5(n4584), .Q(n4583) );
  OA22X1 U4530 ( .IN1(n27633), .IN2(n108), .IN3(n27641), .IN4(n151), .Q(n4584)
         );
  OA221X1 U4531 ( .IN1(n27585), .IN2(n194), .IN3(n27593), .IN4(n237), .IN5(
        n4585), .Q(n4582) );
  OA22X1 U4532 ( .IN1(n27601), .IN2(n280), .IN3(n27609), .IN4(n323), .Q(n4585)
         );
  OA221X1 U4533 ( .IN1(n27553), .IN2(n366), .IN3(n27561), .IN4(n409), .IN5(
        n4586), .Q(n4581) );
  OA22X1 U4534 ( .IN1(n27569), .IN2(n452), .IN3(n27577), .IN4(n495), .Q(n4586)
         );
  OA221X1 U4535 ( .IN1(n27521), .IN2(n538), .IN3(n27529), .IN4(n581), .IN5(
        n4587), .Q(n4580) );
  OA22X1 U4536 ( .IN1(n27537), .IN2(n624), .IN3(n27545), .IN4(n667), .Q(n4587)
         );
  NAND4X0 U4537 ( .IN1(n4588), .IN2(n4589), .IN3(n4590), .IN4(n4591), .QN(
        n4578) );
  OA221X1 U4538 ( .IN1(n27489), .IN2(n22), .IN3(n27497), .IN4(n65), .IN5(n4592), .Q(n4591) );
  OA22X1 U4539 ( .IN1(n27505), .IN2(n108), .IN3(n27513), .IN4(n151), .Q(n4592)
         );
  OA221X1 U4540 ( .IN1(n27457), .IN2(n194), .IN3(n27465), .IN4(n237), .IN5(
        n4593), .Q(n4590) );
  OA22X1 U4541 ( .IN1(n27473), .IN2(n280), .IN3(n27481), .IN4(n323), .Q(n4593)
         );
  OA221X1 U4542 ( .IN1(n27425), .IN2(n366), .IN3(n27433), .IN4(n409), .IN5(
        n4594), .Q(n4589) );
  OA22X1 U4543 ( .IN1(n27441), .IN2(n452), .IN3(n27449), .IN4(n495), .Q(n4594)
         );
  OA221X1 U4544 ( .IN1(n27393), .IN2(n538), .IN3(n27401), .IN4(n581), .IN5(
        n4595), .Q(n4588) );
  OA22X1 U4545 ( .IN1(n27409), .IN2(n624), .IN3(n27417), .IN4(n667), .Q(n4595)
         );
  NAND4X0 U4546 ( .IN1(n4596), .IN2(n4597), .IN3(n4598), .IN4(n4599), .QN(
        n4576) );
  OA221X1 U4547 ( .IN1(n27361), .IN2(n22), .IN3(n27369), .IN4(n65), .IN5(n4600), .Q(n4599) );
  OA22X1 U4548 ( .IN1(n27377), .IN2(n108), .IN3(n27385), .IN4(n151), .Q(n4600)
         );
  OA221X1 U4549 ( .IN1(n27329), .IN2(n194), .IN3(n27337), .IN4(n237), .IN5(
        n4601), .Q(n4598) );
  OA22X1 U4550 ( .IN1(n27345), .IN2(n280), .IN3(n27353), .IN4(n323), .Q(n4601)
         );
  OA221X1 U4551 ( .IN1(n27297), .IN2(n366), .IN3(n27305), .IN4(n409), .IN5(
        n4602), .Q(n4597) );
  OA22X1 U4552 ( .IN1(n27313), .IN2(n452), .IN3(n27321), .IN4(n495), .Q(n4602)
         );
  OA221X1 U4553 ( .IN1(n27265), .IN2(n538), .IN3(n27273), .IN4(n581), .IN5(
        n4603), .Q(n4596) );
  OA22X1 U4554 ( .IN1(n27281), .IN2(n624), .IN3(n27289), .IN4(n667), .Q(n4603)
         );
  NAND4X0 U4555 ( .IN1(n4604), .IN2(n4605), .IN3(n4606), .IN4(n4607), .QN(
        n4575) );
  OA221X1 U4556 ( .IN1(n27233), .IN2(n22), .IN3(n27241), .IN4(n65), .IN5(n4608), .Q(n4607) );
  OA22X1 U4557 ( .IN1(n27249), .IN2(n108), .IN3(n27257), .IN4(n151), .Q(n4608)
         );
  OA221X1 U4558 ( .IN1(n27201), .IN2(n194), .IN3(n27209), .IN4(n237), .IN5(
        n4609), .Q(n4606) );
  OA22X1 U4559 ( .IN1(n27217), .IN2(n280), .IN3(n27225), .IN4(n323), .Q(n4609)
         );
  OA221X1 U4560 ( .IN1(n27169), .IN2(n366), .IN3(n27177), .IN4(n409), .IN5(
        n4610), .Q(n4605) );
  OA22X1 U4561 ( .IN1(n27185), .IN2(n452), .IN3(n27193), .IN4(n495), .Q(n4610)
         );
  OA221X1 U4562 ( .IN1(n27137), .IN2(n538), .IN3(n27145), .IN4(n581), .IN5(
        n4611), .Q(n4604) );
  OA22X1 U4563 ( .IN1(n27153), .IN2(n624), .IN3(n27161), .IN4(n667), .Q(n4611)
         );
  AO221X1 U4564 ( .IN1(n2328), .IN2(n4612), .IN3(n2330), .IN4(n4613), .IN5(
        n4614), .Q(n4497) );
  AO22X1 U4565 ( .IN1(n2333), .IN2(n4615), .IN3(n2335), .IN4(n4616), .Q(n4614)
         );
  NAND4X0 U4566 ( .IN1(n4617), .IN2(n4618), .IN3(n4619), .IN4(n4620), .QN(
        n4616) );
  OA221X1 U4567 ( .IN1(n27105), .IN2(n22), .IN3(n27113), .IN4(n65), .IN5(n4621), .Q(n4620) );
  OA22X1 U4568 ( .IN1(n27121), .IN2(n108), .IN3(n27129), .IN4(n151), .Q(n4621)
         );
  OA221X1 U4569 ( .IN1(n27073), .IN2(n194), .IN3(n27081), .IN4(n237), .IN5(
        n4622), .Q(n4619) );
  OA22X1 U4570 ( .IN1(n27089), .IN2(n280), .IN3(n27097), .IN4(n323), .Q(n4622)
         );
  OA221X1 U4571 ( .IN1(n27041), .IN2(n366), .IN3(n27049), .IN4(n409), .IN5(
        n4623), .Q(n4618) );
  OA22X1 U4572 ( .IN1(n27057), .IN2(n452), .IN3(n27065), .IN4(n495), .Q(n4623)
         );
  OA221X1 U4573 ( .IN1(n27009), .IN2(n538), .IN3(n27017), .IN4(n581), .IN5(
        n4624), .Q(n4617) );
  OA22X1 U4574 ( .IN1(n27025), .IN2(n624), .IN3(n27033), .IN4(n667), .Q(n4624)
         );
  NAND4X0 U4575 ( .IN1(n4625), .IN2(n4626), .IN3(n4627), .IN4(n4628), .QN(
        n4615) );
  OA221X1 U4576 ( .IN1(n26977), .IN2(n22), .IN3(n26985), .IN4(n65), .IN5(n4629), .Q(n4628) );
  OA22X1 U4577 ( .IN1(n26993), .IN2(n108), .IN3(n27001), .IN4(n151), .Q(n4629)
         );
  OA221X1 U4578 ( .IN1(n26945), .IN2(n194), .IN3(n26953), .IN4(n237), .IN5(
        n4630), .Q(n4627) );
  OA22X1 U4579 ( .IN1(n26961), .IN2(n280), .IN3(n26969), .IN4(n323), .Q(n4630)
         );
  OA221X1 U4580 ( .IN1(n26913), .IN2(n366), .IN3(n26921), .IN4(n409), .IN5(
        n4631), .Q(n4626) );
  OA22X1 U4581 ( .IN1(n26929), .IN2(n452), .IN3(n26937), .IN4(n495), .Q(n4631)
         );
  OA221X1 U4582 ( .IN1(n26881), .IN2(n538), .IN3(n26889), .IN4(n581), .IN5(
        n4632), .Q(n4625) );
  OA22X1 U4583 ( .IN1(n26897), .IN2(n624), .IN3(n26905), .IN4(n667), .Q(n4632)
         );
  NAND4X0 U4584 ( .IN1(n4633), .IN2(n4634), .IN3(n4635), .IN4(n4636), .QN(
        n4613) );
  OA221X1 U4585 ( .IN1(n26849), .IN2(n22), .IN3(n26857), .IN4(n65), .IN5(n4637), .Q(n4636) );
  OA22X1 U4586 ( .IN1(n26865), .IN2(n108), .IN3(n26873), .IN4(n151), .Q(n4637)
         );
  OA221X1 U4587 ( .IN1(n26817), .IN2(n194), .IN3(n26825), .IN4(n237), .IN5(
        n4638), .Q(n4635) );
  OA22X1 U4588 ( .IN1(n26833), .IN2(n280), .IN3(n26841), .IN4(n323), .Q(n4638)
         );
  OA221X1 U4589 ( .IN1(n26785), .IN2(n366), .IN3(n26793), .IN4(n409), .IN5(
        n4639), .Q(n4634) );
  OA22X1 U4590 ( .IN1(n26801), .IN2(n452), .IN3(n26809), .IN4(n495), .Q(n4639)
         );
  OA221X1 U4591 ( .IN1(n26753), .IN2(n538), .IN3(n26761), .IN4(n581), .IN5(
        n4640), .Q(n4633) );
  OA22X1 U4592 ( .IN1(n26769), .IN2(n624), .IN3(n26777), .IN4(n667), .Q(n4640)
         );
  NAND4X0 U4593 ( .IN1(n4641), .IN2(n4642), .IN3(n4643), .IN4(n4644), .QN(
        n4612) );
  OA221X1 U4594 ( .IN1(n26721), .IN2(n22), .IN3(n26729), .IN4(n65), .IN5(n4645), .Q(n4644) );
  OA22X1 U4595 ( .IN1(n26737), .IN2(n108), .IN3(n26745), .IN4(n151), .Q(n4645)
         );
  OA221X1 U4596 ( .IN1(n26689), .IN2(n194), .IN3(n26697), .IN4(n237), .IN5(
        n4646), .Q(n4643) );
  OA22X1 U4597 ( .IN1(n26705), .IN2(n280), .IN3(n26713), .IN4(n323), .Q(n4646)
         );
  OA221X1 U4598 ( .IN1(n26657), .IN2(n366), .IN3(n26665), .IN4(n409), .IN5(
        n4647), .Q(n4642) );
  OA22X1 U4599 ( .IN1(n26673), .IN2(n452), .IN3(n26681), .IN4(n495), .Q(n4647)
         );
  OA221X1 U4600 ( .IN1(n26625), .IN2(n538), .IN3(n26633), .IN4(n581), .IN5(
        n4648), .Q(n4641) );
  OA22X1 U4601 ( .IN1(n26641), .IN2(n624), .IN3(n26649), .IN4(n667), .Q(n4648)
         );
  OR4X1 U4602 ( .IN1(n4649), .IN2(n4650), .IN3(n4651), .IN4(n4652), .Q(n2186)
         );
  AO221X1 U4603 ( .IN1(n2157), .IN2(n4653), .IN3(n2159), .IN4(n4654), .IN5(
        n4655), .Q(n4652) );
  AO22X1 U4604 ( .IN1(n2162), .IN2(n4656), .IN3(n2164), .IN4(n4657), .Q(n4655)
         );
  NAND4X0 U4605 ( .IN1(n4658), .IN2(n4659), .IN3(n4660), .IN4(n4661), .QN(
        n4657) );
  OA221X1 U4606 ( .IN1(n30696), .IN2(n22), .IN3(n30704), .IN4(n65), .IN5(n4662), .Q(n4661) );
  OA22X1 U4607 ( .IN1(n30712), .IN2(n108), .IN3(n30720), .IN4(n151), .Q(n4662)
         );
  OA221X1 U4608 ( .IN1(n30664), .IN2(n194), .IN3(n30672), .IN4(n237), .IN5(
        n4663), .Q(n4660) );
  OA22X1 U4609 ( .IN1(n30680), .IN2(n280), .IN3(n30688), .IN4(n323), .Q(n4663)
         );
  OA221X1 U4610 ( .IN1(n30632), .IN2(n366), .IN3(n30640), .IN4(n409), .IN5(
        n4664), .Q(n4659) );
  OA22X1 U4611 ( .IN1(n30648), .IN2(n452), .IN3(n30656), .IN4(n495), .Q(n4664)
         );
  OA221X1 U4612 ( .IN1(n30600), .IN2(n538), .IN3(n30608), .IN4(n581), .IN5(
        n4665), .Q(n4658) );
  OA22X1 U4613 ( .IN1(n30616), .IN2(n624), .IN3(n30624), .IN4(n667), .Q(n4665)
         );
  NAND4X0 U4614 ( .IN1(n4666), .IN2(n4667), .IN3(n4668), .IN4(n4669), .QN(
        n4656) );
  OA221X1 U4615 ( .IN1(n30568), .IN2(n22), .IN3(n30576), .IN4(n65), .IN5(n4670), .Q(n4669) );
  OA22X1 U4616 ( .IN1(n30584), .IN2(n108), .IN3(n30592), .IN4(n151), .Q(n4670)
         );
  OA221X1 U4617 ( .IN1(n30536), .IN2(n194), .IN3(n30544), .IN4(n237), .IN5(
        n4671), .Q(n4668) );
  OA22X1 U4618 ( .IN1(n30552), .IN2(n280), .IN3(n30560), .IN4(n323), .Q(n4671)
         );
  OA221X1 U4619 ( .IN1(n30504), .IN2(n366), .IN3(n30512), .IN4(n409), .IN5(
        n4672), .Q(n4667) );
  OA22X1 U4620 ( .IN1(n30520), .IN2(n452), .IN3(n30528), .IN4(n495), .Q(n4672)
         );
  OA221X1 U4621 ( .IN1(n30472), .IN2(n538), .IN3(n30480), .IN4(n581), .IN5(
        n4673), .Q(n4666) );
  OA22X1 U4622 ( .IN1(n30488), .IN2(n624), .IN3(n30496), .IN4(n667), .Q(n4673)
         );
  NAND4X0 U4623 ( .IN1(n4674), .IN2(n4675), .IN3(n4676), .IN4(n4677), .QN(
        n4654) );
  OA221X1 U4624 ( .IN1(n30440), .IN2(n22), .IN3(n30448), .IN4(n65), .IN5(n4678), .Q(n4677) );
  OA22X1 U4625 ( .IN1(n30456), .IN2(n108), .IN3(n30464), .IN4(n151), .Q(n4678)
         );
  OA221X1 U4626 ( .IN1(n30408), .IN2(n194), .IN3(n30416), .IN4(n237), .IN5(
        n4679), .Q(n4676) );
  OA22X1 U4627 ( .IN1(n30424), .IN2(n280), .IN3(n30432), .IN4(n323), .Q(n4679)
         );
  OA221X1 U4628 ( .IN1(n30376), .IN2(n366), .IN3(n30384), .IN4(n409), .IN5(
        n4680), .Q(n4675) );
  OA22X1 U4629 ( .IN1(n30392), .IN2(n452), .IN3(n30400), .IN4(n495), .Q(n4680)
         );
  OA221X1 U4630 ( .IN1(n30344), .IN2(n538), .IN3(n30352), .IN4(n581), .IN5(
        n4681), .Q(n4674) );
  OA22X1 U4631 ( .IN1(n30360), .IN2(n624), .IN3(n30368), .IN4(n667), .Q(n4681)
         );
  NAND4X0 U4632 ( .IN1(n4682), .IN2(n4683), .IN3(n4684), .IN4(n4685), .QN(
        n4653) );
  OA221X1 U4633 ( .IN1(n30312), .IN2(n22), .IN3(n30320), .IN4(n65), .IN5(n4686), .Q(n4685) );
  OA22X1 U4634 ( .IN1(n30328), .IN2(n108), .IN3(n30336), .IN4(n151), .Q(n4686)
         );
  OA221X1 U4635 ( .IN1(n30280), .IN2(n194), .IN3(n30288), .IN4(n237), .IN5(
        n4687), .Q(n4684) );
  OA22X1 U4636 ( .IN1(n30296), .IN2(n280), .IN3(n30304), .IN4(n323), .Q(n4687)
         );
  OA221X1 U4637 ( .IN1(n30248), .IN2(n366), .IN3(n30256), .IN4(n409), .IN5(
        n4688), .Q(n4683) );
  OA22X1 U4638 ( .IN1(n30264), .IN2(n452), .IN3(n30272), .IN4(n495), .Q(n4688)
         );
  OA221X1 U4639 ( .IN1(n30216), .IN2(n538), .IN3(n30224), .IN4(n581), .IN5(
        n4689), .Q(n4682) );
  OA22X1 U4640 ( .IN1(n30232), .IN2(n624), .IN3(n30240), .IN4(n667), .Q(n4689)
         );
  AO221X1 U4641 ( .IN1(n2246), .IN2(n4690), .IN3(n2248), .IN4(n4691), .IN5(
        n4692), .Q(n4651) );
  AO22X1 U4642 ( .IN1(n2251), .IN2(n4693), .IN3(n2253), .IN4(n4694), .Q(n4692)
         );
  NAND4X0 U4643 ( .IN1(n4695), .IN2(n4696), .IN3(n4697), .IN4(n4698), .QN(
        n4694) );
  OA221X1 U4644 ( .IN1(n30184), .IN2(n21), .IN3(n30192), .IN4(n64), .IN5(n4699), .Q(n4698) );
  OA22X1 U4645 ( .IN1(n30200), .IN2(n107), .IN3(n30208), .IN4(n150), .Q(n4699)
         );
  OA221X1 U4646 ( .IN1(n30152), .IN2(n193), .IN3(n30160), .IN4(n236), .IN5(
        n4700), .Q(n4697) );
  OA22X1 U4647 ( .IN1(n30168), .IN2(n279), .IN3(n30176), .IN4(n322), .Q(n4700)
         );
  OA221X1 U4648 ( .IN1(n30120), .IN2(n365), .IN3(n30128), .IN4(n408), .IN5(
        n4701), .Q(n4696) );
  OA22X1 U4649 ( .IN1(n30136), .IN2(n451), .IN3(n30144), .IN4(n494), .Q(n4701)
         );
  OA221X1 U4650 ( .IN1(n30088), .IN2(n537), .IN3(n30096), .IN4(n580), .IN5(
        n4702), .Q(n4695) );
  OA22X1 U4651 ( .IN1(n30104), .IN2(n623), .IN3(n30112), .IN4(n666), .Q(n4702)
         );
  NAND4X0 U4652 ( .IN1(n4703), .IN2(n4704), .IN3(n4705), .IN4(n4706), .QN(
        n4693) );
  OA221X1 U4653 ( .IN1(n30056), .IN2(n21), .IN3(n30064), .IN4(n64), .IN5(n4707), .Q(n4706) );
  OA22X1 U4654 ( .IN1(n30072), .IN2(n107), .IN3(n30080), .IN4(n150), .Q(n4707)
         );
  OA221X1 U4655 ( .IN1(n30024), .IN2(n193), .IN3(n30032), .IN4(n236), .IN5(
        n4708), .Q(n4705) );
  OA22X1 U4656 ( .IN1(n30040), .IN2(n279), .IN3(n30048), .IN4(n322), .Q(n4708)
         );
  OA221X1 U4657 ( .IN1(n29992), .IN2(n365), .IN3(n30000), .IN4(n408), .IN5(
        n4709), .Q(n4704) );
  OA22X1 U4658 ( .IN1(n30008), .IN2(n451), .IN3(n30016), .IN4(n494), .Q(n4709)
         );
  OA221X1 U4659 ( .IN1(n29960), .IN2(n537), .IN3(n29968), .IN4(n580), .IN5(
        n4710), .Q(n4703) );
  OA22X1 U4660 ( .IN1(n29976), .IN2(n623), .IN3(n29984), .IN4(n666), .Q(n4710)
         );
  NAND4X0 U4661 ( .IN1(n4711), .IN2(n4712), .IN3(n4713), .IN4(n4714), .QN(
        n4691) );
  OA221X1 U4662 ( .IN1(n29928), .IN2(n21), .IN3(n29936), .IN4(n64), .IN5(n4715), .Q(n4714) );
  OA22X1 U4663 ( .IN1(n29944), .IN2(n107), .IN3(n29952), .IN4(n150), .Q(n4715)
         );
  OA221X1 U4664 ( .IN1(n29896), .IN2(n193), .IN3(n29904), .IN4(n236), .IN5(
        n4716), .Q(n4713) );
  OA22X1 U4665 ( .IN1(n29912), .IN2(n279), .IN3(n29920), .IN4(n322), .Q(n4716)
         );
  OA221X1 U4666 ( .IN1(n29864), .IN2(n365), .IN3(n29872), .IN4(n408), .IN5(
        n4717), .Q(n4712) );
  OA22X1 U4667 ( .IN1(n29880), .IN2(n451), .IN3(n29888), .IN4(n494), .Q(n4717)
         );
  OA221X1 U4668 ( .IN1(n29832), .IN2(n537), .IN3(n29840), .IN4(n580), .IN5(
        n4718), .Q(n4711) );
  OA22X1 U4669 ( .IN1(n29848), .IN2(n623), .IN3(n29856), .IN4(n666), .Q(n4718)
         );
  NAND4X0 U4670 ( .IN1(n4719), .IN2(n4720), .IN3(n4721), .IN4(n4722), .QN(
        n4690) );
  OA221X1 U4671 ( .IN1(n29800), .IN2(n21), .IN3(n29808), .IN4(n64), .IN5(n4723), .Q(n4722) );
  OA22X1 U4672 ( .IN1(n29816), .IN2(n107), .IN3(n29824), .IN4(n150), .Q(n4723)
         );
  OA221X1 U4673 ( .IN1(n29768), .IN2(n193), .IN3(n29776), .IN4(n236), .IN5(
        n4724), .Q(n4721) );
  OA22X1 U4674 ( .IN1(n29784), .IN2(n279), .IN3(n29792), .IN4(n322), .Q(n4724)
         );
  OA221X1 U4675 ( .IN1(n29736), .IN2(n365), .IN3(n29744), .IN4(n408), .IN5(
        n4725), .Q(n4720) );
  OA22X1 U4676 ( .IN1(n29752), .IN2(n451), .IN3(n29760), .IN4(n494), .Q(n4725)
         );
  OA221X1 U4677 ( .IN1(n29704), .IN2(n537), .IN3(n29712), .IN4(n580), .IN5(
        n4726), .Q(n4719) );
  OA22X1 U4678 ( .IN1(n29720), .IN2(n623), .IN3(n29728), .IN4(n666), .Q(n4726)
         );
  AO221X1 U4679 ( .IN1(n2287), .IN2(n4727), .IN3(n2289), .IN4(n4728), .IN5(
        n4729), .Q(n4650) );
  AO22X1 U4680 ( .IN1(n2292), .IN2(n4730), .IN3(n2294), .IN4(n4731), .Q(n4729)
         );
  NAND4X0 U4681 ( .IN1(n4732), .IN2(n4733), .IN3(n4734), .IN4(n4735), .QN(
        n4731) );
  OA221X1 U4682 ( .IN1(n31720), .IN2(n21), .IN3(n31728), .IN4(n64), .IN5(n4736), .Q(n4735) );
  OA22X1 U4683 ( .IN1(n31736), .IN2(n107), .IN3(n31744), .IN4(n150), .Q(n4736)
         );
  OA221X1 U4684 ( .IN1(n31688), .IN2(n193), .IN3(n31696), .IN4(n236), .IN5(
        n4737), .Q(n4734) );
  OA22X1 U4685 ( .IN1(n31704), .IN2(n279), .IN3(n31712), .IN4(n322), .Q(n4737)
         );
  OA221X1 U4686 ( .IN1(n31656), .IN2(n365), .IN3(n31664), .IN4(n408), .IN5(
        n4738), .Q(n4733) );
  OA22X1 U4687 ( .IN1(n31672), .IN2(n451), .IN3(n31680), .IN4(n494), .Q(n4738)
         );
  OA221X1 U4688 ( .IN1(n31624), .IN2(n537), .IN3(n31632), .IN4(n580), .IN5(
        n4739), .Q(n4732) );
  OA22X1 U4689 ( .IN1(n31640), .IN2(n623), .IN3(n31648), .IN4(n666), .Q(n4739)
         );
  NAND4X0 U4690 ( .IN1(n4740), .IN2(n4741), .IN3(n4742), .IN4(n4743), .QN(
        n4730) );
  OA221X1 U4691 ( .IN1(n31592), .IN2(n21), .IN3(n31600), .IN4(n64), .IN5(n4744), .Q(n4743) );
  OA22X1 U4692 ( .IN1(n31608), .IN2(n107), .IN3(n31616), .IN4(n150), .Q(n4744)
         );
  OA221X1 U4693 ( .IN1(n31560), .IN2(n193), .IN3(n31568), .IN4(n236), .IN5(
        n4745), .Q(n4742) );
  OA22X1 U4694 ( .IN1(n31576), .IN2(n279), .IN3(n31584), .IN4(n322), .Q(n4745)
         );
  OA221X1 U4695 ( .IN1(n31528), .IN2(n365), .IN3(n31536), .IN4(n408), .IN5(
        n4746), .Q(n4741) );
  OA22X1 U4696 ( .IN1(n31544), .IN2(n451), .IN3(n31552), .IN4(n494), .Q(n4746)
         );
  OA221X1 U4697 ( .IN1(n31496), .IN2(n537), .IN3(n31504), .IN4(n580), .IN5(
        n4747), .Q(n4740) );
  OA22X1 U4698 ( .IN1(n31512), .IN2(n623), .IN3(n31520), .IN4(n666), .Q(n4747)
         );
  NAND4X0 U4699 ( .IN1(n4748), .IN2(n4749), .IN3(n4750), .IN4(n4751), .QN(
        n4728) );
  OA221X1 U4700 ( .IN1(n31464), .IN2(n21), .IN3(n31472), .IN4(n64), .IN5(n4752), .Q(n4751) );
  OA22X1 U4701 ( .IN1(n31480), .IN2(n107), .IN3(n31488), .IN4(n150), .Q(n4752)
         );
  OA221X1 U4702 ( .IN1(n31432), .IN2(n193), .IN3(n31440), .IN4(n236), .IN5(
        n4753), .Q(n4750) );
  OA22X1 U4703 ( .IN1(n31448), .IN2(n279), .IN3(n31456), .IN4(n322), .Q(n4753)
         );
  OA221X1 U4704 ( .IN1(n31400), .IN2(n365), .IN3(n31408), .IN4(n408), .IN5(
        n4754), .Q(n4749) );
  OA22X1 U4705 ( .IN1(n31416), .IN2(n451), .IN3(n31424), .IN4(n494), .Q(n4754)
         );
  OA221X1 U4706 ( .IN1(n31368), .IN2(n537), .IN3(n31376), .IN4(n580), .IN5(
        n4755), .Q(n4748) );
  OA22X1 U4707 ( .IN1(n31384), .IN2(n623), .IN3(n31392), .IN4(n666), .Q(n4755)
         );
  NAND4X0 U4708 ( .IN1(n4756), .IN2(n4757), .IN3(n4758), .IN4(n4759), .QN(
        n4727) );
  OA221X1 U4709 ( .IN1(n31336), .IN2(n21), .IN3(n31344), .IN4(n64), .IN5(n4760), .Q(n4759) );
  OA22X1 U4710 ( .IN1(n31352), .IN2(n107), .IN3(n31360), .IN4(n150), .Q(n4760)
         );
  OA221X1 U4711 ( .IN1(n31304), .IN2(n193), .IN3(n31312), .IN4(n236), .IN5(
        n4761), .Q(n4758) );
  OA22X1 U4712 ( .IN1(n31320), .IN2(n279), .IN3(n31328), .IN4(n322), .Q(n4761)
         );
  OA221X1 U4713 ( .IN1(n31272), .IN2(n365), .IN3(n31280), .IN4(n408), .IN5(
        n4762), .Q(n4757) );
  OA22X1 U4714 ( .IN1(n31288), .IN2(n451), .IN3(n31296), .IN4(n494), .Q(n4762)
         );
  OA221X1 U4715 ( .IN1(n31240), .IN2(n537), .IN3(n31248), .IN4(n580), .IN5(
        n4763), .Q(n4756) );
  OA22X1 U4716 ( .IN1(n31256), .IN2(n623), .IN3(n31264), .IN4(n666), .Q(n4763)
         );
  AO221X1 U4717 ( .IN1(n2328), .IN2(n4764), .IN3(n2330), .IN4(n4765), .IN5(
        n4766), .Q(n4649) );
  AO22X1 U4718 ( .IN1(n2333), .IN2(n4767), .IN3(n2335), .IN4(n4768), .Q(n4766)
         );
  NAND4X0 U4719 ( .IN1(n4769), .IN2(n4770), .IN3(n4771), .IN4(n4772), .QN(
        n4768) );
  OA221X1 U4720 ( .IN1(n31208), .IN2(n21), .IN3(n31216), .IN4(n64), .IN5(n4773), .Q(n4772) );
  OA22X1 U4721 ( .IN1(n31224), .IN2(n107), .IN3(n31232), .IN4(n150), .Q(n4773)
         );
  OA221X1 U4722 ( .IN1(n31176), .IN2(n193), .IN3(n31184), .IN4(n236), .IN5(
        n4774), .Q(n4771) );
  OA22X1 U4723 ( .IN1(n31192), .IN2(n279), .IN3(n31200), .IN4(n322), .Q(n4774)
         );
  OA221X1 U4724 ( .IN1(n31144), .IN2(n365), .IN3(n31152), .IN4(n408), .IN5(
        n4775), .Q(n4770) );
  OA22X1 U4725 ( .IN1(n31160), .IN2(n451), .IN3(n31168), .IN4(n494), .Q(n4775)
         );
  OA221X1 U4726 ( .IN1(n31112), .IN2(n537), .IN3(n31120), .IN4(n580), .IN5(
        n4776), .Q(n4769) );
  OA22X1 U4727 ( .IN1(n31128), .IN2(n623), .IN3(n31136), .IN4(n666), .Q(n4776)
         );
  NAND4X0 U4728 ( .IN1(n4777), .IN2(n4778), .IN3(n4779), .IN4(n4780), .QN(
        n4767) );
  OA221X1 U4729 ( .IN1(n31080), .IN2(n21), .IN3(n31088), .IN4(n64), .IN5(n4781), .Q(n4780) );
  OA22X1 U4730 ( .IN1(n31096), .IN2(n107), .IN3(n31104), .IN4(n150), .Q(n4781)
         );
  OA221X1 U4731 ( .IN1(n31048), .IN2(n193), .IN3(n31056), .IN4(n236), .IN5(
        n4782), .Q(n4779) );
  OA22X1 U4732 ( .IN1(n31064), .IN2(n279), .IN3(n31072), .IN4(n322), .Q(n4782)
         );
  OA221X1 U4733 ( .IN1(n31016), .IN2(n365), .IN3(n31024), .IN4(n408), .IN5(
        n4783), .Q(n4778) );
  OA22X1 U4734 ( .IN1(n31032), .IN2(n451), .IN3(n31040), .IN4(n494), .Q(n4783)
         );
  OA221X1 U4735 ( .IN1(n30984), .IN2(n537), .IN3(n30992), .IN4(n580), .IN5(
        n4784), .Q(n4777) );
  OA22X1 U4736 ( .IN1(n31000), .IN2(n623), .IN3(n31008), .IN4(n666), .Q(n4784)
         );
  NAND4X0 U4737 ( .IN1(n4785), .IN2(n4786), .IN3(n4787), .IN4(n4788), .QN(
        n4765) );
  OA221X1 U4738 ( .IN1(n30952), .IN2(n21), .IN3(n30960), .IN4(n64), .IN5(n4789), .Q(n4788) );
  OA22X1 U4739 ( .IN1(n30968), .IN2(n107), .IN3(n30976), .IN4(n150), .Q(n4789)
         );
  OA221X1 U4740 ( .IN1(n30920), .IN2(n193), .IN3(n30928), .IN4(n236), .IN5(
        n4790), .Q(n4787) );
  OA22X1 U4741 ( .IN1(n30936), .IN2(n279), .IN3(n30944), .IN4(n322), .Q(n4790)
         );
  OA221X1 U4742 ( .IN1(n30888), .IN2(n365), .IN3(n30896), .IN4(n408), .IN5(
        n4791), .Q(n4786) );
  OA22X1 U4743 ( .IN1(n30904), .IN2(n451), .IN3(n30912), .IN4(n494), .Q(n4791)
         );
  OA221X1 U4744 ( .IN1(n30856), .IN2(n537), .IN3(n30864), .IN4(n580), .IN5(
        n4792), .Q(n4785) );
  OA22X1 U4745 ( .IN1(n30872), .IN2(n623), .IN3(n30880), .IN4(n666), .Q(n4792)
         );
  NAND4X0 U4746 ( .IN1(n4793), .IN2(n4794), .IN3(n4795), .IN4(n4796), .QN(
        n4764) );
  OA221X1 U4747 ( .IN1(n30824), .IN2(n21), .IN3(n30832), .IN4(n64), .IN5(n4797), .Q(n4796) );
  OA22X1 U4748 ( .IN1(n30840), .IN2(n107), .IN3(n30848), .IN4(n150), .Q(n4797)
         );
  OA221X1 U4749 ( .IN1(n30792), .IN2(n193), .IN3(n30800), .IN4(n236), .IN5(
        n4798), .Q(n4795) );
  OA22X1 U4750 ( .IN1(n30808), .IN2(n279), .IN3(n30816), .IN4(n322), .Q(n4798)
         );
  OA221X1 U4751 ( .IN1(n30760), .IN2(n365), .IN3(n30768), .IN4(n408), .IN5(
        n4799), .Q(n4794) );
  OA22X1 U4752 ( .IN1(n30776), .IN2(n451), .IN3(n30784), .IN4(n494), .Q(n4799)
         );
  OA221X1 U4753 ( .IN1(n30728), .IN2(n537), .IN3(n30736), .IN4(n580), .IN5(
        n4800), .Q(n4793) );
  OA22X1 U4754 ( .IN1(n30744), .IN2(n623), .IN3(n30752), .IN4(n666), .Q(n4800)
         );
  OR4X1 U4755 ( .IN1(n4801), .IN2(n4802), .IN3(n4803), .IN4(n4804), .Q(n2185)
         );
  AO221X1 U4756 ( .IN1(n2157), .IN2(n4805), .IN3(n2159), .IN4(n4806), .IN5(
        n4807), .Q(n4804) );
  AO22X1 U4757 ( .IN1(n2162), .IN2(n4808), .IN3(n2164), .IN4(n4809), .Q(n4807)
         );
  NAND4X0 U4758 ( .IN1(n4810), .IN2(n4811), .IN3(n4812), .IN4(n4813), .QN(
        n4809) );
  OA221X1 U4759 ( .IN1(n30695), .IN2(n20), .IN3(n30703), .IN4(n63), .IN5(n4814), .Q(n4813) );
  OA22X1 U4760 ( .IN1(n30711), .IN2(n106), .IN3(n30719), .IN4(n149), .Q(n4814)
         );
  OA221X1 U4761 ( .IN1(n30663), .IN2(n192), .IN3(n30671), .IN4(n235), .IN5(
        n4815), .Q(n4812) );
  OA22X1 U4762 ( .IN1(n30679), .IN2(n278), .IN3(n30687), .IN4(n321), .Q(n4815)
         );
  OA221X1 U4763 ( .IN1(n30631), .IN2(n364), .IN3(n30639), .IN4(n407), .IN5(
        n4816), .Q(n4811) );
  OA22X1 U4764 ( .IN1(n30647), .IN2(n450), .IN3(n30655), .IN4(n493), .Q(n4816)
         );
  OA221X1 U4765 ( .IN1(n30599), .IN2(n536), .IN3(n30607), .IN4(n579), .IN5(
        n4817), .Q(n4810) );
  OA22X1 U4766 ( .IN1(n30615), .IN2(n622), .IN3(n30623), .IN4(n665), .Q(n4817)
         );
  NAND4X0 U4767 ( .IN1(n4818), .IN2(n4819), .IN3(n4820), .IN4(n4821), .QN(
        n4808) );
  OA221X1 U4768 ( .IN1(n30567), .IN2(n20), .IN3(n30575), .IN4(n63), .IN5(n4822), .Q(n4821) );
  OA22X1 U4769 ( .IN1(n30583), .IN2(n106), .IN3(n30591), .IN4(n149), .Q(n4822)
         );
  OA221X1 U4770 ( .IN1(n30535), .IN2(n192), .IN3(n30543), .IN4(n235), .IN5(
        n4823), .Q(n4820) );
  OA22X1 U4771 ( .IN1(n30551), .IN2(n278), .IN3(n30559), .IN4(n321), .Q(n4823)
         );
  OA221X1 U4772 ( .IN1(n30503), .IN2(n364), .IN3(n30511), .IN4(n407), .IN5(
        n4824), .Q(n4819) );
  OA22X1 U4773 ( .IN1(n30519), .IN2(n450), .IN3(n30527), .IN4(n493), .Q(n4824)
         );
  OA221X1 U4774 ( .IN1(n30471), .IN2(n536), .IN3(n30479), .IN4(n579), .IN5(
        n4825), .Q(n4818) );
  OA22X1 U4775 ( .IN1(n30487), .IN2(n622), .IN3(n30495), .IN4(n665), .Q(n4825)
         );
  NAND4X0 U4776 ( .IN1(n4826), .IN2(n4827), .IN3(n4828), .IN4(n4829), .QN(
        n4806) );
  OA221X1 U4777 ( .IN1(n30439), .IN2(n20), .IN3(n30447), .IN4(n63), .IN5(n4830), .Q(n4829) );
  OA22X1 U4778 ( .IN1(n30455), .IN2(n106), .IN3(n30463), .IN4(n149), .Q(n4830)
         );
  OA221X1 U4779 ( .IN1(n30407), .IN2(n192), .IN3(n30415), .IN4(n235), .IN5(
        n4831), .Q(n4828) );
  OA22X1 U4780 ( .IN1(n30423), .IN2(n278), .IN3(n30431), .IN4(n321), .Q(n4831)
         );
  OA221X1 U4781 ( .IN1(n30375), .IN2(n364), .IN3(n30383), .IN4(n407), .IN5(
        n4832), .Q(n4827) );
  OA22X1 U4782 ( .IN1(n30391), .IN2(n450), .IN3(n30399), .IN4(n493), .Q(n4832)
         );
  OA221X1 U4783 ( .IN1(n30343), .IN2(n536), .IN3(n30351), .IN4(n579), .IN5(
        n4833), .Q(n4826) );
  OA22X1 U4784 ( .IN1(n30359), .IN2(n622), .IN3(n30367), .IN4(n665), .Q(n4833)
         );
  NAND4X0 U4785 ( .IN1(n4834), .IN2(n4835), .IN3(n4836), .IN4(n4837), .QN(
        n4805) );
  OA221X1 U4786 ( .IN1(n30311), .IN2(n20), .IN3(n30319), .IN4(n63), .IN5(n4838), .Q(n4837) );
  OA22X1 U4787 ( .IN1(n30327), .IN2(n106), .IN3(n30335), .IN4(n149), .Q(n4838)
         );
  OA221X1 U4788 ( .IN1(n30279), .IN2(n192), .IN3(n30287), .IN4(n235), .IN5(
        n4839), .Q(n4836) );
  OA22X1 U4789 ( .IN1(n30295), .IN2(n278), .IN3(n30303), .IN4(n321), .Q(n4839)
         );
  OA221X1 U4790 ( .IN1(n30247), .IN2(n364), .IN3(n30255), .IN4(n407), .IN5(
        n4840), .Q(n4835) );
  OA22X1 U4791 ( .IN1(n30263), .IN2(n450), .IN3(n30271), .IN4(n493), .Q(n4840)
         );
  OA221X1 U4792 ( .IN1(n30215), .IN2(n536), .IN3(n30223), .IN4(n579), .IN5(
        n4841), .Q(n4834) );
  OA22X1 U4793 ( .IN1(n30231), .IN2(n622), .IN3(n30239), .IN4(n665), .Q(n4841)
         );
  AO221X1 U4794 ( .IN1(n2246), .IN2(n4842), .IN3(n2248), .IN4(n4843), .IN5(
        n4844), .Q(n4803) );
  AO22X1 U4795 ( .IN1(n2251), .IN2(n4845), .IN3(n2253), .IN4(n4846), .Q(n4844)
         );
  NAND4X0 U4796 ( .IN1(n4847), .IN2(n4848), .IN3(n4849), .IN4(n4850), .QN(
        n4846) );
  OA221X1 U4797 ( .IN1(n30183), .IN2(n20), .IN3(n30191), .IN4(n63), .IN5(n4851), .Q(n4850) );
  OA22X1 U4798 ( .IN1(n30199), .IN2(n106), .IN3(n30207), .IN4(n149), .Q(n4851)
         );
  OA221X1 U4799 ( .IN1(n30151), .IN2(n192), .IN3(n30159), .IN4(n235), .IN5(
        n4852), .Q(n4849) );
  OA22X1 U4800 ( .IN1(n30167), .IN2(n278), .IN3(n30175), .IN4(n321), .Q(n4852)
         );
  OA221X1 U4801 ( .IN1(n30119), .IN2(n364), .IN3(n30127), .IN4(n407), .IN5(
        n4853), .Q(n4848) );
  OA22X1 U4802 ( .IN1(n30135), .IN2(n450), .IN3(n30143), .IN4(n493), .Q(n4853)
         );
  OA221X1 U4803 ( .IN1(n30087), .IN2(n536), .IN3(n30095), .IN4(n579), .IN5(
        n4854), .Q(n4847) );
  OA22X1 U4804 ( .IN1(n30103), .IN2(n622), .IN3(n30111), .IN4(n665), .Q(n4854)
         );
  NAND4X0 U4805 ( .IN1(n4855), .IN2(n4856), .IN3(n4857), .IN4(n4858), .QN(
        n4845) );
  OA221X1 U4806 ( .IN1(n30055), .IN2(n20), .IN3(n30063), .IN4(n63), .IN5(n4859), .Q(n4858) );
  OA22X1 U4807 ( .IN1(n30071), .IN2(n106), .IN3(n30079), .IN4(n149), .Q(n4859)
         );
  OA221X1 U4808 ( .IN1(n30023), .IN2(n192), .IN3(n30031), .IN4(n235), .IN5(
        n4860), .Q(n4857) );
  OA22X1 U4809 ( .IN1(n30039), .IN2(n278), .IN3(n30047), .IN4(n321), .Q(n4860)
         );
  OA221X1 U4810 ( .IN1(n29991), .IN2(n364), .IN3(n29999), .IN4(n407), .IN5(
        n4861), .Q(n4856) );
  OA22X1 U4811 ( .IN1(n30007), .IN2(n450), .IN3(n30015), .IN4(n493), .Q(n4861)
         );
  OA221X1 U4812 ( .IN1(n29959), .IN2(n536), .IN3(n29967), .IN4(n579), .IN5(
        n4862), .Q(n4855) );
  OA22X1 U4813 ( .IN1(n29975), .IN2(n622), .IN3(n29983), .IN4(n665), .Q(n4862)
         );
  NAND4X0 U4814 ( .IN1(n4863), .IN2(n4864), .IN3(n4865), .IN4(n4866), .QN(
        n4843) );
  OA221X1 U4815 ( .IN1(n29927), .IN2(n20), .IN3(n29935), .IN4(n63), .IN5(n4867), .Q(n4866) );
  OA22X1 U4816 ( .IN1(n29943), .IN2(n106), .IN3(n29951), .IN4(n149), .Q(n4867)
         );
  OA221X1 U4817 ( .IN1(n29895), .IN2(n192), .IN3(n29903), .IN4(n235), .IN5(
        n4868), .Q(n4865) );
  OA22X1 U4818 ( .IN1(n29911), .IN2(n278), .IN3(n29919), .IN4(n321), .Q(n4868)
         );
  OA221X1 U4819 ( .IN1(n29863), .IN2(n364), .IN3(n29871), .IN4(n407), .IN5(
        n4869), .Q(n4864) );
  OA22X1 U4820 ( .IN1(n29879), .IN2(n450), .IN3(n29887), .IN4(n493), .Q(n4869)
         );
  OA221X1 U4821 ( .IN1(n29831), .IN2(n536), .IN3(n29839), .IN4(n579), .IN5(
        n4870), .Q(n4863) );
  OA22X1 U4822 ( .IN1(n29847), .IN2(n622), .IN3(n29855), .IN4(n665), .Q(n4870)
         );
  NAND4X0 U4823 ( .IN1(n4871), .IN2(n4872), .IN3(n4873), .IN4(n4874), .QN(
        n4842) );
  OA221X1 U4824 ( .IN1(n29799), .IN2(n20), .IN3(n29807), .IN4(n63), .IN5(n4875), .Q(n4874) );
  OA22X1 U4825 ( .IN1(n29815), .IN2(n106), .IN3(n29823), .IN4(n149), .Q(n4875)
         );
  OA221X1 U4826 ( .IN1(n29767), .IN2(n192), .IN3(n29775), .IN4(n235), .IN5(
        n4876), .Q(n4873) );
  OA22X1 U4827 ( .IN1(n29783), .IN2(n278), .IN3(n29791), .IN4(n321), .Q(n4876)
         );
  OA221X1 U4828 ( .IN1(n29735), .IN2(n364), .IN3(n29743), .IN4(n407), .IN5(
        n4877), .Q(n4872) );
  OA22X1 U4829 ( .IN1(n29751), .IN2(n450), .IN3(n29759), .IN4(n493), .Q(n4877)
         );
  OA221X1 U4830 ( .IN1(n29703), .IN2(n536), .IN3(n29711), .IN4(n579), .IN5(
        n4878), .Q(n4871) );
  OA22X1 U4831 ( .IN1(n29719), .IN2(n622), .IN3(n29727), .IN4(n665), .Q(n4878)
         );
  AO221X1 U4832 ( .IN1(n2287), .IN2(n4879), .IN3(n2289), .IN4(n4880), .IN5(
        n4881), .Q(n4802) );
  AO22X1 U4833 ( .IN1(n2292), .IN2(n4882), .IN3(n2294), .IN4(n4883), .Q(n4881)
         );
  NAND4X0 U4834 ( .IN1(n4884), .IN2(n4885), .IN3(n4886), .IN4(n4887), .QN(
        n4883) );
  OA221X1 U4835 ( .IN1(n31719), .IN2(n20), .IN3(n31727), .IN4(n63), .IN5(n4888), .Q(n4887) );
  OA22X1 U4836 ( .IN1(n31735), .IN2(n106), .IN3(n31743), .IN4(n149), .Q(n4888)
         );
  OA221X1 U4837 ( .IN1(n31687), .IN2(n192), .IN3(n31695), .IN4(n235), .IN5(
        n4889), .Q(n4886) );
  OA22X1 U4838 ( .IN1(n31703), .IN2(n278), .IN3(n31711), .IN4(n321), .Q(n4889)
         );
  OA221X1 U4839 ( .IN1(n31655), .IN2(n364), .IN3(n31663), .IN4(n407), .IN5(
        n4890), .Q(n4885) );
  OA22X1 U4840 ( .IN1(n31671), .IN2(n450), .IN3(n31679), .IN4(n493), .Q(n4890)
         );
  OA221X1 U4841 ( .IN1(n31623), .IN2(n536), .IN3(n31631), .IN4(n579), .IN5(
        n4891), .Q(n4884) );
  OA22X1 U4842 ( .IN1(n31639), .IN2(n622), .IN3(n31647), .IN4(n665), .Q(n4891)
         );
  NAND4X0 U4843 ( .IN1(n4892), .IN2(n4893), .IN3(n4894), .IN4(n4895), .QN(
        n4882) );
  OA221X1 U4844 ( .IN1(n31591), .IN2(n20), .IN3(n31599), .IN4(n63), .IN5(n4896), .Q(n4895) );
  OA22X1 U4845 ( .IN1(n31607), .IN2(n106), .IN3(n31615), .IN4(n149), .Q(n4896)
         );
  OA221X1 U4846 ( .IN1(n31559), .IN2(n192), .IN3(n31567), .IN4(n235), .IN5(
        n4897), .Q(n4894) );
  OA22X1 U4847 ( .IN1(n31575), .IN2(n278), .IN3(n31583), .IN4(n321), .Q(n4897)
         );
  OA221X1 U4848 ( .IN1(n31527), .IN2(n364), .IN3(n31535), .IN4(n407), .IN5(
        n4898), .Q(n4893) );
  OA22X1 U4849 ( .IN1(n31543), .IN2(n450), .IN3(n31551), .IN4(n493), .Q(n4898)
         );
  OA221X1 U4850 ( .IN1(n31495), .IN2(n536), .IN3(n31503), .IN4(n579), .IN5(
        n4899), .Q(n4892) );
  OA22X1 U4851 ( .IN1(n31511), .IN2(n622), .IN3(n31519), .IN4(n665), .Q(n4899)
         );
  NAND4X0 U4852 ( .IN1(n4900), .IN2(n4901), .IN3(n4902), .IN4(n4903), .QN(
        n4880) );
  OA221X1 U4853 ( .IN1(n31463), .IN2(n20), .IN3(n31471), .IN4(n63), .IN5(n4904), .Q(n4903) );
  OA22X1 U4854 ( .IN1(n31479), .IN2(n106), .IN3(n31487), .IN4(n149), .Q(n4904)
         );
  OA221X1 U4855 ( .IN1(n31431), .IN2(n192), .IN3(n31439), .IN4(n235), .IN5(
        n4905), .Q(n4902) );
  OA22X1 U4856 ( .IN1(n31447), .IN2(n278), .IN3(n31455), .IN4(n321), .Q(n4905)
         );
  OA221X1 U4857 ( .IN1(n31399), .IN2(n364), .IN3(n31407), .IN4(n407), .IN5(
        n4906), .Q(n4901) );
  OA22X1 U4858 ( .IN1(n31415), .IN2(n450), .IN3(n31423), .IN4(n493), .Q(n4906)
         );
  OA221X1 U4859 ( .IN1(n31367), .IN2(n536), .IN3(n31375), .IN4(n579), .IN5(
        n4907), .Q(n4900) );
  OA22X1 U4860 ( .IN1(n31383), .IN2(n622), .IN3(n31391), .IN4(n665), .Q(n4907)
         );
  NAND4X0 U4861 ( .IN1(n4908), .IN2(n4909), .IN3(n4910), .IN4(n4911), .QN(
        n4879) );
  OA221X1 U4862 ( .IN1(n31335), .IN2(n20), .IN3(n31343), .IN4(n63), .IN5(n4912), .Q(n4911) );
  OA22X1 U4863 ( .IN1(n31351), .IN2(n106), .IN3(n31359), .IN4(n149), .Q(n4912)
         );
  OA221X1 U4864 ( .IN1(n31303), .IN2(n192), .IN3(n31311), .IN4(n235), .IN5(
        n4913), .Q(n4910) );
  OA22X1 U4865 ( .IN1(n31319), .IN2(n278), .IN3(n31327), .IN4(n321), .Q(n4913)
         );
  OA221X1 U4866 ( .IN1(n31271), .IN2(n364), .IN3(n31279), .IN4(n407), .IN5(
        n4914), .Q(n4909) );
  OA22X1 U4867 ( .IN1(n31287), .IN2(n450), .IN3(n31295), .IN4(n493), .Q(n4914)
         );
  OA221X1 U4868 ( .IN1(n31239), .IN2(n536), .IN3(n31247), .IN4(n579), .IN5(
        n4915), .Q(n4908) );
  OA22X1 U4869 ( .IN1(n31255), .IN2(n622), .IN3(n31263), .IN4(n665), .Q(n4915)
         );
  AO221X1 U4870 ( .IN1(n2328), .IN2(n4916), .IN3(n2330), .IN4(n4917), .IN5(
        n4918), .Q(n4801) );
  AO22X1 U4871 ( .IN1(n2333), .IN2(n4919), .IN3(n2335), .IN4(n4920), .Q(n4918)
         );
  NAND4X0 U4872 ( .IN1(n4921), .IN2(n4922), .IN3(n4923), .IN4(n4924), .QN(
        n4920) );
  OA221X1 U4873 ( .IN1(n31207), .IN2(n19), .IN3(n31215), .IN4(n62), .IN5(n4925), .Q(n4924) );
  OA22X1 U4874 ( .IN1(n31223), .IN2(n105), .IN3(n31231), .IN4(n148), .Q(n4925)
         );
  OA221X1 U4875 ( .IN1(n31175), .IN2(n191), .IN3(n31183), .IN4(n234), .IN5(
        n4926), .Q(n4923) );
  OA22X1 U4876 ( .IN1(n31191), .IN2(n277), .IN3(n31199), .IN4(n320), .Q(n4926)
         );
  OA221X1 U4877 ( .IN1(n31143), .IN2(n363), .IN3(n31151), .IN4(n406), .IN5(
        n4927), .Q(n4922) );
  OA22X1 U4878 ( .IN1(n31159), .IN2(n449), .IN3(n31167), .IN4(n492), .Q(n4927)
         );
  OA221X1 U4879 ( .IN1(n31111), .IN2(n535), .IN3(n31119), .IN4(n578), .IN5(
        n4928), .Q(n4921) );
  OA22X1 U4880 ( .IN1(n31127), .IN2(n621), .IN3(n31135), .IN4(n664), .Q(n4928)
         );
  NAND4X0 U4881 ( .IN1(n4929), .IN2(n4930), .IN3(n4931), .IN4(n4932), .QN(
        n4919) );
  OA221X1 U4882 ( .IN1(n31079), .IN2(n19), .IN3(n31087), .IN4(n62), .IN5(n4933), .Q(n4932) );
  OA22X1 U4883 ( .IN1(n31095), .IN2(n105), .IN3(n31103), .IN4(n148), .Q(n4933)
         );
  OA221X1 U4884 ( .IN1(n31047), .IN2(n191), .IN3(n31055), .IN4(n234), .IN5(
        n4934), .Q(n4931) );
  OA22X1 U4885 ( .IN1(n31063), .IN2(n277), .IN3(n31071), .IN4(n320), .Q(n4934)
         );
  OA221X1 U4886 ( .IN1(n31015), .IN2(n363), .IN3(n31023), .IN4(n406), .IN5(
        n4935), .Q(n4930) );
  OA22X1 U4887 ( .IN1(n31031), .IN2(n449), .IN3(n31039), .IN4(n492), .Q(n4935)
         );
  OA221X1 U4888 ( .IN1(n30983), .IN2(n535), .IN3(n30991), .IN4(n578), .IN5(
        n4936), .Q(n4929) );
  OA22X1 U4889 ( .IN1(n30999), .IN2(n621), .IN3(n31007), .IN4(n664), .Q(n4936)
         );
  NAND4X0 U4890 ( .IN1(n4937), .IN2(n4938), .IN3(n4939), .IN4(n4940), .QN(
        n4917) );
  OA221X1 U4891 ( .IN1(n30951), .IN2(n19), .IN3(n30959), .IN4(n62), .IN5(n4941), .Q(n4940) );
  OA22X1 U4892 ( .IN1(n30967), .IN2(n105), .IN3(n30975), .IN4(n148), .Q(n4941)
         );
  OA221X1 U4893 ( .IN1(n30919), .IN2(n191), .IN3(n30927), .IN4(n234), .IN5(
        n4942), .Q(n4939) );
  OA22X1 U4894 ( .IN1(n30935), .IN2(n277), .IN3(n30943), .IN4(n320), .Q(n4942)
         );
  OA221X1 U4895 ( .IN1(n30887), .IN2(n363), .IN3(n30895), .IN4(n406), .IN5(
        n4943), .Q(n4938) );
  OA22X1 U4896 ( .IN1(n30903), .IN2(n449), .IN3(n30911), .IN4(n492), .Q(n4943)
         );
  OA221X1 U4897 ( .IN1(n30855), .IN2(n535), .IN3(n30863), .IN4(n578), .IN5(
        n4944), .Q(n4937) );
  OA22X1 U4898 ( .IN1(n30871), .IN2(n621), .IN3(n30879), .IN4(n664), .Q(n4944)
         );
  NAND4X0 U4899 ( .IN1(n4945), .IN2(n4946), .IN3(n4947), .IN4(n4948), .QN(
        n4916) );
  OA221X1 U4900 ( .IN1(n30823), .IN2(n19), .IN3(n30831), .IN4(n62), .IN5(n4949), .Q(n4948) );
  OA22X1 U4901 ( .IN1(n30839), .IN2(n105), .IN3(n30847), .IN4(n148), .Q(n4949)
         );
  OA221X1 U4902 ( .IN1(n30791), .IN2(n191), .IN3(n30799), .IN4(n234), .IN5(
        n4950), .Q(n4947) );
  OA22X1 U4903 ( .IN1(n30807), .IN2(n277), .IN3(n30815), .IN4(n320), .Q(n4950)
         );
  OA221X1 U4904 ( .IN1(n30759), .IN2(n363), .IN3(n30767), .IN4(n406), .IN5(
        n4951), .Q(n4946) );
  OA22X1 U4905 ( .IN1(n30775), .IN2(n449), .IN3(n30783), .IN4(n492), .Q(n4951)
         );
  OA221X1 U4906 ( .IN1(n30727), .IN2(n535), .IN3(n30735), .IN4(n578), .IN5(
        n4952), .Q(n4945) );
  OA22X1 U4907 ( .IN1(n30743), .IN2(n621), .IN3(n30751), .IN4(n664), .Q(n4952)
         );
  OR4X1 U4908 ( .IN1(n4953), .IN2(n4954), .IN3(n4955), .IN4(n4956), .Q(n2184)
         );
  AO221X1 U4909 ( .IN1(n2157), .IN2(n4957), .IN3(n2159), .IN4(n4958), .IN5(
        n4959), .Q(n4956) );
  AO22X1 U4910 ( .IN1(n2162), .IN2(n4960), .IN3(n2164), .IN4(n4961), .Q(n4959)
         );
  NAND4X0 U4911 ( .IN1(n4962), .IN2(n4963), .IN3(n4964), .IN4(n4965), .QN(
        n4961) );
  OA221X1 U4912 ( .IN1(n30694), .IN2(n19), .IN3(n30702), .IN4(n62), .IN5(n4966), .Q(n4965) );
  OA22X1 U4913 ( .IN1(n30710), .IN2(n105), .IN3(n30718), .IN4(n148), .Q(n4966)
         );
  OA221X1 U4914 ( .IN1(n30662), .IN2(n191), .IN3(n30670), .IN4(n234), .IN5(
        n4967), .Q(n4964) );
  OA22X1 U4915 ( .IN1(n30678), .IN2(n277), .IN3(n30686), .IN4(n320), .Q(n4967)
         );
  OA221X1 U4916 ( .IN1(n30630), .IN2(n363), .IN3(n30638), .IN4(n406), .IN5(
        n4968), .Q(n4963) );
  OA22X1 U4917 ( .IN1(n30646), .IN2(n449), .IN3(n30654), .IN4(n492), .Q(n4968)
         );
  OA221X1 U4918 ( .IN1(n30598), .IN2(n535), .IN3(n30606), .IN4(n578), .IN5(
        n4969), .Q(n4962) );
  OA22X1 U4919 ( .IN1(n30614), .IN2(n621), .IN3(n30622), .IN4(n664), .Q(n4969)
         );
  NAND4X0 U4920 ( .IN1(n4970), .IN2(n4971), .IN3(n4972), .IN4(n4973), .QN(
        n4960) );
  OA221X1 U4921 ( .IN1(n30566), .IN2(n19), .IN3(n30574), .IN4(n62), .IN5(n4974), .Q(n4973) );
  OA22X1 U4922 ( .IN1(n30582), .IN2(n105), .IN3(n30590), .IN4(n148), .Q(n4974)
         );
  OA221X1 U4923 ( .IN1(n30534), .IN2(n191), .IN3(n30542), .IN4(n234), .IN5(
        n4975), .Q(n4972) );
  OA22X1 U4924 ( .IN1(n30550), .IN2(n277), .IN3(n30558), .IN4(n320), .Q(n4975)
         );
  OA221X1 U4925 ( .IN1(n30502), .IN2(n363), .IN3(n30510), .IN4(n406), .IN5(
        n4976), .Q(n4971) );
  OA22X1 U4926 ( .IN1(n30518), .IN2(n449), .IN3(n30526), .IN4(n492), .Q(n4976)
         );
  OA221X1 U4927 ( .IN1(n30470), .IN2(n535), .IN3(n30478), .IN4(n578), .IN5(
        n4977), .Q(n4970) );
  OA22X1 U4928 ( .IN1(n30486), .IN2(n621), .IN3(n30494), .IN4(n664), .Q(n4977)
         );
  NAND4X0 U4929 ( .IN1(n4978), .IN2(n4979), .IN3(n4980), .IN4(n4981), .QN(
        n4958) );
  OA221X1 U4930 ( .IN1(n30438), .IN2(n19), .IN3(n30446), .IN4(n62), .IN5(n4982), .Q(n4981) );
  OA22X1 U4931 ( .IN1(n30454), .IN2(n105), .IN3(n30462), .IN4(n148), .Q(n4982)
         );
  OA221X1 U4932 ( .IN1(n30406), .IN2(n191), .IN3(n30414), .IN4(n234), .IN5(
        n4983), .Q(n4980) );
  OA22X1 U4933 ( .IN1(n30422), .IN2(n277), .IN3(n30430), .IN4(n320), .Q(n4983)
         );
  OA221X1 U4934 ( .IN1(n30374), .IN2(n363), .IN3(n30382), .IN4(n406), .IN5(
        n4984), .Q(n4979) );
  OA22X1 U4935 ( .IN1(n30390), .IN2(n449), .IN3(n30398), .IN4(n492), .Q(n4984)
         );
  OA221X1 U4936 ( .IN1(n30342), .IN2(n535), .IN3(n30350), .IN4(n578), .IN5(
        n4985), .Q(n4978) );
  OA22X1 U4937 ( .IN1(n30358), .IN2(n621), .IN3(n30366), .IN4(n664), .Q(n4985)
         );
  NAND4X0 U4938 ( .IN1(n4986), .IN2(n4987), .IN3(n4988), .IN4(n4989), .QN(
        n4957) );
  OA221X1 U4939 ( .IN1(n30310), .IN2(n19), .IN3(n30318), .IN4(n62), .IN5(n4990), .Q(n4989) );
  OA22X1 U4940 ( .IN1(n30326), .IN2(n105), .IN3(n30334), .IN4(n148), .Q(n4990)
         );
  OA221X1 U4941 ( .IN1(n30278), .IN2(n191), .IN3(n30286), .IN4(n234), .IN5(
        n4991), .Q(n4988) );
  OA22X1 U4942 ( .IN1(n30294), .IN2(n277), .IN3(n30302), .IN4(n320), .Q(n4991)
         );
  OA221X1 U4943 ( .IN1(n30246), .IN2(n363), .IN3(n30254), .IN4(n406), .IN5(
        n4992), .Q(n4987) );
  OA22X1 U4944 ( .IN1(n30262), .IN2(n449), .IN3(n30270), .IN4(n492), .Q(n4992)
         );
  OA221X1 U4945 ( .IN1(n30214), .IN2(n535), .IN3(n30222), .IN4(n578), .IN5(
        n4993), .Q(n4986) );
  OA22X1 U4946 ( .IN1(n30230), .IN2(n621), .IN3(n30238), .IN4(n664), .Q(n4993)
         );
  AO221X1 U4947 ( .IN1(n2246), .IN2(n4994), .IN3(n2248), .IN4(n4995), .IN5(
        n4996), .Q(n4955) );
  AO22X1 U4948 ( .IN1(n2251), .IN2(n4997), .IN3(n2253), .IN4(n4998), .Q(n4996)
         );
  NAND4X0 U4949 ( .IN1(n4999), .IN2(n5000), .IN3(n5001), .IN4(n5002), .QN(
        n4998) );
  OA221X1 U4950 ( .IN1(n30182), .IN2(n19), .IN3(n30190), .IN4(n62), .IN5(n5003), .Q(n5002) );
  OA22X1 U4951 ( .IN1(n30198), .IN2(n105), .IN3(n30206), .IN4(n148), .Q(n5003)
         );
  OA221X1 U4952 ( .IN1(n30150), .IN2(n191), .IN3(n30158), .IN4(n234), .IN5(
        n5004), .Q(n5001) );
  OA22X1 U4953 ( .IN1(n30166), .IN2(n277), .IN3(n30174), .IN4(n320), .Q(n5004)
         );
  OA221X1 U4954 ( .IN1(n30118), .IN2(n363), .IN3(n30126), .IN4(n406), .IN5(
        n5005), .Q(n5000) );
  OA22X1 U4955 ( .IN1(n30134), .IN2(n449), .IN3(n30142), .IN4(n492), .Q(n5005)
         );
  OA221X1 U4956 ( .IN1(n30086), .IN2(n535), .IN3(n30094), .IN4(n578), .IN5(
        n5006), .Q(n4999) );
  OA22X1 U4957 ( .IN1(n30102), .IN2(n621), .IN3(n30110), .IN4(n664), .Q(n5006)
         );
  NAND4X0 U4958 ( .IN1(n5007), .IN2(n5008), .IN3(n5009), .IN4(n5010), .QN(
        n4997) );
  OA221X1 U4959 ( .IN1(n30054), .IN2(n19), .IN3(n30062), .IN4(n62), .IN5(n5011), .Q(n5010) );
  OA22X1 U4960 ( .IN1(n30070), .IN2(n105), .IN3(n30078), .IN4(n148), .Q(n5011)
         );
  OA221X1 U4961 ( .IN1(n30022), .IN2(n191), .IN3(n30030), .IN4(n234), .IN5(
        n5012), .Q(n5009) );
  OA22X1 U4962 ( .IN1(n30038), .IN2(n277), .IN3(n30046), .IN4(n320), .Q(n5012)
         );
  OA221X1 U4963 ( .IN1(n29990), .IN2(n363), .IN3(n29998), .IN4(n406), .IN5(
        n5013), .Q(n5008) );
  OA22X1 U4964 ( .IN1(n30006), .IN2(n449), .IN3(n30014), .IN4(n492), .Q(n5013)
         );
  OA221X1 U4965 ( .IN1(n29958), .IN2(n535), .IN3(n29966), .IN4(n578), .IN5(
        n5014), .Q(n5007) );
  OA22X1 U4966 ( .IN1(n29974), .IN2(n621), .IN3(n29982), .IN4(n664), .Q(n5014)
         );
  NAND4X0 U4967 ( .IN1(n5015), .IN2(n5016), .IN3(n5017), .IN4(n5018), .QN(
        n4995) );
  OA221X1 U4968 ( .IN1(n29926), .IN2(n19), .IN3(n29934), .IN4(n62), .IN5(n5019), .Q(n5018) );
  OA22X1 U4969 ( .IN1(n29942), .IN2(n105), .IN3(n29950), .IN4(n148), .Q(n5019)
         );
  OA221X1 U4970 ( .IN1(n29894), .IN2(n191), .IN3(n29902), .IN4(n234), .IN5(
        n5020), .Q(n5017) );
  OA22X1 U4971 ( .IN1(n29910), .IN2(n277), .IN3(n29918), .IN4(n320), .Q(n5020)
         );
  OA221X1 U4972 ( .IN1(n29862), .IN2(n363), .IN3(n29870), .IN4(n406), .IN5(
        n5021), .Q(n5016) );
  OA22X1 U4973 ( .IN1(n29878), .IN2(n449), .IN3(n29886), .IN4(n492), .Q(n5021)
         );
  OA221X1 U4974 ( .IN1(n29830), .IN2(n535), .IN3(n29838), .IN4(n578), .IN5(
        n5022), .Q(n5015) );
  OA22X1 U4975 ( .IN1(n29846), .IN2(n621), .IN3(n29854), .IN4(n664), .Q(n5022)
         );
  NAND4X0 U4976 ( .IN1(n5023), .IN2(n5024), .IN3(n5025), .IN4(n5026), .QN(
        n4994) );
  OA221X1 U4977 ( .IN1(n29798), .IN2(n19), .IN3(n29806), .IN4(n62), .IN5(n5027), .Q(n5026) );
  OA22X1 U4978 ( .IN1(n29814), .IN2(n105), .IN3(n29822), .IN4(n148), .Q(n5027)
         );
  OA221X1 U4979 ( .IN1(n29766), .IN2(n191), .IN3(n29774), .IN4(n234), .IN5(
        n5028), .Q(n5025) );
  OA22X1 U4980 ( .IN1(n29782), .IN2(n277), .IN3(n29790), .IN4(n320), .Q(n5028)
         );
  OA221X1 U4981 ( .IN1(n29734), .IN2(n363), .IN3(n29742), .IN4(n406), .IN5(
        n5029), .Q(n5024) );
  OA22X1 U4982 ( .IN1(n29750), .IN2(n449), .IN3(n29758), .IN4(n492), .Q(n5029)
         );
  OA221X1 U4983 ( .IN1(n29702), .IN2(n535), .IN3(n29710), .IN4(n578), .IN5(
        n5030), .Q(n5023) );
  OA22X1 U4984 ( .IN1(n29718), .IN2(n621), .IN3(n29726), .IN4(n664), .Q(n5030)
         );
  AO221X1 U4985 ( .IN1(n2287), .IN2(n5031), .IN3(n2289), .IN4(n5032), .IN5(
        n5033), .Q(n4954) );
  AO22X1 U4986 ( .IN1(n2292), .IN2(n5034), .IN3(n2294), .IN4(n5035), .Q(n5033)
         );
  NAND4X0 U4987 ( .IN1(n5036), .IN2(n5037), .IN3(n5038), .IN4(n5039), .QN(
        n5035) );
  OA221X1 U4988 ( .IN1(n31718), .IN2(n18), .IN3(n31726), .IN4(n61), .IN5(n5040), .Q(n5039) );
  OA22X1 U4989 ( .IN1(n31734), .IN2(n104), .IN3(n31742), .IN4(n147), .Q(n5040)
         );
  OA221X1 U4990 ( .IN1(n31686), .IN2(n190), .IN3(n31694), .IN4(n233), .IN5(
        n5041), .Q(n5038) );
  OA22X1 U4991 ( .IN1(n31702), .IN2(n276), .IN3(n31710), .IN4(n319), .Q(n5041)
         );
  OA221X1 U4992 ( .IN1(n31654), .IN2(n362), .IN3(n31662), .IN4(n405), .IN5(
        n5042), .Q(n5037) );
  OA22X1 U4993 ( .IN1(n31670), .IN2(n448), .IN3(n31678), .IN4(n491), .Q(n5042)
         );
  OA221X1 U4994 ( .IN1(n31622), .IN2(n534), .IN3(n31630), .IN4(n577), .IN5(
        n5043), .Q(n5036) );
  OA22X1 U4995 ( .IN1(n31638), .IN2(n620), .IN3(n31646), .IN4(n663), .Q(n5043)
         );
  NAND4X0 U4996 ( .IN1(n5044), .IN2(n5045), .IN3(n5046), .IN4(n5047), .QN(
        n5034) );
  OA221X1 U4997 ( .IN1(n31590), .IN2(n18), .IN3(n31598), .IN4(n61), .IN5(n5048), .Q(n5047) );
  OA22X1 U4998 ( .IN1(n31606), .IN2(n104), .IN3(n31614), .IN4(n147), .Q(n5048)
         );
  OA221X1 U4999 ( .IN1(n31558), .IN2(n190), .IN3(n31566), .IN4(n233), .IN5(
        n5049), .Q(n5046) );
  OA22X1 U5000 ( .IN1(n31574), .IN2(n276), .IN3(n31582), .IN4(n319), .Q(n5049)
         );
  OA221X1 U5001 ( .IN1(n31526), .IN2(n362), .IN3(n31534), .IN4(n405), .IN5(
        n5050), .Q(n5045) );
  OA22X1 U5002 ( .IN1(n31542), .IN2(n448), .IN3(n31550), .IN4(n491), .Q(n5050)
         );
  OA221X1 U5003 ( .IN1(n31494), .IN2(n534), .IN3(n31502), .IN4(n577), .IN5(
        n5051), .Q(n5044) );
  OA22X1 U5004 ( .IN1(n31510), .IN2(n620), .IN3(n31518), .IN4(n663), .Q(n5051)
         );
  NAND4X0 U5005 ( .IN1(n5052), .IN2(n5053), .IN3(n5054), .IN4(n5055), .QN(
        n5032) );
  OA221X1 U5006 ( .IN1(n31462), .IN2(n18), .IN3(n31470), .IN4(n61), .IN5(n5056), .Q(n5055) );
  OA22X1 U5007 ( .IN1(n31478), .IN2(n104), .IN3(n31486), .IN4(n147), .Q(n5056)
         );
  OA221X1 U5008 ( .IN1(n31430), .IN2(n190), .IN3(n31438), .IN4(n233), .IN5(
        n5057), .Q(n5054) );
  OA22X1 U5009 ( .IN1(n31446), .IN2(n276), .IN3(n31454), .IN4(n319), .Q(n5057)
         );
  OA221X1 U5010 ( .IN1(n31398), .IN2(n362), .IN3(n31406), .IN4(n405), .IN5(
        n5058), .Q(n5053) );
  OA22X1 U5011 ( .IN1(n31414), .IN2(n448), .IN3(n31422), .IN4(n491), .Q(n5058)
         );
  OA221X1 U5012 ( .IN1(n31366), .IN2(n534), .IN3(n31374), .IN4(n577), .IN5(
        n5059), .Q(n5052) );
  OA22X1 U5013 ( .IN1(n31382), .IN2(n620), .IN3(n31390), .IN4(n663), .Q(n5059)
         );
  NAND4X0 U5014 ( .IN1(n5060), .IN2(n5061), .IN3(n5062), .IN4(n5063), .QN(
        n5031) );
  OA221X1 U5015 ( .IN1(n31334), .IN2(n18), .IN3(n31342), .IN4(n61), .IN5(n5064), .Q(n5063) );
  OA22X1 U5016 ( .IN1(n31350), .IN2(n104), .IN3(n31358), .IN4(n147), .Q(n5064)
         );
  OA221X1 U5017 ( .IN1(n31302), .IN2(n190), .IN3(n31310), .IN4(n233), .IN5(
        n5065), .Q(n5062) );
  OA22X1 U5018 ( .IN1(n31318), .IN2(n276), .IN3(n31326), .IN4(n319), .Q(n5065)
         );
  OA221X1 U5019 ( .IN1(n31270), .IN2(n362), .IN3(n31278), .IN4(n405), .IN5(
        n5066), .Q(n5061) );
  OA22X1 U5020 ( .IN1(n31286), .IN2(n448), .IN3(n31294), .IN4(n491), .Q(n5066)
         );
  OA221X1 U5021 ( .IN1(n31238), .IN2(n534), .IN3(n31246), .IN4(n577), .IN5(
        n5067), .Q(n5060) );
  OA22X1 U5022 ( .IN1(n31254), .IN2(n620), .IN3(n31262), .IN4(n663), .Q(n5067)
         );
  AO221X1 U5023 ( .IN1(n2328), .IN2(n5068), .IN3(n2330), .IN4(n5069), .IN5(
        n5070), .Q(n4953) );
  AO22X1 U5024 ( .IN1(n2333), .IN2(n5071), .IN3(n2335), .IN4(n5072), .Q(n5070)
         );
  NAND4X0 U5025 ( .IN1(n5073), .IN2(n5074), .IN3(n5075), .IN4(n5076), .QN(
        n5072) );
  OA221X1 U5026 ( .IN1(n31206), .IN2(n18), .IN3(n31214), .IN4(n61), .IN5(n5077), .Q(n5076) );
  OA22X1 U5027 ( .IN1(n31222), .IN2(n104), .IN3(n31230), .IN4(n147), .Q(n5077)
         );
  OA221X1 U5028 ( .IN1(n31174), .IN2(n190), .IN3(n31182), .IN4(n233), .IN5(
        n5078), .Q(n5075) );
  OA22X1 U5029 ( .IN1(n31190), .IN2(n276), .IN3(n31198), .IN4(n319), .Q(n5078)
         );
  OA221X1 U5030 ( .IN1(n31142), .IN2(n362), .IN3(n31150), .IN4(n405), .IN5(
        n5079), .Q(n5074) );
  OA22X1 U5031 ( .IN1(n31158), .IN2(n448), .IN3(n31166), .IN4(n491), .Q(n5079)
         );
  OA221X1 U5032 ( .IN1(n31110), .IN2(n534), .IN3(n31118), .IN4(n577), .IN5(
        n5080), .Q(n5073) );
  OA22X1 U5033 ( .IN1(n31126), .IN2(n620), .IN3(n31134), .IN4(n663), .Q(n5080)
         );
  NAND4X0 U5034 ( .IN1(n5081), .IN2(n5082), .IN3(n5083), .IN4(n5084), .QN(
        n5071) );
  OA221X1 U5035 ( .IN1(n31078), .IN2(n18), .IN3(n31086), .IN4(n61), .IN5(n5085), .Q(n5084) );
  OA22X1 U5036 ( .IN1(n31094), .IN2(n104), .IN3(n31102), .IN4(n147), .Q(n5085)
         );
  OA221X1 U5037 ( .IN1(n31046), .IN2(n190), .IN3(n31054), .IN4(n233), .IN5(
        n5086), .Q(n5083) );
  OA22X1 U5038 ( .IN1(n31062), .IN2(n276), .IN3(n31070), .IN4(n319), .Q(n5086)
         );
  OA221X1 U5039 ( .IN1(n31014), .IN2(n362), .IN3(n31022), .IN4(n405), .IN5(
        n5087), .Q(n5082) );
  OA22X1 U5040 ( .IN1(n31030), .IN2(n448), .IN3(n31038), .IN4(n491), .Q(n5087)
         );
  OA221X1 U5041 ( .IN1(n30982), .IN2(n534), .IN3(n30990), .IN4(n577), .IN5(
        n5088), .Q(n5081) );
  OA22X1 U5042 ( .IN1(n30998), .IN2(n620), .IN3(n31006), .IN4(n663), .Q(n5088)
         );
  NAND4X0 U5043 ( .IN1(n5089), .IN2(n5090), .IN3(n5091), .IN4(n5092), .QN(
        n5069) );
  OA221X1 U5044 ( .IN1(n30950), .IN2(n18), .IN3(n30958), .IN4(n61), .IN5(n5093), .Q(n5092) );
  OA22X1 U5045 ( .IN1(n30966), .IN2(n104), .IN3(n30974), .IN4(n147), .Q(n5093)
         );
  OA221X1 U5046 ( .IN1(n30918), .IN2(n190), .IN3(n30926), .IN4(n233), .IN5(
        n5094), .Q(n5091) );
  OA22X1 U5047 ( .IN1(n30934), .IN2(n276), .IN3(n30942), .IN4(n319), .Q(n5094)
         );
  OA221X1 U5048 ( .IN1(n30886), .IN2(n362), .IN3(n30894), .IN4(n405), .IN5(
        n5095), .Q(n5090) );
  OA22X1 U5049 ( .IN1(n30902), .IN2(n448), .IN3(n30910), .IN4(n491), .Q(n5095)
         );
  OA221X1 U5050 ( .IN1(n30854), .IN2(n534), .IN3(n30862), .IN4(n577), .IN5(
        n5096), .Q(n5089) );
  OA22X1 U5051 ( .IN1(n30870), .IN2(n620), .IN3(n30878), .IN4(n663), .Q(n5096)
         );
  NAND4X0 U5052 ( .IN1(n5097), .IN2(n5098), .IN3(n5099), .IN4(n5100), .QN(
        n5068) );
  OA221X1 U5053 ( .IN1(n30822), .IN2(n18), .IN3(n30830), .IN4(n61), .IN5(n5101), .Q(n5100) );
  OA22X1 U5054 ( .IN1(n30838), .IN2(n104), .IN3(n30846), .IN4(n147), .Q(n5101)
         );
  OA221X1 U5055 ( .IN1(n30790), .IN2(n190), .IN3(n30798), .IN4(n233), .IN5(
        n5102), .Q(n5099) );
  OA22X1 U5056 ( .IN1(n30806), .IN2(n276), .IN3(n30814), .IN4(n319), .Q(n5102)
         );
  OA221X1 U5057 ( .IN1(n30758), .IN2(n362), .IN3(n30766), .IN4(n405), .IN5(
        n5103), .Q(n5098) );
  OA22X1 U5058 ( .IN1(n30774), .IN2(n448), .IN3(n30782), .IN4(n491), .Q(n5103)
         );
  OA221X1 U5059 ( .IN1(n30726), .IN2(n534), .IN3(n30734), .IN4(n577), .IN5(
        n5104), .Q(n5097) );
  OA22X1 U5060 ( .IN1(n30742), .IN2(n620), .IN3(n30750), .IN4(n663), .Q(n5104)
         );
  OR4X1 U5061 ( .IN1(n5105), .IN2(n5106), .IN3(n5107), .IN4(n5108), .Q(n2183)
         );
  AO221X1 U5062 ( .IN1(n2157), .IN2(n5109), .IN3(n2159), .IN4(n5110), .IN5(
        n5111), .Q(n5108) );
  AO22X1 U5063 ( .IN1(n2162), .IN2(n5112), .IN3(n2164), .IN4(n5113), .Q(n5111)
         );
  NAND4X0 U5064 ( .IN1(n5114), .IN2(n5115), .IN3(n5116), .IN4(n5117), .QN(
        n5113) );
  OA221X1 U5065 ( .IN1(n30693), .IN2(n18), .IN3(n30701), .IN4(n61), .IN5(n5118), .Q(n5117) );
  OA22X1 U5066 ( .IN1(n30709), .IN2(n104), .IN3(n30717), .IN4(n147), .Q(n5118)
         );
  OA221X1 U5067 ( .IN1(n30661), .IN2(n190), .IN3(n30669), .IN4(n233), .IN5(
        n5119), .Q(n5116) );
  OA22X1 U5068 ( .IN1(n30677), .IN2(n276), .IN3(n30685), .IN4(n319), .Q(n5119)
         );
  OA221X1 U5069 ( .IN1(n30629), .IN2(n362), .IN3(n30637), .IN4(n405), .IN5(
        n5120), .Q(n5115) );
  OA22X1 U5070 ( .IN1(n30645), .IN2(n448), .IN3(n30653), .IN4(n491), .Q(n5120)
         );
  OA221X1 U5071 ( .IN1(n30597), .IN2(n534), .IN3(n30605), .IN4(n577), .IN5(
        n5121), .Q(n5114) );
  OA22X1 U5072 ( .IN1(n30613), .IN2(n620), .IN3(n30621), .IN4(n663), .Q(n5121)
         );
  NAND4X0 U5073 ( .IN1(n5122), .IN2(n5123), .IN3(n5124), .IN4(n5125), .QN(
        n5112) );
  OA221X1 U5074 ( .IN1(n30565), .IN2(n18), .IN3(n30573), .IN4(n61), .IN5(n5126), .Q(n5125) );
  OA22X1 U5075 ( .IN1(n30581), .IN2(n104), .IN3(n30589), .IN4(n147), .Q(n5126)
         );
  OA221X1 U5076 ( .IN1(n30533), .IN2(n190), .IN3(n30541), .IN4(n233), .IN5(
        n5127), .Q(n5124) );
  OA22X1 U5077 ( .IN1(n30549), .IN2(n276), .IN3(n30557), .IN4(n319), .Q(n5127)
         );
  OA221X1 U5078 ( .IN1(n30501), .IN2(n362), .IN3(n30509), .IN4(n405), .IN5(
        n5128), .Q(n5123) );
  OA22X1 U5079 ( .IN1(n30517), .IN2(n448), .IN3(n30525), .IN4(n491), .Q(n5128)
         );
  OA221X1 U5080 ( .IN1(n30469), .IN2(n534), .IN3(n30477), .IN4(n577), .IN5(
        n5129), .Q(n5122) );
  OA22X1 U5081 ( .IN1(n30485), .IN2(n620), .IN3(n30493), .IN4(n663), .Q(n5129)
         );
  NAND4X0 U5082 ( .IN1(n5130), .IN2(n5131), .IN3(n5132), .IN4(n5133), .QN(
        n5110) );
  OA221X1 U5083 ( .IN1(n30437), .IN2(n18), .IN3(n30445), .IN4(n61), .IN5(n5134), .Q(n5133) );
  OA22X1 U5084 ( .IN1(n30453), .IN2(n104), .IN3(n30461), .IN4(n147), .Q(n5134)
         );
  OA221X1 U5085 ( .IN1(n30405), .IN2(n190), .IN3(n30413), .IN4(n233), .IN5(
        n5135), .Q(n5132) );
  OA22X1 U5086 ( .IN1(n30421), .IN2(n276), .IN3(n30429), .IN4(n319), .Q(n5135)
         );
  OA221X1 U5087 ( .IN1(n30373), .IN2(n362), .IN3(n30381), .IN4(n405), .IN5(
        n5136), .Q(n5131) );
  OA22X1 U5088 ( .IN1(n30389), .IN2(n448), .IN3(n30397), .IN4(n491), .Q(n5136)
         );
  OA221X1 U5089 ( .IN1(n30341), .IN2(n534), .IN3(n30349), .IN4(n577), .IN5(
        n5137), .Q(n5130) );
  OA22X1 U5090 ( .IN1(n30357), .IN2(n620), .IN3(n30365), .IN4(n663), .Q(n5137)
         );
  NAND4X0 U5091 ( .IN1(n5138), .IN2(n5139), .IN3(n5140), .IN4(n5141), .QN(
        n5109) );
  OA221X1 U5092 ( .IN1(n30309), .IN2(n18), .IN3(n30317), .IN4(n61), .IN5(n5142), .Q(n5141) );
  OA22X1 U5093 ( .IN1(n30325), .IN2(n104), .IN3(n30333), .IN4(n147), .Q(n5142)
         );
  OA221X1 U5094 ( .IN1(n30277), .IN2(n190), .IN3(n30285), .IN4(n233), .IN5(
        n5143), .Q(n5140) );
  OA22X1 U5095 ( .IN1(n30293), .IN2(n276), .IN3(n30301), .IN4(n319), .Q(n5143)
         );
  OA221X1 U5096 ( .IN1(n30245), .IN2(n362), .IN3(n30253), .IN4(n405), .IN5(
        n5144), .Q(n5139) );
  OA22X1 U5097 ( .IN1(n30261), .IN2(n448), .IN3(n30269), .IN4(n491), .Q(n5144)
         );
  OA221X1 U5098 ( .IN1(n30213), .IN2(n534), .IN3(n30221), .IN4(n577), .IN5(
        n5145), .Q(n5138) );
  OA22X1 U5099 ( .IN1(n30229), .IN2(n620), .IN3(n30237), .IN4(n663), .Q(n5145)
         );
  AO221X1 U5100 ( .IN1(n2246), .IN2(n5146), .IN3(n2248), .IN4(n5147), .IN5(
        n5148), .Q(n5107) );
  AO22X1 U5101 ( .IN1(n2251), .IN2(n5149), .IN3(n2253), .IN4(n5150), .Q(n5148)
         );
  NAND4X0 U5102 ( .IN1(n5151), .IN2(n5152), .IN3(n5153), .IN4(n5154), .QN(
        n5150) );
  OA221X1 U5103 ( .IN1(n30181), .IN2(n17), .IN3(n30189), .IN4(n60), .IN5(n5155), .Q(n5154) );
  OA22X1 U5104 ( .IN1(n30197), .IN2(n103), .IN3(n30205), .IN4(n146), .Q(n5155)
         );
  OA221X1 U5105 ( .IN1(n30149), .IN2(n189), .IN3(n30157), .IN4(n232), .IN5(
        n5156), .Q(n5153) );
  OA22X1 U5106 ( .IN1(n30165), .IN2(n275), .IN3(n30173), .IN4(n318), .Q(n5156)
         );
  OA221X1 U5107 ( .IN1(n30117), .IN2(n361), .IN3(n30125), .IN4(n404), .IN5(
        n5157), .Q(n5152) );
  OA22X1 U5108 ( .IN1(n30133), .IN2(n447), .IN3(n30141), .IN4(n490), .Q(n5157)
         );
  OA221X1 U5109 ( .IN1(n30085), .IN2(n533), .IN3(n30093), .IN4(n576), .IN5(
        n5158), .Q(n5151) );
  OA22X1 U5110 ( .IN1(n30101), .IN2(n619), .IN3(n30109), .IN4(n662), .Q(n5158)
         );
  NAND4X0 U5111 ( .IN1(n5159), .IN2(n5160), .IN3(n5161), .IN4(n5162), .QN(
        n5149) );
  OA221X1 U5112 ( .IN1(n30053), .IN2(n17), .IN3(n30061), .IN4(n60), .IN5(n5163), .Q(n5162) );
  OA22X1 U5113 ( .IN1(n30069), .IN2(n103), .IN3(n30077), .IN4(n146), .Q(n5163)
         );
  OA221X1 U5114 ( .IN1(n30021), .IN2(n189), .IN3(n30029), .IN4(n232), .IN5(
        n5164), .Q(n5161) );
  OA22X1 U5115 ( .IN1(n30037), .IN2(n275), .IN3(n30045), .IN4(n318), .Q(n5164)
         );
  OA221X1 U5116 ( .IN1(n29989), .IN2(n361), .IN3(n29997), .IN4(n404), .IN5(
        n5165), .Q(n5160) );
  OA22X1 U5117 ( .IN1(n30005), .IN2(n447), .IN3(n30013), .IN4(n490), .Q(n5165)
         );
  OA221X1 U5118 ( .IN1(n29957), .IN2(n533), .IN3(n29965), .IN4(n576), .IN5(
        n5166), .Q(n5159) );
  OA22X1 U5119 ( .IN1(n29973), .IN2(n619), .IN3(n29981), .IN4(n662), .Q(n5166)
         );
  NAND4X0 U5120 ( .IN1(n5167), .IN2(n5168), .IN3(n5169), .IN4(n5170), .QN(
        n5147) );
  OA221X1 U5121 ( .IN1(n29925), .IN2(n17), .IN3(n29933), .IN4(n60), .IN5(n5171), .Q(n5170) );
  OA22X1 U5122 ( .IN1(n29941), .IN2(n103), .IN3(n29949), .IN4(n146), .Q(n5171)
         );
  OA221X1 U5123 ( .IN1(n29893), .IN2(n189), .IN3(n29901), .IN4(n232), .IN5(
        n5172), .Q(n5169) );
  OA22X1 U5124 ( .IN1(n29909), .IN2(n275), .IN3(n29917), .IN4(n318), .Q(n5172)
         );
  OA221X1 U5125 ( .IN1(n29861), .IN2(n361), .IN3(n29869), .IN4(n404), .IN5(
        n5173), .Q(n5168) );
  OA22X1 U5126 ( .IN1(n29877), .IN2(n447), .IN3(n29885), .IN4(n490), .Q(n5173)
         );
  OA221X1 U5127 ( .IN1(n29829), .IN2(n533), .IN3(n29837), .IN4(n576), .IN5(
        n5174), .Q(n5167) );
  OA22X1 U5128 ( .IN1(n29845), .IN2(n619), .IN3(n29853), .IN4(n662), .Q(n5174)
         );
  NAND4X0 U5129 ( .IN1(n5175), .IN2(n5176), .IN3(n5177), .IN4(n5178), .QN(
        n5146) );
  OA221X1 U5130 ( .IN1(n29797), .IN2(n17), .IN3(n29805), .IN4(n60), .IN5(n5179), .Q(n5178) );
  OA22X1 U5131 ( .IN1(n29813), .IN2(n103), .IN3(n29821), .IN4(n146), .Q(n5179)
         );
  OA221X1 U5132 ( .IN1(n29765), .IN2(n189), .IN3(n29773), .IN4(n232), .IN5(
        n5180), .Q(n5177) );
  OA22X1 U5133 ( .IN1(n29781), .IN2(n275), .IN3(n29789), .IN4(n318), .Q(n5180)
         );
  OA221X1 U5134 ( .IN1(n29733), .IN2(n361), .IN3(n29741), .IN4(n404), .IN5(
        n5181), .Q(n5176) );
  OA22X1 U5135 ( .IN1(n29749), .IN2(n447), .IN3(n29757), .IN4(n490), .Q(n5181)
         );
  OA221X1 U5136 ( .IN1(n29701), .IN2(n533), .IN3(n29709), .IN4(n576), .IN5(
        n5182), .Q(n5175) );
  OA22X1 U5137 ( .IN1(n29717), .IN2(n619), .IN3(n29725), .IN4(n662), .Q(n5182)
         );
  AO221X1 U5138 ( .IN1(n2287), .IN2(n5183), .IN3(n2289), .IN4(n5184), .IN5(
        n5185), .Q(n5106) );
  AO22X1 U5139 ( .IN1(n2292), .IN2(n5186), .IN3(n2294), .IN4(n5187), .Q(n5185)
         );
  NAND4X0 U5140 ( .IN1(n5188), .IN2(n5189), .IN3(n5190), .IN4(n5191), .QN(
        n5187) );
  OA221X1 U5141 ( .IN1(n31717), .IN2(n17), .IN3(n31725), .IN4(n60), .IN5(n5192), .Q(n5191) );
  OA22X1 U5142 ( .IN1(n31733), .IN2(n103), .IN3(n31741), .IN4(n146), .Q(n5192)
         );
  OA221X1 U5143 ( .IN1(n31685), .IN2(n189), .IN3(n31693), .IN4(n232), .IN5(
        n5193), .Q(n5190) );
  OA22X1 U5144 ( .IN1(n31701), .IN2(n275), .IN3(n31709), .IN4(n318), .Q(n5193)
         );
  OA221X1 U5145 ( .IN1(n31653), .IN2(n361), .IN3(n31661), .IN4(n404), .IN5(
        n5194), .Q(n5189) );
  OA22X1 U5146 ( .IN1(n31669), .IN2(n447), .IN3(n31677), .IN4(n490), .Q(n5194)
         );
  OA221X1 U5147 ( .IN1(n31621), .IN2(n533), .IN3(n31629), .IN4(n576), .IN5(
        n5195), .Q(n5188) );
  OA22X1 U5148 ( .IN1(n31637), .IN2(n619), .IN3(n31645), .IN4(n662), .Q(n5195)
         );
  NAND4X0 U5149 ( .IN1(n5196), .IN2(n5197), .IN3(n5198), .IN4(n5199), .QN(
        n5186) );
  OA221X1 U5150 ( .IN1(n31589), .IN2(n17), .IN3(n31597), .IN4(n60), .IN5(n5200), .Q(n5199) );
  OA22X1 U5151 ( .IN1(n31605), .IN2(n103), .IN3(n31613), .IN4(n146), .Q(n5200)
         );
  OA221X1 U5152 ( .IN1(n31557), .IN2(n189), .IN3(n31565), .IN4(n232), .IN5(
        n5201), .Q(n5198) );
  OA22X1 U5153 ( .IN1(n31573), .IN2(n275), .IN3(n31581), .IN4(n318), .Q(n5201)
         );
  OA221X1 U5154 ( .IN1(n31525), .IN2(n361), .IN3(n31533), .IN4(n404), .IN5(
        n5202), .Q(n5197) );
  OA22X1 U5155 ( .IN1(n31541), .IN2(n447), .IN3(n31549), .IN4(n490), .Q(n5202)
         );
  OA221X1 U5156 ( .IN1(n31493), .IN2(n533), .IN3(n31501), .IN4(n576), .IN5(
        n5203), .Q(n5196) );
  OA22X1 U5157 ( .IN1(n31509), .IN2(n619), .IN3(n31517), .IN4(n662), .Q(n5203)
         );
  NAND4X0 U5158 ( .IN1(n5204), .IN2(n5205), .IN3(n5206), .IN4(n5207), .QN(
        n5184) );
  OA221X1 U5159 ( .IN1(n31461), .IN2(n17), .IN3(n31469), .IN4(n60), .IN5(n5208), .Q(n5207) );
  OA22X1 U5160 ( .IN1(n31477), .IN2(n103), .IN3(n31485), .IN4(n146), .Q(n5208)
         );
  OA221X1 U5161 ( .IN1(n31429), .IN2(n189), .IN3(n31437), .IN4(n232), .IN5(
        n5209), .Q(n5206) );
  OA22X1 U5162 ( .IN1(n31445), .IN2(n275), .IN3(n31453), .IN4(n318), .Q(n5209)
         );
  OA221X1 U5163 ( .IN1(n31397), .IN2(n361), .IN3(n31405), .IN4(n404), .IN5(
        n5210), .Q(n5205) );
  OA22X1 U5164 ( .IN1(n31413), .IN2(n447), .IN3(n31421), .IN4(n490), .Q(n5210)
         );
  OA221X1 U5165 ( .IN1(n31365), .IN2(n533), .IN3(n31373), .IN4(n576), .IN5(
        n5211), .Q(n5204) );
  OA22X1 U5166 ( .IN1(n31381), .IN2(n619), .IN3(n31389), .IN4(n662), .Q(n5211)
         );
  NAND4X0 U5167 ( .IN1(n5212), .IN2(n5213), .IN3(n5214), .IN4(n5215), .QN(
        n5183) );
  OA221X1 U5168 ( .IN1(n31333), .IN2(n17), .IN3(n31341), .IN4(n60), .IN5(n5216), .Q(n5215) );
  OA22X1 U5169 ( .IN1(n31349), .IN2(n103), .IN3(n31357), .IN4(n146), .Q(n5216)
         );
  OA221X1 U5170 ( .IN1(n31301), .IN2(n189), .IN3(n31309), .IN4(n232), .IN5(
        n5217), .Q(n5214) );
  OA22X1 U5171 ( .IN1(n31317), .IN2(n275), .IN3(n31325), .IN4(n318), .Q(n5217)
         );
  OA221X1 U5172 ( .IN1(n31269), .IN2(n361), .IN3(n31277), .IN4(n404), .IN5(
        n5218), .Q(n5213) );
  OA22X1 U5173 ( .IN1(n31285), .IN2(n447), .IN3(n31293), .IN4(n490), .Q(n5218)
         );
  OA221X1 U5174 ( .IN1(n31237), .IN2(n533), .IN3(n31245), .IN4(n576), .IN5(
        n5219), .Q(n5212) );
  OA22X1 U5175 ( .IN1(n31253), .IN2(n619), .IN3(n31261), .IN4(n662), .Q(n5219)
         );
  AO221X1 U5176 ( .IN1(n2328), .IN2(n5220), .IN3(n2330), .IN4(n5221), .IN5(
        n5222), .Q(n5105) );
  AO22X1 U5177 ( .IN1(n2333), .IN2(n5223), .IN3(n2335), .IN4(n5224), .Q(n5222)
         );
  NAND4X0 U5178 ( .IN1(n5225), .IN2(n5226), .IN3(n5227), .IN4(n5228), .QN(
        n5224) );
  OA221X1 U5179 ( .IN1(n31205), .IN2(n17), .IN3(n31213), .IN4(n60), .IN5(n5229), .Q(n5228) );
  OA22X1 U5180 ( .IN1(n31221), .IN2(n103), .IN3(n31229), .IN4(n146), .Q(n5229)
         );
  OA221X1 U5181 ( .IN1(n31173), .IN2(n189), .IN3(n31181), .IN4(n232), .IN5(
        n5230), .Q(n5227) );
  OA22X1 U5182 ( .IN1(n31189), .IN2(n275), .IN3(n31197), .IN4(n318), .Q(n5230)
         );
  OA221X1 U5183 ( .IN1(n31141), .IN2(n361), .IN3(n31149), .IN4(n404), .IN5(
        n5231), .Q(n5226) );
  OA22X1 U5184 ( .IN1(n31157), .IN2(n447), .IN3(n31165), .IN4(n490), .Q(n5231)
         );
  OA221X1 U5185 ( .IN1(n31109), .IN2(n533), .IN3(n31117), .IN4(n576), .IN5(
        n5232), .Q(n5225) );
  OA22X1 U5186 ( .IN1(n31125), .IN2(n619), .IN3(n31133), .IN4(n662), .Q(n5232)
         );
  NAND4X0 U5187 ( .IN1(n5233), .IN2(n5234), .IN3(n5235), .IN4(n5236), .QN(
        n5223) );
  OA221X1 U5188 ( .IN1(n31077), .IN2(n17), .IN3(n31085), .IN4(n60), .IN5(n5237), .Q(n5236) );
  OA22X1 U5189 ( .IN1(n31093), .IN2(n103), .IN3(n31101), .IN4(n146), .Q(n5237)
         );
  OA221X1 U5190 ( .IN1(n31045), .IN2(n189), .IN3(n31053), .IN4(n232), .IN5(
        n5238), .Q(n5235) );
  OA22X1 U5191 ( .IN1(n31061), .IN2(n275), .IN3(n31069), .IN4(n318), .Q(n5238)
         );
  OA221X1 U5192 ( .IN1(n31013), .IN2(n361), .IN3(n31021), .IN4(n404), .IN5(
        n5239), .Q(n5234) );
  OA22X1 U5193 ( .IN1(n31029), .IN2(n447), .IN3(n31037), .IN4(n490), .Q(n5239)
         );
  OA221X1 U5194 ( .IN1(n30981), .IN2(n533), .IN3(n30989), .IN4(n576), .IN5(
        n5240), .Q(n5233) );
  OA22X1 U5195 ( .IN1(n30997), .IN2(n619), .IN3(n31005), .IN4(n662), .Q(n5240)
         );
  NAND4X0 U5196 ( .IN1(n5241), .IN2(n5242), .IN3(n5243), .IN4(n5244), .QN(
        n5221) );
  OA221X1 U5197 ( .IN1(n30949), .IN2(n17), .IN3(n30957), .IN4(n60), .IN5(n5245), .Q(n5244) );
  OA22X1 U5198 ( .IN1(n30965), .IN2(n103), .IN3(n30973), .IN4(n146), .Q(n5245)
         );
  OA221X1 U5199 ( .IN1(n30917), .IN2(n189), .IN3(n30925), .IN4(n232), .IN5(
        n5246), .Q(n5243) );
  OA22X1 U5200 ( .IN1(n30933), .IN2(n275), .IN3(n30941), .IN4(n318), .Q(n5246)
         );
  OA221X1 U5201 ( .IN1(n30885), .IN2(n361), .IN3(n30893), .IN4(n404), .IN5(
        n5247), .Q(n5242) );
  OA22X1 U5202 ( .IN1(n30901), .IN2(n447), .IN3(n30909), .IN4(n490), .Q(n5247)
         );
  OA221X1 U5203 ( .IN1(n30853), .IN2(n533), .IN3(n30861), .IN4(n576), .IN5(
        n5248), .Q(n5241) );
  OA22X1 U5204 ( .IN1(n30869), .IN2(n619), .IN3(n30877), .IN4(n662), .Q(n5248)
         );
  NAND4X0 U5205 ( .IN1(n5249), .IN2(n5250), .IN3(n5251), .IN4(n5252), .QN(
        n5220) );
  OA221X1 U5206 ( .IN1(n30821), .IN2(n17), .IN3(n30829), .IN4(n60), .IN5(n5253), .Q(n5252) );
  OA22X1 U5207 ( .IN1(n30837), .IN2(n103), .IN3(n30845), .IN4(n146), .Q(n5253)
         );
  OA221X1 U5208 ( .IN1(n30789), .IN2(n189), .IN3(n30797), .IN4(n232), .IN5(
        n5254), .Q(n5251) );
  OA22X1 U5209 ( .IN1(n30805), .IN2(n275), .IN3(n30813), .IN4(n318), .Q(n5254)
         );
  OA221X1 U5210 ( .IN1(n30757), .IN2(n361), .IN3(n30765), .IN4(n404), .IN5(
        n5255), .Q(n5250) );
  OA22X1 U5211 ( .IN1(n30773), .IN2(n447), .IN3(n30781), .IN4(n490), .Q(n5255)
         );
  OA221X1 U5212 ( .IN1(n30725), .IN2(n533), .IN3(n30733), .IN4(n576), .IN5(
        n5256), .Q(n5249) );
  OA22X1 U5213 ( .IN1(n30741), .IN2(n619), .IN3(n30749), .IN4(n662), .Q(n5256)
         );
  OR4X1 U5214 ( .IN1(n5257), .IN2(n5258), .IN3(n5259), .IN4(n5260), .Q(n2182)
         );
  AO221X1 U5215 ( .IN1(n2157), .IN2(n5261), .IN3(n2159), .IN4(n5262), .IN5(
        n5263), .Q(n5260) );
  AO22X1 U5216 ( .IN1(n2162), .IN2(n5264), .IN3(n2164), .IN4(n5265), .Q(n5263)
         );
  NAND4X0 U5217 ( .IN1(n5266), .IN2(n5267), .IN3(n5268), .IN4(n5269), .QN(
        n5265) );
  OA221X1 U5218 ( .IN1(n30692), .IN2(n16), .IN3(n30700), .IN4(n59), .IN5(n5270), .Q(n5269) );
  OA22X1 U5219 ( .IN1(n30708), .IN2(n102), .IN3(n30716), .IN4(n145), .Q(n5270)
         );
  OA221X1 U5220 ( .IN1(n30660), .IN2(n188), .IN3(n30668), .IN4(n231), .IN5(
        n5271), .Q(n5268) );
  OA22X1 U5221 ( .IN1(n30676), .IN2(n274), .IN3(n30684), .IN4(n317), .Q(n5271)
         );
  OA221X1 U5222 ( .IN1(n30628), .IN2(n360), .IN3(n30636), .IN4(n403), .IN5(
        n5272), .Q(n5267) );
  OA22X1 U5223 ( .IN1(n30644), .IN2(n446), .IN3(n30652), .IN4(n489), .Q(n5272)
         );
  OA221X1 U5224 ( .IN1(n30596), .IN2(n532), .IN3(n30604), .IN4(n575), .IN5(
        n5273), .Q(n5266) );
  OA22X1 U5225 ( .IN1(n30612), .IN2(n618), .IN3(n30620), .IN4(n661), .Q(n5273)
         );
  NAND4X0 U5226 ( .IN1(n5274), .IN2(n5275), .IN3(n5276), .IN4(n5277), .QN(
        n5264) );
  OA221X1 U5227 ( .IN1(n30564), .IN2(n16), .IN3(n30572), .IN4(n59), .IN5(n5278), .Q(n5277) );
  OA22X1 U5228 ( .IN1(n30580), .IN2(n102), .IN3(n30588), .IN4(n145), .Q(n5278)
         );
  OA221X1 U5229 ( .IN1(n30532), .IN2(n188), .IN3(n30540), .IN4(n231), .IN5(
        n5279), .Q(n5276) );
  OA22X1 U5230 ( .IN1(n30548), .IN2(n274), .IN3(n30556), .IN4(n317), .Q(n5279)
         );
  OA221X1 U5231 ( .IN1(n30500), .IN2(n360), .IN3(n30508), .IN4(n403), .IN5(
        n5280), .Q(n5275) );
  OA22X1 U5232 ( .IN1(n30516), .IN2(n446), .IN3(n30524), .IN4(n489), .Q(n5280)
         );
  OA221X1 U5233 ( .IN1(n30468), .IN2(n532), .IN3(n30476), .IN4(n575), .IN5(
        n5281), .Q(n5274) );
  OA22X1 U5234 ( .IN1(n30484), .IN2(n618), .IN3(n30492), .IN4(n661), .Q(n5281)
         );
  NAND4X0 U5235 ( .IN1(n5282), .IN2(n5283), .IN3(n5284), .IN4(n5285), .QN(
        n5262) );
  OA221X1 U5236 ( .IN1(n30436), .IN2(n16), .IN3(n30444), .IN4(n59), .IN5(n5286), .Q(n5285) );
  OA22X1 U5237 ( .IN1(n30452), .IN2(n102), .IN3(n30460), .IN4(n145), .Q(n5286)
         );
  OA221X1 U5238 ( .IN1(n30404), .IN2(n188), .IN3(n30412), .IN4(n231), .IN5(
        n5287), .Q(n5284) );
  OA22X1 U5239 ( .IN1(n30420), .IN2(n274), .IN3(n30428), .IN4(n317), .Q(n5287)
         );
  OA221X1 U5240 ( .IN1(n30372), .IN2(n360), .IN3(n30380), .IN4(n403), .IN5(
        n5288), .Q(n5283) );
  OA22X1 U5241 ( .IN1(n30388), .IN2(n446), .IN3(n30396), .IN4(n489), .Q(n5288)
         );
  OA221X1 U5242 ( .IN1(n30340), .IN2(n532), .IN3(n30348), .IN4(n575), .IN5(
        n5289), .Q(n5282) );
  OA22X1 U5243 ( .IN1(n30356), .IN2(n618), .IN3(n30364), .IN4(n661), .Q(n5289)
         );
  NAND4X0 U5244 ( .IN1(n5290), .IN2(n5291), .IN3(n5292), .IN4(n5293), .QN(
        n5261) );
  OA221X1 U5245 ( .IN1(n30308), .IN2(n16), .IN3(n30316), .IN4(n59), .IN5(n5294), .Q(n5293) );
  OA22X1 U5246 ( .IN1(n30324), .IN2(n102), .IN3(n30332), .IN4(n145), .Q(n5294)
         );
  OA221X1 U5247 ( .IN1(n30276), .IN2(n188), .IN3(n30284), .IN4(n231), .IN5(
        n5295), .Q(n5292) );
  OA22X1 U5248 ( .IN1(n30292), .IN2(n274), .IN3(n30300), .IN4(n317), .Q(n5295)
         );
  OA221X1 U5249 ( .IN1(n30244), .IN2(n360), .IN3(n30252), .IN4(n403), .IN5(
        n5296), .Q(n5291) );
  OA22X1 U5250 ( .IN1(n30260), .IN2(n446), .IN3(n30268), .IN4(n489), .Q(n5296)
         );
  OA221X1 U5251 ( .IN1(n30212), .IN2(n532), .IN3(n30220), .IN4(n575), .IN5(
        n5297), .Q(n5290) );
  OA22X1 U5252 ( .IN1(n30228), .IN2(n618), .IN3(n30236), .IN4(n661), .Q(n5297)
         );
  AO221X1 U5253 ( .IN1(n2246), .IN2(n5298), .IN3(n2248), .IN4(n5299), .IN5(
        n5300), .Q(n5259) );
  AO22X1 U5254 ( .IN1(n2251), .IN2(n5301), .IN3(n2253), .IN4(n5302), .Q(n5300)
         );
  NAND4X0 U5255 ( .IN1(n5303), .IN2(n5304), .IN3(n5305), .IN4(n5306), .QN(
        n5302) );
  OA221X1 U5256 ( .IN1(n30180), .IN2(n16), .IN3(n30188), .IN4(n59), .IN5(n5307), .Q(n5306) );
  OA22X1 U5257 ( .IN1(n30196), .IN2(n102), .IN3(n30204), .IN4(n145), .Q(n5307)
         );
  OA221X1 U5258 ( .IN1(n30148), .IN2(n188), .IN3(n30156), .IN4(n231), .IN5(
        n5308), .Q(n5305) );
  OA22X1 U5259 ( .IN1(n30164), .IN2(n274), .IN3(n30172), .IN4(n317), .Q(n5308)
         );
  OA221X1 U5260 ( .IN1(n30116), .IN2(n360), .IN3(n30124), .IN4(n403), .IN5(
        n5309), .Q(n5304) );
  OA22X1 U5261 ( .IN1(n30132), .IN2(n446), .IN3(n30140), .IN4(n489), .Q(n5309)
         );
  OA221X1 U5262 ( .IN1(n30084), .IN2(n532), .IN3(n30092), .IN4(n575), .IN5(
        n5310), .Q(n5303) );
  OA22X1 U5263 ( .IN1(n30100), .IN2(n618), .IN3(n30108), .IN4(n661), .Q(n5310)
         );
  NAND4X0 U5264 ( .IN1(n5311), .IN2(n5312), .IN3(n5313), .IN4(n5314), .QN(
        n5301) );
  OA221X1 U5265 ( .IN1(n30052), .IN2(n16), .IN3(n30060), .IN4(n59), .IN5(n5315), .Q(n5314) );
  OA22X1 U5266 ( .IN1(n30068), .IN2(n102), .IN3(n30076), .IN4(n145), .Q(n5315)
         );
  OA221X1 U5267 ( .IN1(n30020), .IN2(n188), .IN3(n30028), .IN4(n231), .IN5(
        n5316), .Q(n5313) );
  OA22X1 U5268 ( .IN1(n30036), .IN2(n274), .IN3(n30044), .IN4(n317), .Q(n5316)
         );
  OA221X1 U5269 ( .IN1(n29988), .IN2(n360), .IN3(n29996), .IN4(n403), .IN5(
        n5317), .Q(n5312) );
  OA22X1 U5270 ( .IN1(n30004), .IN2(n446), .IN3(n30012), .IN4(n489), .Q(n5317)
         );
  OA221X1 U5271 ( .IN1(n29956), .IN2(n532), .IN3(n29964), .IN4(n575), .IN5(
        n5318), .Q(n5311) );
  OA22X1 U5272 ( .IN1(n29972), .IN2(n618), .IN3(n29980), .IN4(n661), .Q(n5318)
         );
  NAND4X0 U5273 ( .IN1(n5319), .IN2(n5320), .IN3(n5321), .IN4(n5322), .QN(
        n5299) );
  OA221X1 U5274 ( .IN1(n29924), .IN2(n16), .IN3(n29932), .IN4(n59), .IN5(n5323), .Q(n5322) );
  OA22X1 U5275 ( .IN1(n29940), .IN2(n102), .IN3(n29948), .IN4(n145), .Q(n5323)
         );
  OA221X1 U5276 ( .IN1(n29892), .IN2(n188), .IN3(n29900), .IN4(n231), .IN5(
        n5324), .Q(n5321) );
  OA22X1 U5277 ( .IN1(n29908), .IN2(n274), .IN3(n29916), .IN4(n317), .Q(n5324)
         );
  OA221X1 U5278 ( .IN1(n29860), .IN2(n360), .IN3(n29868), .IN4(n403), .IN5(
        n5325), .Q(n5320) );
  OA22X1 U5279 ( .IN1(n29876), .IN2(n446), .IN3(n29884), .IN4(n489), .Q(n5325)
         );
  OA221X1 U5280 ( .IN1(n29828), .IN2(n532), .IN3(n29836), .IN4(n575), .IN5(
        n5326), .Q(n5319) );
  OA22X1 U5281 ( .IN1(n29844), .IN2(n618), .IN3(n29852), .IN4(n661), .Q(n5326)
         );
  NAND4X0 U5282 ( .IN1(n5327), .IN2(n5328), .IN3(n5329), .IN4(n5330), .QN(
        n5298) );
  OA221X1 U5283 ( .IN1(n29796), .IN2(n16), .IN3(n29804), .IN4(n59), .IN5(n5331), .Q(n5330) );
  OA22X1 U5284 ( .IN1(n29812), .IN2(n102), .IN3(n29820), .IN4(n145), .Q(n5331)
         );
  OA221X1 U5285 ( .IN1(n29764), .IN2(n188), .IN3(n29772), .IN4(n231), .IN5(
        n5332), .Q(n5329) );
  OA22X1 U5286 ( .IN1(n29780), .IN2(n274), .IN3(n29788), .IN4(n317), .Q(n5332)
         );
  OA221X1 U5287 ( .IN1(n29732), .IN2(n360), .IN3(n29740), .IN4(n403), .IN5(
        n5333), .Q(n5328) );
  OA22X1 U5288 ( .IN1(n29748), .IN2(n446), .IN3(n29756), .IN4(n489), .Q(n5333)
         );
  OA221X1 U5289 ( .IN1(n29700), .IN2(n532), .IN3(n29708), .IN4(n575), .IN5(
        n5334), .Q(n5327) );
  OA22X1 U5290 ( .IN1(n29716), .IN2(n618), .IN3(n29724), .IN4(n661), .Q(n5334)
         );
  AO221X1 U5291 ( .IN1(n2287), .IN2(n5335), .IN3(n2289), .IN4(n5336), .IN5(
        n5337), .Q(n5258) );
  AO22X1 U5292 ( .IN1(n2292), .IN2(n5338), .IN3(n2294), .IN4(n5339), .Q(n5337)
         );
  NAND4X0 U5293 ( .IN1(n5340), .IN2(n5341), .IN3(n5342), .IN4(n5343), .QN(
        n5339) );
  OA221X1 U5294 ( .IN1(n31716), .IN2(n16), .IN3(n31724), .IN4(n59), .IN5(n5344), .Q(n5343) );
  OA22X1 U5295 ( .IN1(n31732), .IN2(n102), .IN3(n31740), .IN4(n145), .Q(n5344)
         );
  OA221X1 U5296 ( .IN1(n31684), .IN2(n188), .IN3(n31692), .IN4(n231), .IN5(
        n5345), .Q(n5342) );
  OA22X1 U5297 ( .IN1(n31700), .IN2(n274), .IN3(n31708), .IN4(n317), .Q(n5345)
         );
  OA221X1 U5298 ( .IN1(n31652), .IN2(n360), .IN3(n31660), .IN4(n403), .IN5(
        n5346), .Q(n5341) );
  OA22X1 U5299 ( .IN1(n31668), .IN2(n446), .IN3(n31676), .IN4(n489), .Q(n5346)
         );
  OA221X1 U5300 ( .IN1(n31620), .IN2(n532), .IN3(n31628), .IN4(n575), .IN5(
        n5347), .Q(n5340) );
  OA22X1 U5301 ( .IN1(n31636), .IN2(n618), .IN3(n31644), .IN4(n661), .Q(n5347)
         );
  NAND4X0 U5302 ( .IN1(n5348), .IN2(n5349), .IN3(n5350), .IN4(n5351), .QN(
        n5338) );
  OA221X1 U5303 ( .IN1(n31588), .IN2(n16), .IN3(n31596), .IN4(n59), .IN5(n5352), .Q(n5351) );
  OA22X1 U5304 ( .IN1(n31604), .IN2(n102), .IN3(n31612), .IN4(n145), .Q(n5352)
         );
  OA221X1 U5305 ( .IN1(n31556), .IN2(n188), .IN3(n31564), .IN4(n231), .IN5(
        n5353), .Q(n5350) );
  OA22X1 U5306 ( .IN1(n31572), .IN2(n274), .IN3(n31580), .IN4(n317), .Q(n5353)
         );
  OA221X1 U5307 ( .IN1(n31524), .IN2(n360), .IN3(n31532), .IN4(n403), .IN5(
        n5354), .Q(n5349) );
  OA22X1 U5308 ( .IN1(n31540), .IN2(n446), .IN3(n31548), .IN4(n489), .Q(n5354)
         );
  OA221X1 U5309 ( .IN1(n31492), .IN2(n532), .IN3(n31500), .IN4(n575), .IN5(
        n5355), .Q(n5348) );
  OA22X1 U5310 ( .IN1(n31508), .IN2(n618), .IN3(n31516), .IN4(n661), .Q(n5355)
         );
  NAND4X0 U5311 ( .IN1(n5356), .IN2(n5357), .IN3(n5358), .IN4(n5359), .QN(
        n5336) );
  OA221X1 U5312 ( .IN1(n31460), .IN2(n16), .IN3(n31468), .IN4(n59), .IN5(n5360), .Q(n5359) );
  OA22X1 U5313 ( .IN1(n31476), .IN2(n102), .IN3(n31484), .IN4(n145), .Q(n5360)
         );
  OA221X1 U5314 ( .IN1(n31428), .IN2(n188), .IN3(n31436), .IN4(n231), .IN5(
        n5361), .Q(n5358) );
  OA22X1 U5315 ( .IN1(n31444), .IN2(n274), .IN3(n31452), .IN4(n317), .Q(n5361)
         );
  OA221X1 U5316 ( .IN1(n31396), .IN2(n360), .IN3(n31404), .IN4(n403), .IN5(
        n5362), .Q(n5357) );
  OA22X1 U5317 ( .IN1(n31412), .IN2(n446), .IN3(n31420), .IN4(n489), .Q(n5362)
         );
  OA221X1 U5318 ( .IN1(n31364), .IN2(n532), .IN3(n31372), .IN4(n575), .IN5(
        n5363), .Q(n5356) );
  OA22X1 U5319 ( .IN1(n31380), .IN2(n618), .IN3(n31388), .IN4(n661), .Q(n5363)
         );
  NAND4X0 U5320 ( .IN1(n5364), .IN2(n5365), .IN3(n5366), .IN4(n5367), .QN(
        n5335) );
  OA221X1 U5321 ( .IN1(n31332), .IN2(n16), .IN3(n31340), .IN4(n59), .IN5(n5368), .Q(n5367) );
  OA22X1 U5322 ( .IN1(n31348), .IN2(n102), .IN3(n31356), .IN4(n145), .Q(n5368)
         );
  OA221X1 U5323 ( .IN1(n31300), .IN2(n188), .IN3(n31308), .IN4(n231), .IN5(
        n5369), .Q(n5366) );
  OA22X1 U5324 ( .IN1(n31316), .IN2(n274), .IN3(n31324), .IN4(n317), .Q(n5369)
         );
  OA221X1 U5325 ( .IN1(n31268), .IN2(n360), .IN3(n31276), .IN4(n403), .IN5(
        n5370), .Q(n5365) );
  OA22X1 U5326 ( .IN1(n31284), .IN2(n446), .IN3(n31292), .IN4(n489), .Q(n5370)
         );
  OA221X1 U5327 ( .IN1(n31236), .IN2(n532), .IN3(n31244), .IN4(n575), .IN5(
        n5371), .Q(n5364) );
  OA22X1 U5328 ( .IN1(n31252), .IN2(n618), .IN3(n31260), .IN4(n661), .Q(n5371)
         );
  AO221X1 U5329 ( .IN1(n2328), .IN2(n5372), .IN3(n2330), .IN4(n5373), .IN5(
        n5374), .Q(n5257) );
  AO22X1 U5330 ( .IN1(n2333), .IN2(n5375), .IN3(n2335), .IN4(n5376), .Q(n5374)
         );
  NAND4X0 U5331 ( .IN1(n5377), .IN2(n5378), .IN3(n5379), .IN4(n5380), .QN(
        n5376) );
  OA221X1 U5332 ( .IN1(n31204), .IN2(n15), .IN3(n31212), .IN4(n58), .IN5(n5381), .Q(n5380) );
  OA22X1 U5333 ( .IN1(n31220), .IN2(n101), .IN3(n31228), .IN4(n144), .Q(n5381)
         );
  OA221X1 U5334 ( .IN1(n31172), .IN2(n187), .IN3(n31180), .IN4(n230), .IN5(
        n5382), .Q(n5379) );
  OA22X1 U5335 ( .IN1(n31188), .IN2(n273), .IN3(n31196), .IN4(n316), .Q(n5382)
         );
  OA221X1 U5336 ( .IN1(n31140), .IN2(n359), .IN3(n31148), .IN4(n402), .IN5(
        n5383), .Q(n5378) );
  OA22X1 U5337 ( .IN1(n31156), .IN2(n445), .IN3(n31164), .IN4(n488), .Q(n5383)
         );
  OA221X1 U5338 ( .IN1(n31108), .IN2(n531), .IN3(n31116), .IN4(n574), .IN5(
        n5384), .Q(n5377) );
  OA22X1 U5339 ( .IN1(n31124), .IN2(n617), .IN3(n31132), .IN4(n660), .Q(n5384)
         );
  NAND4X0 U5340 ( .IN1(n5385), .IN2(n5386), .IN3(n5387), .IN4(n5388), .QN(
        n5375) );
  OA221X1 U5341 ( .IN1(n31076), .IN2(n15), .IN3(n31084), .IN4(n58), .IN5(n5389), .Q(n5388) );
  OA22X1 U5342 ( .IN1(n31092), .IN2(n101), .IN3(n31100), .IN4(n144), .Q(n5389)
         );
  OA221X1 U5343 ( .IN1(n31044), .IN2(n187), .IN3(n31052), .IN4(n230), .IN5(
        n5390), .Q(n5387) );
  OA22X1 U5344 ( .IN1(n31060), .IN2(n273), .IN3(n31068), .IN4(n316), .Q(n5390)
         );
  OA221X1 U5345 ( .IN1(n31012), .IN2(n359), .IN3(n31020), .IN4(n402), .IN5(
        n5391), .Q(n5386) );
  OA22X1 U5346 ( .IN1(n31028), .IN2(n445), .IN3(n31036), .IN4(n488), .Q(n5391)
         );
  OA221X1 U5347 ( .IN1(n30980), .IN2(n531), .IN3(n30988), .IN4(n574), .IN5(
        n5392), .Q(n5385) );
  OA22X1 U5348 ( .IN1(n30996), .IN2(n617), .IN3(n31004), .IN4(n660), .Q(n5392)
         );
  NAND4X0 U5349 ( .IN1(n5393), .IN2(n5394), .IN3(n5395), .IN4(n5396), .QN(
        n5373) );
  OA221X1 U5350 ( .IN1(n30948), .IN2(n15), .IN3(n30956), .IN4(n58), .IN5(n5397), .Q(n5396) );
  OA22X1 U5351 ( .IN1(n30964), .IN2(n101), .IN3(n30972), .IN4(n144), .Q(n5397)
         );
  OA221X1 U5352 ( .IN1(n30916), .IN2(n187), .IN3(n30924), .IN4(n230), .IN5(
        n5398), .Q(n5395) );
  OA22X1 U5353 ( .IN1(n30932), .IN2(n273), .IN3(n30940), .IN4(n316), .Q(n5398)
         );
  OA221X1 U5354 ( .IN1(n30884), .IN2(n359), .IN3(n30892), .IN4(n402), .IN5(
        n5399), .Q(n5394) );
  OA22X1 U5355 ( .IN1(n30900), .IN2(n445), .IN3(n30908), .IN4(n488), .Q(n5399)
         );
  OA221X1 U5356 ( .IN1(n30852), .IN2(n531), .IN3(n30860), .IN4(n574), .IN5(
        n5400), .Q(n5393) );
  OA22X1 U5357 ( .IN1(n30868), .IN2(n617), .IN3(n30876), .IN4(n660), .Q(n5400)
         );
  NAND4X0 U5358 ( .IN1(n5401), .IN2(n5402), .IN3(n5403), .IN4(n5404), .QN(
        n5372) );
  OA221X1 U5359 ( .IN1(n30820), .IN2(n15), .IN3(n30828), .IN4(n58), .IN5(n5405), .Q(n5404) );
  OA22X1 U5360 ( .IN1(n30836), .IN2(n101), .IN3(n30844), .IN4(n144), .Q(n5405)
         );
  OA221X1 U5361 ( .IN1(n30788), .IN2(n187), .IN3(n30796), .IN4(n230), .IN5(
        n5406), .Q(n5403) );
  OA22X1 U5362 ( .IN1(n30804), .IN2(n273), .IN3(n30812), .IN4(n316), .Q(n5406)
         );
  OA221X1 U5363 ( .IN1(n30756), .IN2(n359), .IN3(n30764), .IN4(n402), .IN5(
        n5407), .Q(n5402) );
  OA22X1 U5364 ( .IN1(n30772), .IN2(n445), .IN3(n30780), .IN4(n488), .Q(n5407)
         );
  OA221X1 U5365 ( .IN1(n30724), .IN2(n531), .IN3(n30732), .IN4(n574), .IN5(
        n5408), .Q(n5401) );
  OA22X1 U5366 ( .IN1(n30740), .IN2(n617), .IN3(n30748), .IN4(n660), .Q(n5408)
         );
  OR4X1 U5367 ( .IN1(n5409), .IN2(n5410), .IN3(n5411), .IN4(n5412), .Q(n2181)
         );
  AO221X1 U5368 ( .IN1(n2157), .IN2(n5413), .IN3(n2159), .IN4(n5414), .IN5(
        n5415), .Q(n5412) );
  AO22X1 U5369 ( .IN1(n2162), .IN2(n5416), .IN3(n2164), .IN4(n5417), .Q(n5415)
         );
  NAND4X0 U5370 ( .IN1(n5418), .IN2(n5419), .IN3(n5420), .IN4(n5421), .QN(
        n5417) );
  OA221X1 U5371 ( .IN1(n30691), .IN2(n15), .IN3(n30699), .IN4(n58), .IN5(n5422), .Q(n5421) );
  OA22X1 U5372 ( .IN1(n30707), .IN2(n101), .IN3(n30715), .IN4(n144), .Q(n5422)
         );
  OA221X1 U5373 ( .IN1(n30659), .IN2(n187), .IN3(n30667), .IN4(n230), .IN5(
        n5423), .Q(n5420) );
  OA22X1 U5374 ( .IN1(n30675), .IN2(n273), .IN3(n30683), .IN4(n316), .Q(n5423)
         );
  OA221X1 U5375 ( .IN1(n30627), .IN2(n359), .IN3(n30635), .IN4(n402), .IN5(
        n5424), .Q(n5419) );
  OA22X1 U5376 ( .IN1(n30643), .IN2(n445), .IN3(n30651), .IN4(n488), .Q(n5424)
         );
  OA221X1 U5377 ( .IN1(n30595), .IN2(n531), .IN3(n30603), .IN4(n574), .IN5(
        n5425), .Q(n5418) );
  OA22X1 U5378 ( .IN1(n30611), .IN2(n617), .IN3(n30619), .IN4(n660), .Q(n5425)
         );
  NAND4X0 U5379 ( .IN1(n5426), .IN2(n5427), .IN3(n5428), .IN4(n5429), .QN(
        n5416) );
  OA221X1 U5380 ( .IN1(n30563), .IN2(n15), .IN3(n30571), .IN4(n58), .IN5(n5430), .Q(n5429) );
  OA22X1 U5381 ( .IN1(n30579), .IN2(n101), .IN3(n30587), .IN4(n144), .Q(n5430)
         );
  OA221X1 U5382 ( .IN1(n30531), .IN2(n187), .IN3(n30539), .IN4(n230), .IN5(
        n5431), .Q(n5428) );
  OA22X1 U5383 ( .IN1(n30547), .IN2(n273), .IN3(n30555), .IN4(n316), .Q(n5431)
         );
  OA221X1 U5384 ( .IN1(n30499), .IN2(n359), .IN3(n30507), .IN4(n402), .IN5(
        n5432), .Q(n5427) );
  OA22X1 U5385 ( .IN1(n30515), .IN2(n445), .IN3(n30523), .IN4(n488), .Q(n5432)
         );
  OA221X1 U5386 ( .IN1(n30467), .IN2(n531), .IN3(n30475), .IN4(n574), .IN5(
        n5433), .Q(n5426) );
  OA22X1 U5387 ( .IN1(n30483), .IN2(n617), .IN3(n30491), .IN4(n660), .Q(n5433)
         );
  NAND4X0 U5388 ( .IN1(n5434), .IN2(n5435), .IN3(n5436), .IN4(n5437), .QN(
        n5414) );
  OA221X1 U5389 ( .IN1(n30435), .IN2(n15), .IN3(n30443), .IN4(n58), .IN5(n5438), .Q(n5437) );
  OA22X1 U5390 ( .IN1(n30451), .IN2(n101), .IN3(n30459), .IN4(n144), .Q(n5438)
         );
  OA221X1 U5391 ( .IN1(n30403), .IN2(n187), .IN3(n30411), .IN4(n230), .IN5(
        n5439), .Q(n5436) );
  OA22X1 U5392 ( .IN1(n30419), .IN2(n273), .IN3(n30427), .IN4(n316), .Q(n5439)
         );
  OA221X1 U5393 ( .IN1(n30371), .IN2(n359), .IN3(n30379), .IN4(n402), .IN5(
        n5440), .Q(n5435) );
  OA22X1 U5394 ( .IN1(n30387), .IN2(n445), .IN3(n30395), .IN4(n488), .Q(n5440)
         );
  OA221X1 U5395 ( .IN1(n30339), .IN2(n531), .IN3(n30347), .IN4(n574), .IN5(
        n5441), .Q(n5434) );
  OA22X1 U5396 ( .IN1(n30355), .IN2(n617), .IN3(n30363), .IN4(n660), .Q(n5441)
         );
  NAND4X0 U5397 ( .IN1(n5442), .IN2(n5443), .IN3(n5444), .IN4(n5445), .QN(
        n5413) );
  OA221X1 U5398 ( .IN1(n30307), .IN2(n15), .IN3(n30315), .IN4(n58), .IN5(n5446), .Q(n5445) );
  OA22X1 U5399 ( .IN1(n30323), .IN2(n101), .IN3(n30331), .IN4(n144), .Q(n5446)
         );
  OA221X1 U5400 ( .IN1(n30275), .IN2(n187), .IN3(n30283), .IN4(n230), .IN5(
        n5447), .Q(n5444) );
  OA22X1 U5401 ( .IN1(n30291), .IN2(n273), .IN3(n30299), .IN4(n316), .Q(n5447)
         );
  OA221X1 U5402 ( .IN1(n30243), .IN2(n359), .IN3(n30251), .IN4(n402), .IN5(
        n5448), .Q(n5443) );
  OA22X1 U5403 ( .IN1(n30259), .IN2(n445), .IN3(n30267), .IN4(n488), .Q(n5448)
         );
  OA221X1 U5404 ( .IN1(n30211), .IN2(n531), .IN3(n30219), .IN4(n574), .IN5(
        n5449), .Q(n5442) );
  OA22X1 U5405 ( .IN1(n30227), .IN2(n617), .IN3(n30235), .IN4(n660), .Q(n5449)
         );
  AO221X1 U5406 ( .IN1(n2246), .IN2(n5450), .IN3(n2248), .IN4(n5451), .IN5(
        n5452), .Q(n5411) );
  AO22X1 U5407 ( .IN1(n2251), .IN2(n5453), .IN3(n2253), .IN4(n5454), .Q(n5452)
         );
  NAND4X0 U5408 ( .IN1(n5455), .IN2(n5456), .IN3(n5457), .IN4(n5458), .QN(
        n5454) );
  OA221X1 U5409 ( .IN1(n30179), .IN2(n15), .IN3(n30187), .IN4(n58), .IN5(n5459), .Q(n5458) );
  OA22X1 U5410 ( .IN1(n30195), .IN2(n101), .IN3(n30203), .IN4(n144), .Q(n5459)
         );
  OA221X1 U5411 ( .IN1(n30147), .IN2(n187), .IN3(n30155), .IN4(n230), .IN5(
        n5460), .Q(n5457) );
  OA22X1 U5412 ( .IN1(n30163), .IN2(n273), .IN3(n30171), .IN4(n316), .Q(n5460)
         );
  OA221X1 U5413 ( .IN1(n30115), .IN2(n359), .IN3(n30123), .IN4(n402), .IN5(
        n5461), .Q(n5456) );
  OA22X1 U5414 ( .IN1(n30131), .IN2(n445), .IN3(n30139), .IN4(n488), .Q(n5461)
         );
  OA221X1 U5415 ( .IN1(n30083), .IN2(n531), .IN3(n30091), .IN4(n574), .IN5(
        n5462), .Q(n5455) );
  OA22X1 U5416 ( .IN1(n30099), .IN2(n617), .IN3(n30107), .IN4(n660), .Q(n5462)
         );
  NAND4X0 U5417 ( .IN1(n5463), .IN2(n5464), .IN3(n5465), .IN4(n5466), .QN(
        n5453) );
  OA221X1 U5418 ( .IN1(n30051), .IN2(n15), .IN3(n30059), .IN4(n58), .IN5(n5467), .Q(n5466) );
  OA22X1 U5419 ( .IN1(n30067), .IN2(n101), .IN3(n30075), .IN4(n144), .Q(n5467)
         );
  OA221X1 U5420 ( .IN1(n30019), .IN2(n187), .IN3(n30027), .IN4(n230), .IN5(
        n5468), .Q(n5465) );
  OA22X1 U5421 ( .IN1(n30035), .IN2(n273), .IN3(n30043), .IN4(n316), .Q(n5468)
         );
  OA221X1 U5422 ( .IN1(n29987), .IN2(n359), .IN3(n29995), .IN4(n402), .IN5(
        n5469), .Q(n5464) );
  OA22X1 U5423 ( .IN1(n30003), .IN2(n445), .IN3(n30011), .IN4(n488), .Q(n5469)
         );
  OA221X1 U5424 ( .IN1(n29955), .IN2(n531), .IN3(n29963), .IN4(n574), .IN5(
        n5470), .Q(n5463) );
  OA22X1 U5425 ( .IN1(n29971), .IN2(n617), .IN3(n29979), .IN4(n660), .Q(n5470)
         );
  NAND4X0 U5426 ( .IN1(n5471), .IN2(n5472), .IN3(n5473), .IN4(n5474), .QN(
        n5451) );
  OA221X1 U5427 ( .IN1(n29923), .IN2(n15), .IN3(n29931), .IN4(n58), .IN5(n5475), .Q(n5474) );
  OA22X1 U5428 ( .IN1(n29939), .IN2(n101), .IN3(n29947), .IN4(n144), .Q(n5475)
         );
  OA221X1 U5429 ( .IN1(n29891), .IN2(n187), .IN3(n29899), .IN4(n230), .IN5(
        n5476), .Q(n5473) );
  OA22X1 U5430 ( .IN1(n29907), .IN2(n273), .IN3(n29915), .IN4(n316), .Q(n5476)
         );
  OA221X1 U5431 ( .IN1(n29859), .IN2(n359), .IN3(n29867), .IN4(n402), .IN5(
        n5477), .Q(n5472) );
  OA22X1 U5432 ( .IN1(n29875), .IN2(n445), .IN3(n29883), .IN4(n488), .Q(n5477)
         );
  OA221X1 U5433 ( .IN1(n29827), .IN2(n531), .IN3(n29835), .IN4(n574), .IN5(
        n5478), .Q(n5471) );
  OA22X1 U5434 ( .IN1(n29843), .IN2(n617), .IN3(n29851), .IN4(n660), .Q(n5478)
         );
  NAND4X0 U5435 ( .IN1(n5479), .IN2(n5480), .IN3(n5481), .IN4(n5482), .QN(
        n5450) );
  OA221X1 U5436 ( .IN1(n29795), .IN2(n15), .IN3(n29803), .IN4(n58), .IN5(n5483), .Q(n5482) );
  OA22X1 U5437 ( .IN1(n29811), .IN2(n101), .IN3(n29819), .IN4(n144), .Q(n5483)
         );
  OA221X1 U5438 ( .IN1(n29763), .IN2(n187), .IN3(n29771), .IN4(n230), .IN5(
        n5484), .Q(n5481) );
  OA22X1 U5439 ( .IN1(n29779), .IN2(n273), .IN3(n29787), .IN4(n316), .Q(n5484)
         );
  OA221X1 U5440 ( .IN1(n29731), .IN2(n359), .IN3(n29739), .IN4(n402), .IN5(
        n5485), .Q(n5480) );
  OA22X1 U5441 ( .IN1(n29747), .IN2(n445), .IN3(n29755), .IN4(n488), .Q(n5485)
         );
  OA221X1 U5442 ( .IN1(n29699), .IN2(n531), .IN3(n29707), .IN4(n574), .IN5(
        n5486), .Q(n5479) );
  OA22X1 U5443 ( .IN1(n29715), .IN2(n617), .IN3(n29723), .IN4(n660), .Q(n5486)
         );
  AO221X1 U5444 ( .IN1(n2287), .IN2(n5487), .IN3(n2289), .IN4(n5488), .IN5(
        n5489), .Q(n5410) );
  AO22X1 U5445 ( .IN1(n2292), .IN2(n5490), .IN3(n2294), .IN4(n5491), .Q(n5489)
         );
  NAND4X0 U5446 ( .IN1(n5492), .IN2(n5493), .IN3(n5494), .IN4(n5495), .QN(
        n5491) );
  OA221X1 U5447 ( .IN1(n31715), .IN2(n14), .IN3(n31723), .IN4(n57), .IN5(n5496), .Q(n5495) );
  OA22X1 U5448 ( .IN1(n31731), .IN2(n100), .IN3(n31739), .IN4(n143), .Q(n5496)
         );
  OA221X1 U5449 ( .IN1(n31683), .IN2(n186), .IN3(n31691), .IN4(n229), .IN5(
        n5497), .Q(n5494) );
  OA22X1 U5450 ( .IN1(n31699), .IN2(n272), .IN3(n31707), .IN4(n315), .Q(n5497)
         );
  OA221X1 U5451 ( .IN1(n31651), .IN2(n358), .IN3(n31659), .IN4(n401), .IN5(
        n5498), .Q(n5493) );
  OA22X1 U5452 ( .IN1(n31667), .IN2(n444), .IN3(n31675), .IN4(n487), .Q(n5498)
         );
  OA221X1 U5453 ( .IN1(n31619), .IN2(n530), .IN3(n31627), .IN4(n573), .IN5(
        n5499), .Q(n5492) );
  OA22X1 U5454 ( .IN1(n31635), .IN2(n616), .IN3(n31643), .IN4(n659), .Q(n5499)
         );
  NAND4X0 U5455 ( .IN1(n5500), .IN2(n5501), .IN3(n5502), .IN4(n5503), .QN(
        n5490) );
  OA221X1 U5456 ( .IN1(n31587), .IN2(n14), .IN3(n31595), .IN4(n57), .IN5(n5504), .Q(n5503) );
  OA22X1 U5457 ( .IN1(n31603), .IN2(n100), .IN3(n31611), .IN4(n143), .Q(n5504)
         );
  OA221X1 U5458 ( .IN1(n31555), .IN2(n186), .IN3(n31563), .IN4(n229), .IN5(
        n5505), .Q(n5502) );
  OA22X1 U5459 ( .IN1(n31571), .IN2(n272), .IN3(n31579), .IN4(n315), .Q(n5505)
         );
  OA221X1 U5460 ( .IN1(n31523), .IN2(n358), .IN3(n31531), .IN4(n401), .IN5(
        n5506), .Q(n5501) );
  OA22X1 U5461 ( .IN1(n31539), .IN2(n444), .IN3(n31547), .IN4(n487), .Q(n5506)
         );
  OA221X1 U5462 ( .IN1(n31491), .IN2(n530), .IN3(n31499), .IN4(n573), .IN5(
        n5507), .Q(n5500) );
  OA22X1 U5463 ( .IN1(n31507), .IN2(n616), .IN3(n31515), .IN4(n659), .Q(n5507)
         );
  NAND4X0 U5464 ( .IN1(n5508), .IN2(n5509), .IN3(n5510), .IN4(n5511), .QN(
        n5488) );
  OA221X1 U5465 ( .IN1(n31459), .IN2(n14), .IN3(n31467), .IN4(n57), .IN5(n5512), .Q(n5511) );
  OA22X1 U5466 ( .IN1(n31475), .IN2(n100), .IN3(n31483), .IN4(n143), .Q(n5512)
         );
  OA221X1 U5467 ( .IN1(n31427), .IN2(n186), .IN3(n31435), .IN4(n229), .IN5(
        n5513), .Q(n5510) );
  OA22X1 U5468 ( .IN1(n31443), .IN2(n272), .IN3(n31451), .IN4(n315), .Q(n5513)
         );
  OA221X1 U5469 ( .IN1(n31395), .IN2(n358), .IN3(n31403), .IN4(n401), .IN5(
        n5514), .Q(n5509) );
  OA22X1 U5470 ( .IN1(n31411), .IN2(n444), .IN3(n31419), .IN4(n487), .Q(n5514)
         );
  OA221X1 U5471 ( .IN1(n31363), .IN2(n530), .IN3(n31371), .IN4(n573), .IN5(
        n5515), .Q(n5508) );
  OA22X1 U5472 ( .IN1(n31379), .IN2(n616), .IN3(n31387), .IN4(n659), .Q(n5515)
         );
  NAND4X0 U5473 ( .IN1(n5516), .IN2(n5517), .IN3(n5518), .IN4(n5519), .QN(
        n5487) );
  OA221X1 U5474 ( .IN1(n31331), .IN2(n14), .IN3(n31339), .IN4(n57), .IN5(n5520), .Q(n5519) );
  OA22X1 U5475 ( .IN1(n31347), .IN2(n100), .IN3(n31355), .IN4(n143), .Q(n5520)
         );
  OA221X1 U5476 ( .IN1(n31299), .IN2(n186), .IN3(n31307), .IN4(n229), .IN5(
        n5521), .Q(n5518) );
  OA22X1 U5477 ( .IN1(n31315), .IN2(n272), .IN3(n31323), .IN4(n315), .Q(n5521)
         );
  OA221X1 U5478 ( .IN1(n31267), .IN2(n358), .IN3(n31275), .IN4(n401), .IN5(
        n5522), .Q(n5517) );
  OA22X1 U5479 ( .IN1(n31283), .IN2(n444), .IN3(n31291), .IN4(n487), .Q(n5522)
         );
  OA221X1 U5480 ( .IN1(n31235), .IN2(n530), .IN3(n31243), .IN4(n573), .IN5(
        n5523), .Q(n5516) );
  OA22X1 U5481 ( .IN1(n31251), .IN2(n616), .IN3(n31259), .IN4(n659), .Q(n5523)
         );
  AO221X1 U5482 ( .IN1(n2328), .IN2(n5524), .IN3(n2330), .IN4(n5525), .IN5(
        n5526), .Q(n5409) );
  AO22X1 U5483 ( .IN1(n2333), .IN2(n5527), .IN3(n2335), .IN4(n5528), .Q(n5526)
         );
  NAND4X0 U5484 ( .IN1(n5529), .IN2(n5530), .IN3(n5531), .IN4(n5532), .QN(
        n5528) );
  OA221X1 U5485 ( .IN1(n31203), .IN2(n14), .IN3(n31211), .IN4(n57), .IN5(n5533), .Q(n5532) );
  OA22X1 U5486 ( .IN1(n31219), .IN2(n100), .IN3(n31227), .IN4(n143), .Q(n5533)
         );
  OA221X1 U5487 ( .IN1(n31171), .IN2(n186), .IN3(n31179), .IN4(n229), .IN5(
        n5534), .Q(n5531) );
  OA22X1 U5488 ( .IN1(n31187), .IN2(n272), .IN3(n31195), .IN4(n315), .Q(n5534)
         );
  OA221X1 U5489 ( .IN1(n31139), .IN2(n358), .IN3(n31147), .IN4(n401), .IN5(
        n5535), .Q(n5530) );
  OA22X1 U5490 ( .IN1(n31155), .IN2(n444), .IN3(n31163), .IN4(n487), .Q(n5535)
         );
  OA221X1 U5491 ( .IN1(n31107), .IN2(n530), .IN3(n31115), .IN4(n573), .IN5(
        n5536), .Q(n5529) );
  OA22X1 U5492 ( .IN1(n31123), .IN2(n616), .IN3(n31131), .IN4(n659), .Q(n5536)
         );
  NAND4X0 U5493 ( .IN1(n5537), .IN2(n5538), .IN3(n5539), .IN4(n5540), .QN(
        n5527) );
  OA221X1 U5494 ( .IN1(n31075), .IN2(n14), .IN3(n31083), .IN4(n57), .IN5(n5541), .Q(n5540) );
  OA22X1 U5495 ( .IN1(n31091), .IN2(n100), .IN3(n31099), .IN4(n143), .Q(n5541)
         );
  OA221X1 U5496 ( .IN1(n31043), .IN2(n186), .IN3(n31051), .IN4(n229), .IN5(
        n5542), .Q(n5539) );
  OA22X1 U5497 ( .IN1(n31059), .IN2(n272), .IN3(n31067), .IN4(n315), .Q(n5542)
         );
  OA221X1 U5498 ( .IN1(n31011), .IN2(n358), .IN3(n31019), .IN4(n401), .IN5(
        n5543), .Q(n5538) );
  OA22X1 U5499 ( .IN1(n31027), .IN2(n444), .IN3(n31035), .IN4(n487), .Q(n5543)
         );
  OA221X1 U5500 ( .IN1(n30979), .IN2(n530), .IN3(n30987), .IN4(n573), .IN5(
        n5544), .Q(n5537) );
  OA22X1 U5501 ( .IN1(n30995), .IN2(n616), .IN3(n31003), .IN4(n659), .Q(n5544)
         );
  NAND4X0 U5502 ( .IN1(n5545), .IN2(n5546), .IN3(n5547), .IN4(n5548), .QN(
        n5525) );
  OA221X1 U5503 ( .IN1(n30947), .IN2(n14), .IN3(n30955), .IN4(n57), .IN5(n5549), .Q(n5548) );
  OA22X1 U5504 ( .IN1(n30963), .IN2(n100), .IN3(n30971), .IN4(n143), .Q(n5549)
         );
  OA221X1 U5505 ( .IN1(n30915), .IN2(n186), .IN3(n30923), .IN4(n229), .IN5(
        n5550), .Q(n5547) );
  OA22X1 U5506 ( .IN1(n30931), .IN2(n272), .IN3(n30939), .IN4(n315), .Q(n5550)
         );
  OA221X1 U5507 ( .IN1(n30883), .IN2(n358), .IN3(n30891), .IN4(n401), .IN5(
        n5551), .Q(n5546) );
  OA22X1 U5508 ( .IN1(n30899), .IN2(n444), .IN3(n30907), .IN4(n487), .Q(n5551)
         );
  OA221X1 U5509 ( .IN1(n30851), .IN2(n530), .IN3(n30859), .IN4(n573), .IN5(
        n5552), .Q(n5545) );
  OA22X1 U5510 ( .IN1(n30867), .IN2(n616), .IN3(n30875), .IN4(n659), .Q(n5552)
         );
  NAND4X0 U5511 ( .IN1(n5553), .IN2(n5554), .IN3(n5555), .IN4(n5556), .QN(
        n5524) );
  OA221X1 U5512 ( .IN1(n30819), .IN2(n14), .IN3(n30827), .IN4(n57), .IN5(n5557), .Q(n5556) );
  OA22X1 U5513 ( .IN1(n30835), .IN2(n100), .IN3(n30843), .IN4(n143), .Q(n5557)
         );
  OA221X1 U5514 ( .IN1(n30787), .IN2(n186), .IN3(n30795), .IN4(n229), .IN5(
        n5558), .Q(n5555) );
  OA22X1 U5515 ( .IN1(n30803), .IN2(n272), .IN3(n30811), .IN4(n315), .Q(n5558)
         );
  OA221X1 U5516 ( .IN1(n30755), .IN2(n358), .IN3(n30763), .IN4(n401), .IN5(
        n5559), .Q(n5554) );
  OA22X1 U5517 ( .IN1(n30771), .IN2(n444), .IN3(n30779), .IN4(n487), .Q(n5559)
         );
  OA221X1 U5518 ( .IN1(n30723), .IN2(n530), .IN3(n30731), .IN4(n573), .IN5(
        n5560), .Q(n5553) );
  OA22X1 U5519 ( .IN1(n30739), .IN2(n616), .IN3(n30747), .IN4(n659), .Q(n5560)
         );
  OR4X1 U5520 ( .IN1(n5561), .IN2(n5562), .IN3(n5563), .IN4(n5564), .Q(n2180)
         );
  AO221X1 U5521 ( .IN1(n2157), .IN2(n5565), .IN3(n2159), .IN4(n5566), .IN5(
        n5567), .Q(n5564) );
  AO22X1 U5522 ( .IN1(n2162), .IN2(n5568), .IN3(n2164), .IN4(n5569), .Q(n5567)
         );
  NAND4X0 U5523 ( .IN1(n5570), .IN2(n5571), .IN3(n5572), .IN4(n5573), .QN(
        n5569) );
  OA221X1 U5524 ( .IN1(n30690), .IN2(n14), .IN3(n30698), .IN4(n57), .IN5(n5574), .Q(n5573) );
  OA22X1 U5525 ( .IN1(n30706), .IN2(n100), .IN3(n30714), .IN4(n143), .Q(n5574)
         );
  OA221X1 U5526 ( .IN1(n30658), .IN2(n186), .IN3(n30666), .IN4(n229), .IN5(
        n5575), .Q(n5572) );
  OA22X1 U5527 ( .IN1(n30674), .IN2(n272), .IN3(n30682), .IN4(n315), .Q(n5575)
         );
  OA221X1 U5528 ( .IN1(n30626), .IN2(n358), .IN3(n30634), .IN4(n401), .IN5(
        n5576), .Q(n5571) );
  OA22X1 U5529 ( .IN1(n30642), .IN2(n444), .IN3(n30650), .IN4(n487), .Q(n5576)
         );
  OA221X1 U5530 ( .IN1(n30594), .IN2(n530), .IN3(n30602), .IN4(n573), .IN5(
        n5577), .Q(n5570) );
  OA22X1 U5531 ( .IN1(n30610), .IN2(n616), .IN3(n30618), .IN4(n659), .Q(n5577)
         );
  NAND4X0 U5532 ( .IN1(n5578), .IN2(n5579), .IN3(n5580), .IN4(n5581), .QN(
        n5568) );
  OA221X1 U5533 ( .IN1(n30562), .IN2(n14), .IN3(n30570), .IN4(n57), .IN5(n5582), .Q(n5581) );
  OA22X1 U5534 ( .IN1(n30578), .IN2(n100), .IN3(n30586), .IN4(n143), .Q(n5582)
         );
  OA221X1 U5535 ( .IN1(n30530), .IN2(n186), .IN3(n30538), .IN4(n229), .IN5(
        n5583), .Q(n5580) );
  OA22X1 U5536 ( .IN1(n30546), .IN2(n272), .IN3(n30554), .IN4(n315), .Q(n5583)
         );
  OA221X1 U5537 ( .IN1(n30498), .IN2(n358), .IN3(n30506), .IN4(n401), .IN5(
        n5584), .Q(n5579) );
  OA22X1 U5538 ( .IN1(n30514), .IN2(n444), .IN3(n30522), .IN4(n487), .Q(n5584)
         );
  OA221X1 U5539 ( .IN1(n30466), .IN2(n530), .IN3(n30474), .IN4(n573), .IN5(
        n5585), .Q(n5578) );
  OA22X1 U5540 ( .IN1(n30482), .IN2(n616), .IN3(n30490), .IN4(n659), .Q(n5585)
         );
  NAND4X0 U5541 ( .IN1(n5586), .IN2(n5587), .IN3(n5588), .IN4(n5589), .QN(
        n5566) );
  OA221X1 U5542 ( .IN1(n30434), .IN2(n14), .IN3(n30442), .IN4(n57), .IN5(n5590), .Q(n5589) );
  OA22X1 U5543 ( .IN1(n30450), .IN2(n100), .IN3(n30458), .IN4(n143), .Q(n5590)
         );
  OA221X1 U5544 ( .IN1(n30402), .IN2(n186), .IN3(n30410), .IN4(n229), .IN5(
        n5591), .Q(n5588) );
  OA22X1 U5545 ( .IN1(n30418), .IN2(n272), .IN3(n30426), .IN4(n315), .Q(n5591)
         );
  OA221X1 U5546 ( .IN1(n30370), .IN2(n358), .IN3(n30378), .IN4(n401), .IN5(
        n5592), .Q(n5587) );
  OA22X1 U5547 ( .IN1(n30386), .IN2(n444), .IN3(n30394), .IN4(n487), .Q(n5592)
         );
  OA221X1 U5548 ( .IN1(n30338), .IN2(n530), .IN3(n30346), .IN4(n573), .IN5(
        n5593), .Q(n5586) );
  OA22X1 U5549 ( .IN1(n30354), .IN2(n616), .IN3(n30362), .IN4(n659), .Q(n5593)
         );
  NAND4X0 U5550 ( .IN1(n5594), .IN2(n5595), .IN3(n5596), .IN4(n5597), .QN(
        n5565) );
  OA221X1 U5551 ( .IN1(n30306), .IN2(n14), .IN3(n30314), .IN4(n57), .IN5(n5598), .Q(n5597) );
  OA22X1 U5552 ( .IN1(n30322), .IN2(n100), .IN3(n30330), .IN4(n143), .Q(n5598)
         );
  OA221X1 U5553 ( .IN1(n30274), .IN2(n186), .IN3(n30282), .IN4(n229), .IN5(
        n5599), .Q(n5596) );
  OA22X1 U5554 ( .IN1(n30290), .IN2(n272), .IN3(n30298), .IN4(n315), .Q(n5599)
         );
  OA221X1 U5555 ( .IN1(n30242), .IN2(n358), .IN3(n30250), .IN4(n401), .IN5(
        n5600), .Q(n5595) );
  OA22X1 U5556 ( .IN1(n30258), .IN2(n444), .IN3(n30266), .IN4(n487), .Q(n5600)
         );
  OA221X1 U5557 ( .IN1(n30210), .IN2(n530), .IN3(n30218), .IN4(n573), .IN5(
        n5601), .Q(n5594) );
  OA22X1 U5558 ( .IN1(n30226), .IN2(n616), .IN3(n30234), .IN4(n659), .Q(n5601)
         );
  AO221X1 U5559 ( .IN1(n2246), .IN2(n5602), .IN3(n2248), .IN4(n5603), .IN5(
        n5604), .Q(n5563) );
  AO22X1 U5560 ( .IN1(n2251), .IN2(n5605), .IN3(n2253), .IN4(n5606), .Q(n5604)
         );
  NAND4X0 U5561 ( .IN1(n5607), .IN2(n5608), .IN3(n5609), .IN4(n5610), .QN(
        n5606) );
  OA221X1 U5562 ( .IN1(n30178), .IN2(n13), .IN3(n30186), .IN4(n56), .IN5(n5611), .Q(n5610) );
  OA22X1 U5563 ( .IN1(n30194), .IN2(n99), .IN3(n30202), .IN4(n142), .Q(n5611)
         );
  OA221X1 U5564 ( .IN1(n30146), .IN2(n185), .IN3(n30154), .IN4(n228), .IN5(
        n5612), .Q(n5609) );
  OA22X1 U5565 ( .IN1(n30162), .IN2(n271), .IN3(n30170), .IN4(n314), .Q(n5612)
         );
  OA221X1 U5566 ( .IN1(n30114), .IN2(n357), .IN3(n30122), .IN4(n400), .IN5(
        n5613), .Q(n5608) );
  OA22X1 U5567 ( .IN1(n30130), .IN2(n443), .IN3(n30138), .IN4(n486), .Q(n5613)
         );
  OA221X1 U5568 ( .IN1(n30082), .IN2(n529), .IN3(n30090), .IN4(n572), .IN5(
        n5614), .Q(n5607) );
  OA22X1 U5569 ( .IN1(n30098), .IN2(n615), .IN3(n30106), .IN4(n658), .Q(n5614)
         );
  NAND4X0 U5570 ( .IN1(n5615), .IN2(n5616), .IN3(n5617), .IN4(n5618), .QN(
        n5605) );
  OA221X1 U5571 ( .IN1(n30050), .IN2(n13), .IN3(n30058), .IN4(n56), .IN5(n5619), .Q(n5618) );
  OA22X1 U5572 ( .IN1(n30066), .IN2(n99), .IN3(n30074), .IN4(n142), .Q(n5619)
         );
  OA221X1 U5573 ( .IN1(n30018), .IN2(n185), .IN3(n30026), .IN4(n228), .IN5(
        n5620), .Q(n5617) );
  OA22X1 U5574 ( .IN1(n30034), .IN2(n271), .IN3(n30042), .IN4(n314), .Q(n5620)
         );
  OA221X1 U5575 ( .IN1(n29986), .IN2(n357), .IN3(n29994), .IN4(n400), .IN5(
        n5621), .Q(n5616) );
  OA22X1 U5576 ( .IN1(n30002), .IN2(n443), .IN3(n30010), .IN4(n486), .Q(n5621)
         );
  OA221X1 U5577 ( .IN1(n29954), .IN2(n529), .IN3(n29962), .IN4(n572), .IN5(
        n5622), .Q(n5615) );
  OA22X1 U5578 ( .IN1(n29970), .IN2(n615), .IN3(n29978), .IN4(n658), .Q(n5622)
         );
  NAND4X0 U5579 ( .IN1(n5623), .IN2(n5624), .IN3(n5625), .IN4(n5626), .QN(
        n5603) );
  OA221X1 U5580 ( .IN1(n29922), .IN2(n13), .IN3(n29930), .IN4(n56), .IN5(n5627), .Q(n5626) );
  OA22X1 U5581 ( .IN1(n29938), .IN2(n99), .IN3(n29946), .IN4(n142), .Q(n5627)
         );
  OA221X1 U5582 ( .IN1(n29890), .IN2(n185), .IN3(n29898), .IN4(n228), .IN5(
        n5628), .Q(n5625) );
  OA22X1 U5583 ( .IN1(n29906), .IN2(n271), .IN3(n29914), .IN4(n314), .Q(n5628)
         );
  OA221X1 U5584 ( .IN1(n29858), .IN2(n357), .IN3(n29866), .IN4(n400), .IN5(
        n5629), .Q(n5624) );
  OA22X1 U5585 ( .IN1(n29874), .IN2(n443), .IN3(n29882), .IN4(n486), .Q(n5629)
         );
  OA221X1 U5586 ( .IN1(n29826), .IN2(n529), .IN3(n29834), .IN4(n572), .IN5(
        n5630), .Q(n5623) );
  OA22X1 U5587 ( .IN1(n29842), .IN2(n615), .IN3(n29850), .IN4(n658), .Q(n5630)
         );
  NAND4X0 U5588 ( .IN1(n5631), .IN2(n5632), .IN3(n5633), .IN4(n5634), .QN(
        n5602) );
  OA221X1 U5589 ( .IN1(n29794), .IN2(n13), .IN3(n29802), .IN4(n56), .IN5(n5635), .Q(n5634) );
  OA22X1 U5590 ( .IN1(n29810), .IN2(n99), .IN3(n29818), .IN4(n142), .Q(n5635)
         );
  OA221X1 U5591 ( .IN1(n29762), .IN2(n185), .IN3(n29770), .IN4(n228), .IN5(
        n5636), .Q(n5633) );
  OA22X1 U5592 ( .IN1(n29778), .IN2(n271), .IN3(n29786), .IN4(n314), .Q(n5636)
         );
  OA221X1 U5593 ( .IN1(n29730), .IN2(n357), .IN3(n29738), .IN4(n400), .IN5(
        n5637), .Q(n5632) );
  OA22X1 U5594 ( .IN1(n29746), .IN2(n443), .IN3(n29754), .IN4(n486), .Q(n5637)
         );
  OA221X1 U5595 ( .IN1(n29698), .IN2(n529), .IN3(n29706), .IN4(n572), .IN5(
        n5638), .Q(n5631) );
  OA22X1 U5596 ( .IN1(n29714), .IN2(n615), .IN3(n29722), .IN4(n658), .Q(n5638)
         );
  AO221X1 U5597 ( .IN1(n2287), .IN2(n5639), .IN3(n2289), .IN4(n5640), .IN5(
        n5641), .Q(n5562) );
  AO22X1 U5598 ( .IN1(n2292), .IN2(n5642), .IN3(n2294), .IN4(n5643), .Q(n5641)
         );
  NAND4X0 U5599 ( .IN1(n5644), .IN2(n5645), .IN3(n5646), .IN4(n5647), .QN(
        n5643) );
  OA221X1 U5600 ( .IN1(n31714), .IN2(n13), .IN3(n31722), .IN4(n56), .IN5(n5648), .Q(n5647) );
  OA22X1 U5601 ( .IN1(n31730), .IN2(n99), .IN3(n31738), .IN4(n142), .Q(n5648)
         );
  OA221X1 U5602 ( .IN1(n31682), .IN2(n185), .IN3(n31690), .IN4(n228), .IN5(
        n5649), .Q(n5646) );
  OA22X1 U5603 ( .IN1(n31698), .IN2(n271), .IN3(n31706), .IN4(n314), .Q(n5649)
         );
  OA221X1 U5604 ( .IN1(n31650), .IN2(n357), .IN3(n31658), .IN4(n400), .IN5(
        n5650), .Q(n5645) );
  OA22X1 U5605 ( .IN1(n31666), .IN2(n443), .IN3(n31674), .IN4(n486), .Q(n5650)
         );
  OA221X1 U5606 ( .IN1(n31618), .IN2(n529), .IN3(n31626), .IN4(n572), .IN5(
        n5651), .Q(n5644) );
  OA22X1 U5607 ( .IN1(n31634), .IN2(n615), .IN3(n31642), .IN4(n658), .Q(n5651)
         );
  NAND4X0 U5608 ( .IN1(n5652), .IN2(n5653), .IN3(n5654), .IN4(n5655), .QN(
        n5642) );
  OA221X1 U5609 ( .IN1(n31586), .IN2(n13), .IN3(n31594), .IN4(n56), .IN5(n5656), .Q(n5655) );
  OA22X1 U5610 ( .IN1(n31602), .IN2(n99), .IN3(n31610), .IN4(n142), .Q(n5656)
         );
  OA221X1 U5611 ( .IN1(n31554), .IN2(n185), .IN3(n31562), .IN4(n228), .IN5(
        n5657), .Q(n5654) );
  OA22X1 U5612 ( .IN1(n31570), .IN2(n271), .IN3(n31578), .IN4(n314), .Q(n5657)
         );
  OA221X1 U5613 ( .IN1(n31522), .IN2(n357), .IN3(n31530), .IN4(n400), .IN5(
        n5658), .Q(n5653) );
  OA22X1 U5614 ( .IN1(n31538), .IN2(n443), .IN3(n31546), .IN4(n486), .Q(n5658)
         );
  OA221X1 U5615 ( .IN1(n31490), .IN2(n529), .IN3(n31498), .IN4(n572), .IN5(
        n5659), .Q(n5652) );
  OA22X1 U5616 ( .IN1(n31506), .IN2(n615), .IN3(n31514), .IN4(n658), .Q(n5659)
         );
  NAND4X0 U5617 ( .IN1(n5660), .IN2(n5661), .IN3(n5662), .IN4(n5663), .QN(
        n5640) );
  OA221X1 U5618 ( .IN1(n31458), .IN2(n13), .IN3(n31466), .IN4(n56), .IN5(n5664), .Q(n5663) );
  OA22X1 U5619 ( .IN1(n31474), .IN2(n99), .IN3(n31482), .IN4(n142), .Q(n5664)
         );
  OA221X1 U5620 ( .IN1(n31426), .IN2(n185), .IN3(n31434), .IN4(n228), .IN5(
        n5665), .Q(n5662) );
  OA22X1 U5621 ( .IN1(n31442), .IN2(n271), .IN3(n31450), .IN4(n314), .Q(n5665)
         );
  OA221X1 U5622 ( .IN1(n31394), .IN2(n357), .IN3(n31402), .IN4(n400), .IN5(
        n5666), .Q(n5661) );
  OA22X1 U5623 ( .IN1(n31410), .IN2(n443), .IN3(n31418), .IN4(n486), .Q(n5666)
         );
  OA221X1 U5624 ( .IN1(n31362), .IN2(n529), .IN3(n31370), .IN4(n572), .IN5(
        n5667), .Q(n5660) );
  OA22X1 U5625 ( .IN1(n31378), .IN2(n615), .IN3(n31386), .IN4(n658), .Q(n5667)
         );
  NAND4X0 U5626 ( .IN1(n5668), .IN2(n5669), .IN3(n5670), .IN4(n5671), .QN(
        n5639) );
  OA221X1 U5627 ( .IN1(n31330), .IN2(n13), .IN3(n31338), .IN4(n56), .IN5(n5672), .Q(n5671) );
  OA22X1 U5628 ( .IN1(n31346), .IN2(n99), .IN3(n31354), .IN4(n142), .Q(n5672)
         );
  OA221X1 U5629 ( .IN1(n31298), .IN2(n185), .IN3(n31306), .IN4(n228), .IN5(
        n5673), .Q(n5670) );
  OA22X1 U5630 ( .IN1(n31314), .IN2(n271), .IN3(n31322), .IN4(n314), .Q(n5673)
         );
  OA221X1 U5631 ( .IN1(n31266), .IN2(n357), .IN3(n31274), .IN4(n400), .IN5(
        n5674), .Q(n5669) );
  OA22X1 U5632 ( .IN1(n31282), .IN2(n443), .IN3(n31290), .IN4(n486), .Q(n5674)
         );
  OA221X1 U5633 ( .IN1(n31234), .IN2(n529), .IN3(n31242), .IN4(n572), .IN5(
        n5675), .Q(n5668) );
  OA22X1 U5634 ( .IN1(n31250), .IN2(n615), .IN3(n31258), .IN4(n658), .Q(n5675)
         );
  AO221X1 U5635 ( .IN1(n2328), .IN2(n5676), .IN3(n2330), .IN4(n5677), .IN5(
        n5678), .Q(n5561) );
  AO22X1 U5636 ( .IN1(n2333), .IN2(n5679), .IN3(n2335), .IN4(n5680), .Q(n5678)
         );
  NAND4X0 U5637 ( .IN1(n5681), .IN2(n5682), .IN3(n5683), .IN4(n5684), .QN(
        n5680) );
  OA221X1 U5638 ( .IN1(n31202), .IN2(n13), .IN3(n31210), .IN4(n56), .IN5(n5685), .Q(n5684) );
  OA22X1 U5639 ( .IN1(n31218), .IN2(n99), .IN3(n31226), .IN4(n142), .Q(n5685)
         );
  OA221X1 U5640 ( .IN1(n31170), .IN2(n185), .IN3(n31178), .IN4(n228), .IN5(
        n5686), .Q(n5683) );
  OA22X1 U5641 ( .IN1(n31186), .IN2(n271), .IN3(n31194), .IN4(n314), .Q(n5686)
         );
  OA221X1 U5642 ( .IN1(n31138), .IN2(n357), .IN3(n31146), .IN4(n400), .IN5(
        n5687), .Q(n5682) );
  OA22X1 U5643 ( .IN1(n31154), .IN2(n443), .IN3(n31162), .IN4(n486), .Q(n5687)
         );
  OA221X1 U5644 ( .IN1(n31106), .IN2(n529), .IN3(n31114), .IN4(n572), .IN5(
        n5688), .Q(n5681) );
  OA22X1 U5645 ( .IN1(n31122), .IN2(n615), .IN3(n31130), .IN4(n658), .Q(n5688)
         );
  NAND4X0 U5646 ( .IN1(n5689), .IN2(n5690), .IN3(n5691), .IN4(n5692), .QN(
        n5679) );
  OA221X1 U5647 ( .IN1(n31074), .IN2(n13), .IN3(n31082), .IN4(n56), .IN5(n5693), .Q(n5692) );
  OA22X1 U5648 ( .IN1(n31090), .IN2(n99), .IN3(n31098), .IN4(n142), .Q(n5693)
         );
  OA221X1 U5649 ( .IN1(n31042), .IN2(n185), .IN3(n31050), .IN4(n228), .IN5(
        n5694), .Q(n5691) );
  OA22X1 U5650 ( .IN1(n31058), .IN2(n271), .IN3(n31066), .IN4(n314), .Q(n5694)
         );
  OA221X1 U5651 ( .IN1(n31010), .IN2(n357), .IN3(n31018), .IN4(n400), .IN5(
        n5695), .Q(n5690) );
  OA22X1 U5652 ( .IN1(n31026), .IN2(n443), .IN3(n31034), .IN4(n486), .Q(n5695)
         );
  OA221X1 U5653 ( .IN1(n30978), .IN2(n529), .IN3(n30986), .IN4(n572), .IN5(
        n5696), .Q(n5689) );
  OA22X1 U5654 ( .IN1(n30994), .IN2(n615), .IN3(n31002), .IN4(n658), .Q(n5696)
         );
  NAND4X0 U5655 ( .IN1(n5697), .IN2(n5698), .IN3(n5699), .IN4(n5700), .QN(
        n5677) );
  OA221X1 U5656 ( .IN1(n30946), .IN2(n13), .IN3(n30954), .IN4(n56), .IN5(n5701), .Q(n5700) );
  OA22X1 U5657 ( .IN1(n30962), .IN2(n99), .IN3(n30970), .IN4(n142), .Q(n5701)
         );
  OA221X1 U5658 ( .IN1(n30914), .IN2(n185), .IN3(n30922), .IN4(n228), .IN5(
        n5702), .Q(n5699) );
  OA22X1 U5659 ( .IN1(n30930), .IN2(n271), .IN3(n30938), .IN4(n314), .Q(n5702)
         );
  OA221X1 U5660 ( .IN1(n30882), .IN2(n357), .IN3(n30890), .IN4(n400), .IN5(
        n5703), .Q(n5698) );
  OA22X1 U5661 ( .IN1(n30898), .IN2(n443), .IN3(n30906), .IN4(n486), .Q(n5703)
         );
  OA221X1 U5662 ( .IN1(n30850), .IN2(n529), .IN3(n30858), .IN4(n572), .IN5(
        n5704), .Q(n5697) );
  OA22X1 U5663 ( .IN1(n30866), .IN2(n615), .IN3(n30874), .IN4(n658), .Q(n5704)
         );
  NAND4X0 U5664 ( .IN1(n5705), .IN2(n5706), .IN3(n5707), .IN4(n5708), .QN(
        n5676) );
  OA221X1 U5665 ( .IN1(n30818), .IN2(n13), .IN3(n30826), .IN4(n56), .IN5(n5709), .Q(n5708) );
  OA22X1 U5666 ( .IN1(n30834), .IN2(n99), .IN3(n30842), .IN4(n142), .Q(n5709)
         );
  OA221X1 U5667 ( .IN1(n30786), .IN2(n185), .IN3(n30794), .IN4(n228), .IN5(
        n5710), .Q(n5707) );
  OA22X1 U5668 ( .IN1(n30802), .IN2(n271), .IN3(n30810), .IN4(n314), .Q(n5710)
         );
  OA221X1 U5669 ( .IN1(n30754), .IN2(n357), .IN3(n30762), .IN4(n400), .IN5(
        n5711), .Q(n5706) );
  OA22X1 U5670 ( .IN1(n30770), .IN2(n443), .IN3(n30778), .IN4(n486), .Q(n5711)
         );
  OA221X1 U5671 ( .IN1(n30722), .IN2(n529), .IN3(n30730), .IN4(n572), .IN5(
        n5712), .Q(n5705) );
  OA22X1 U5672 ( .IN1(n30738), .IN2(n615), .IN3(n30746), .IN4(n658), .Q(n5712)
         );
  OR4X1 U5673 ( .IN1(n5713), .IN2(n5714), .IN3(n5715), .IN4(n5716), .Q(n2179)
         );
  AO221X1 U5674 ( .IN1(n2157), .IN2(n5717), .IN3(n2159), .IN4(n5718), .IN5(
        n5719), .Q(n5716) );
  AO22X1 U5675 ( .IN1(n2162), .IN2(n5720), .IN3(n2164), .IN4(n5721), .Q(n5719)
         );
  NAND4X0 U5676 ( .IN1(n5722), .IN2(n5723), .IN3(n5724), .IN4(n5725), .QN(
        n5721) );
  OA221X1 U5677 ( .IN1(n30689), .IN2(n12), .IN3(n30697), .IN4(n55), .IN5(n5726), .Q(n5725) );
  OA22X1 U5678 ( .IN1(n30705), .IN2(n98), .IN3(n30713), .IN4(n141), .Q(n5726)
         );
  OA221X1 U5679 ( .IN1(n30657), .IN2(n184), .IN3(n30665), .IN4(n227), .IN5(
        n5727), .Q(n5724) );
  OA22X1 U5680 ( .IN1(n30673), .IN2(n270), .IN3(n30681), .IN4(n313), .Q(n5727)
         );
  OA221X1 U5681 ( .IN1(n30625), .IN2(n356), .IN3(n30633), .IN4(n399), .IN5(
        n5728), .Q(n5723) );
  OA22X1 U5682 ( .IN1(n30641), .IN2(n442), .IN3(n30649), .IN4(n485), .Q(n5728)
         );
  OA221X1 U5683 ( .IN1(n30593), .IN2(n528), .IN3(n30601), .IN4(n571), .IN5(
        n5729), .Q(n5722) );
  OA22X1 U5684 ( .IN1(n30609), .IN2(n614), .IN3(n30617), .IN4(n657), .Q(n5729)
         );
  NAND4X0 U5685 ( .IN1(n5730), .IN2(n5731), .IN3(n5732), .IN4(n5733), .QN(
        n5720) );
  OA221X1 U5686 ( .IN1(n30561), .IN2(n12), .IN3(n30569), .IN4(n55), .IN5(n5734), .Q(n5733) );
  OA22X1 U5687 ( .IN1(n30577), .IN2(n98), .IN3(n30585), .IN4(n141), .Q(n5734)
         );
  OA221X1 U5688 ( .IN1(n30529), .IN2(n184), .IN3(n30537), .IN4(n227), .IN5(
        n5735), .Q(n5732) );
  OA22X1 U5689 ( .IN1(n30545), .IN2(n270), .IN3(n30553), .IN4(n313), .Q(n5735)
         );
  OA221X1 U5690 ( .IN1(n30497), .IN2(n356), .IN3(n30505), .IN4(n399), .IN5(
        n5736), .Q(n5731) );
  OA22X1 U5691 ( .IN1(n30513), .IN2(n442), .IN3(n30521), .IN4(n485), .Q(n5736)
         );
  OA221X1 U5692 ( .IN1(n30465), .IN2(n528), .IN3(n30473), .IN4(n571), .IN5(
        n5737), .Q(n5730) );
  OA22X1 U5693 ( .IN1(n30481), .IN2(n614), .IN3(n30489), .IN4(n657), .Q(n5737)
         );
  NAND4X0 U5694 ( .IN1(n5738), .IN2(n5739), .IN3(n5740), .IN4(n5741), .QN(
        n5718) );
  OA221X1 U5695 ( .IN1(n30433), .IN2(n12), .IN3(n30441), .IN4(n55), .IN5(n5742), .Q(n5741) );
  OA22X1 U5696 ( .IN1(n30449), .IN2(n98), .IN3(n30457), .IN4(n141), .Q(n5742)
         );
  OA221X1 U5697 ( .IN1(n30401), .IN2(n184), .IN3(n30409), .IN4(n227), .IN5(
        n5743), .Q(n5740) );
  OA22X1 U5698 ( .IN1(n30417), .IN2(n270), .IN3(n30425), .IN4(n313), .Q(n5743)
         );
  OA221X1 U5699 ( .IN1(n30369), .IN2(n356), .IN3(n30377), .IN4(n399), .IN5(
        n5744), .Q(n5739) );
  OA22X1 U5700 ( .IN1(n30385), .IN2(n442), .IN3(n30393), .IN4(n485), .Q(n5744)
         );
  OA221X1 U5701 ( .IN1(n30337), .IN2(n528), .IN3(n30345), .IN4(n571), .IN5(
        n5745), .Q(n5738) );
  OA22X1 U5702 ( .IN1(n30353), .IN2(n614), .IN3(n30361), .IN4(n657), .Q(n5745)
         );
  NAND4X0 U5703 ( .IN1(n5746), .IN2(n5747), .IN3(n5748), .IN4(n5749), .QN(
        n5717) );
  OA221X1 U5704 ( .IN1(n30305), .IN2(n12), .IN3(n30313), .IN4(n55), .IN5(n5750), .Q(n5749) );
  OA22X1 U5705 ( .IN1(n30321), .IN2(n98), .IN3(n30329), .IN4(n141), .Q(n5750)
         );
  OA221X1 U5706 ( .IN1(n30273), .IN2(n184), .IN3(n30281), .IN4(n227), .IN5(
        n5751), .Q(n5748) );
  OA22X1 U5707 ( .IN1(n30289), .IN2(n270), .IN3(n30297), .IN4(n313), .Q(n5751)
         );
  OA221X1 U5708 ( .IN1(n30241), .IN2(n356), .IN3(n30249), .IN4(n399), .IN5(
        n5752), .Q(n5747) );
  OA22X1 U5709 ( .IN1(n30257), .IN2(n442), .IN3(n30265), .IN4(n485), .Q(n5752)
         );
  OA221X1 U5710 ( .IN1(n30209), .IN2(n528), .IN3(n30217), .IN4(n571), .IN5(
        n5753), .Q(n5746) );
  OA22X1 U5711 ( .IN1(n30225), .IN2(n614), .IN3(n30233), .IN4(n657), .Q(n5753)
         );
  AO221X1 U5712 ( .IN1(n2246), .IN2(n5754), .IN3(n2248), .IN4(n5755), .IN5(
        n5756), .Q(n5715) );
  AO22X1 U5713 ( .IN1(n2251), .IN2(n5757), .IN3(n2253), .IN4(n5758), .Q(n5756)
         );
  NAND4X0 U5714 ( .IN1(n5759), .IN2(n5760), .IN3(n5761), .IN4(n5762), .QN(
        n5758) );
  OA221X1 U5715 ( .IN1(n30177), .IN2(n12), .IN3(n30185), .IN4(n55), .IN5(n5763), .Q(n5762) );
  OA22X1 U5716 ( .IN1(n30193), .IN2(n98), .IN3(n30201), .IN4(n141), .Q(n5763)
         );
  OA221X1 U5717 ( .IN1(n30145), .IN2(n184), .IN3(n30153), .IN4(n227), .IN5(
        n5764), .Q(n5761) );
  OA22X1 U5718 ( .IN1(n30161), .IN2(n270), .IN3(n30169), .IN4(n313), .Q(n5764)
         );
  OA221X1 U5719 ( .IN1(n30113), .IN2(n356), .IN3(n30121), .IN4(n399), .IN5(
        n5765), .Q(n5760) );
  OA22X1 U5720 ( .IN1(n30129), .IN2(n442), .IN3(n30137), .IN4(n485), .Q(n5765)
         );
  OA221X1 U5721 ( .IN1(n30081), .IN2(n528), .IN3(n30089), .IN4(n571), .IN5(
        n5766), .Q(n5759) );
  OA22X1 U5722 ( .IN1(n30097), .IN2(n614), .IN3(n30105), .IN4(n657), .Q(n5766)
         );
  NAND4X0 U5723 ( .IN1(n5767), .IN2(n5768), .IN3(n5769), .IN4(n5770), .QN(
        n5757) );
  OA221X1 U5724 ( .IN1(n30049), .IN2(n12), .IN3(n30057), .IN4(n55), .IN5(n5771), .Q(n5770) );
  OA22X1 U5725 ( .IN1(n30065), .IN2(n98), .IN3(n30073), .IN4(n141), .Q(n5771)
         );
  OA221X1 U5726 ( .IN1(n30017), .IN2(n184), .IN3(n30025), .IN4(n227), .IN5(
        n5772), .Q(n5769) );
  OA22X1 U5727 ( .IN1(n30033), .IN2(n270), .IN3(n30041), .IN4(n313), .Q(n5772)
         );
  OA221X1 U5728 ( .IN1(n29985), .IN2(n356), .IN3(n29993), .IN4(n399), .IN5(
        n5773), .Q(n5768) );
  OA22X1 U5729 ( .IN1(n30001), .IN2(n442), .IN3(n30009), .IN4(n485), .Q(n5773)
         );
  OA221X1 U5730 ( .IN1(n29953), .IN2(n528), .IN3(n29961), .IN4(n571), .IN5(
        n5774), .Q(n5767) );
  OA22X1 U5731 ( .IN1(n29969), .IN2(n614), .IN3(n29977), .IN4(n657), .Q(n5774)
         );
  NAND4X0 U5732 ( .IN1(n5775), .IN2(n5776), .IN3(n5777), .IN4(n5778), .QN(
        n5755) );
  OA221X1 U5733 ( .IN1(n29921), .IN2(n12), .IN3(n29929), .IN4(n55), .IN5(n5779), .Q(n5778) );
  OA22X1 U5734 ( .IN1(n29937), .IN2(n98), .IN3(n29945), .IN4(n141), .Q(n5779)
         );
  OA221X1 U5735 ( .IN1(n29889), .IN2(n184), .IN3(n29897), .IN4(n227), .IN5(
        n5780), .Q(n5777) );
  OA22X1 U5736 ( .IN1(n29905), .IN2(n270), .IN3(n29913), .IN4(n313), .Q(n5780)
         );
  OA221X1 U5737 ( .IN1(n29857), .IN2(n356), .IN3(n29865), .IN4(n399), .IN5(
        n5781), .Q(n5776) );
  OA22X1 U5738 ( .IN1(n29873), .IN2(n442), .IN3(n29881), .IN4(n485), .Q(n5781)
         );
  OA221X1 U5739 ( .IN1(n29825), .IN2(n528), .IN3(n29833), .IN4(n571), .IN5(
        n5782), .Q(n5775) );
  OA22X1 U5740 ( .IN1(n29841), .IN2(n614), .IN3(n29849), .IN4(n657), .Q(n5782)
         );
  NAND4X0 U5741 ( .IN1(n5783), .IN2(n5784), .IN3(n5785), .IN4(n5786), .QN(
        n5754) );
  OA221X1 U5742 ( .IN1(n29793), .IN2(n12), .IN3(n29801), .IN4(n55), .IN5(n5787), .Q(n5786) );
  OA22X1 U5743 ( .IN1(n29809), .IN2(n98), .IN3(n29817), .IN4(n141), .Q(n5787)
         );
  OA221X1 U5744 ( .IN1(n29761), .IN2(n184), .IN3(n29769), .IN4(n227), .IN5(
        n5788), .Q(n5785) );
  OA22X1 U5745 ( .IN1(n29777), .IN2(n270), .IN3(n29785), .IN4(n313), .Q(n5788)
         );
  OA221X1 U5746 ( .IN1(n29729), .IN2(n356), .IN3(n29737), .IN4(n399), .IN5(
        n5789), .Q(n5784) );
  OA22X1 U5747 ( .IN1(n29745), .IN2(n442), .IN3(n29753), .IN4(n485), .Q(n5789)
         );
  OA221X1 U5748 ( .IN1(n29697), .IN2(n528), .IN3(n29705), .IN4(n571), .IN5(
        n5790), .Q(n5783) );
  OA22X1 U5749 ( .IN1(n29713), .IN2(n614), .IN3(n29721), .IN4(n657), .Q(n5790)
         );
  AO221X1 U5750 ( .IN1(n2287), .IN2(n5791), .IN3(n2289), .IN4(n5792), .IN5(
        n5793), .Q(n5714) );
  AO22X1 U5751 ( .IN1(n2292), .IN2(n5794), .IN3(n2294), .IN4(n5795), .Q(n5793)
         );
  NAND4X0 U5752 ( .IN1(n5796), .IN2(n5797), .IN3(n5798), .IN4(n5799), .QN(
        n5795) );
  OA221X1 U5753 ( .IN1(n31713), .IN2(n12), .IN3(n31721), .IN4(n55), .IN5(n5800), .Q(n5799) );
  OA22X1 U5754 ( .IN1(n31729), .IN2(n98), .IN3(n31737), .IN4(n141), .Q(n5800)
         );
  OA221X1 U5755 ( .IN1(n31681), .IN2(n184), .IN3(n31689), .IN4(n227), .IN5(
        n5801), .Q(n5798) );
  OA22X1 U5756 ( .IN1(n31697), .IN2(n270), .IN3(n31705), .IN4(n313), .Q(n5801)
         );
  OA221X1 U5757 ( .IN1(n31649), .IN2(n356), .IN3(n31657), .IN4(n399), .IN5(
        n5802), .Q(n5797) );
  OA22X1 U5758 ( .IN1(n31665), .IN2(n442), .IN3(n31673), .IN4(n485), .Q(n5802)
         );
  OA221X1 U5759 ( .IN1(n31617), .IN2(n528), .IN3(n31625), .IN4(n571), .IN5(
        n5803), .Q(n5796) );
  OA22X1 U5760 ( .IN1(n31633), .IN2(n614), .IN3(n31641), .IN4(n657), .Q(n5803)
         );
  NAND4X0 U5761 ( .IN1(n5804), .IN2(n5805), .IN3(n5806), .IN4(n5807), .QN(
        n5794) );
  OA221X1 U5762 ( .IN1(n31585), .IN2(n12), .IN3(n31593), .IN4(n55), .IN5(n5808), .Q(n5807) );
  OA22X1 U5763 ( .IN1(n31601), .IN2(n98), .IN3(n31609), .IN4(n141), .Q(n5808)
         );
  OA221X1 U5764 ( .IN1(n31553), .IN2(n184), .IN3(n31561), .IN4(n227), .IN5(
        n5809), .Q(n5806) );
  OA22X1 U5765 ( .IN1(n31569), .IN2(n270), .IN3(n31577), .IN4(n313), .Q(n5809)
         );
  OA221X1 U5766 ( .IN1(n31521), .IN2(n356), .IN3(n31529), .IN4(n399), .IN5(
        n5810), .Q(n5805) );
  OA22X1 U5767 ( .IN1(n31537), .IN2(n442), .IN3(n31545), .IN4(n485), .Q(n5810)
         );
  OA221X1 U5768 ( .IN1(n31489), .IN2(n528), .IN3(n31497), .IN4(n571), .IN5(
        n5811), .Q(n5804) );
  OA22X1 U5769 ( .IN1(n31505), .IN2(n614), .IN3(n31513), .IN4(n657), .Q(n5811)
         );
  NAND4X0 U5770 ( .IN1(n5812), .IN2(n5813), .IN3(n5814), .IN4(n5815), .QN(
        n5792) );
  OA221X1 U5771 ( .IN1(n31457), .IN2(n12), .IN3(n31465), .IN4(n55), .IN5(n5816), .Q(n5815) );
  OA22X1 U5772 ( .IN1(n31473), .IN2(n98), .IN3(n31481), .IN4(n141), .Q(n5816)
         );
  OA221X1 U5773 ( .IN1(n31425), .IN2(n184), .IN3(n31433), .IN4(n227), .IN5(
        n5817), .Q(n5814) );
  OA22X1 U5774 ( .IN1(n31441), .IN2(n270), .IN3(n31449), .IN4(n313), .Q(n5817)
         );
  OA221X1 U5775 ( .IN1(n31393), .IN2(n356), .IN3(n31401), .IN4(n399), .IN5(
        n5818), .Q(n5813) );
  OA22X1 U5776 ( .IN1(n31409), .IN2(n442), .IN3(n31417), .IN4(n485), .Q(n5818)
         );
  OA221X1 U5777 ( .IN1(n31361), .IN2(n528), .IN3(n31369), .IN4(n571), .IN5(
        n5819), .Q(n5812) );
  OA22X1 U5778 ( .IN1(n31377), .IN2(n614), .IN3(n31385), .IN4(n657), .Q(n5819)
         );
  NAND4X0 U5779 ( .IN1(n5820), .IN2(n5821), .IN3(n5822), .IN4(n5823), .QN(
        n5791) );
  OA221X1 U5780 ( .IN1(n31329), .IN2(n12), .IN3(n31337), .IN4(n55), .IN5(n5824), .Q(n5823) );
  OA22X1 U5781 ( .IN1(n31345), .IN2(n98), .IN3(n31353), .IN4(n141), .Q(n5824)
         );
  OA221X1 U5782 ( .IN1(n31297), .IN2(n184), .IN3(n31305), .IN4(n227), .IN5(
        n5825), .Q(n5822) );
  OA22X1 U5783 ( .IN1(n31313), .IN2(n270), .IN3(n31321), .IN4(n313), .Q(n5825)
         );
  OA221X1 U5784 ( .IN1(n31265), .IN2(n356), .IN3(n31273), .IN4(n399), .IN5(
        n5826), .Q(n5821) );
  OA22X1 U5785 ( .IN1(n31281), .IN2(n442), .IN3(n31289), .IN4(n485), .Q(n5826)
         );
  OA221X1 U5786 ( .IN1(n31233), .IN2(n528), .IN3(n31241), .IN4(n571), .IN5(
        n5827), .Q(n5820) );
  OA22X1 U5787 ( .IN1(n31249), .IN2(n614), .IN3(n31257), .IN4(n657), .Q(n5827)
         );
  AO221X1 U5788 ( .IN1(n2328), .IN2(n5828), .IN3(n2330), .IN4(n5829), .IN5(
        n5830), .Q(n5713) );
  AO22X1 U5789 ( .IN1(n2333), .IN2(n5831), .IN3(n2335), .IN4(n5832), .Q(n5830)
         );
  NAND4X0 U5790 ( .IN1(n5833), .IN2(n5834), .IN3(n5835), .IN4(n5836), .QN(
        n5832) );
  OA221X1 U5791 ( .IN1(n31201), .IN2(n11), .IN3(n31209), .IN4(n54), .IN5(n5837), .Q(n5836) );
  OA22X1 U5792 ( .IN1(n31217), .IN2(n97), .IN3(n31225), .IN4(n140), .Q(n5837)
         );
  OA221X1 U5793 ( .IN1(n31169), .IN2(n183), .IN3(n31177), .IN4(n226), .IN5(
        n5838), .Q(n5835) );
  OA22X1 U5794 ( .IN1(n31185), .IN2(n269), .IN3(n31193), .IN4(n312), .Q(n5838)
         );
  OA221X1 U5795 ( .IN1(n31137), .IN2(n355), .IN3(n31145), .IN4(n398), .IN5(
        n5839), .Q(n5834) );
  OA22X1 U5796 ( .IN1(n31153), .IN2(n441), .IN3(n31161), .IN4(n484), .Q(n5839)
         );
  OA221X1 U5797 ( .IN1(n31105), .IN2(n527), .IN3(n31113), .IN4(n570), .IN5(
        n5840), .Q(n5833) );
  OA22X1 U5798 ( .IN1(n31121), .IN2(n613), .IN3(n31129), .IN4(n656), .Q(n5840)
         );
  NAND4X0 U5799 ( .IN1(n5841), .IN2(n5842), .IN3(n5843), .IN4(n5844), .QN(
        n5831) );
  OA221X1 U5800 ( .IN1(n31073), .IN2(n11), .IN3(n31081), .IN4(n54), .IN5(n5845), .Q(n5844) );
  OA22X1 U5801 ( .IN1(n31089), .IN2(n97), .IN3(n31097), .IN4(n140), .Q(n5845)
         );
  OA221X1 U5802 ( .IN1(n31041), .IN2(n183), .IN3(n31049), .IN4(n226), .IN5(
        n5846), .Q(n5843) );
  OA22X1 U5803 ( .IN1(n31057), .IN2(n269), .IN3(n31065), .IN4(n312), .Q(n5846)
         );
  OA221X1 U5804 ( .IN1(n31009), .IN2(n355), .IN3(n31017), .IN4(n398), .IN5(
        n5847), .Q(n5842) );
  OA22X1 U5805 ( .IN1(n31025), .IN2(n441), .IN3(n31033), .IN4(n484), .Q(n5847)
         );
  OA221X1 U5806 ( .IN1(n30977), .IN2(n527), .IN3(n30985), .IN4(n570), .IN5(
        n5848), .Q(n5841) );
  OA22X1 U5807 ( .IN1(n30993), .IN2(n613), .IN3(n31001), .IN4(n656), .Q(n5848)
         );
  NAND4X0 U5808 ( .IN1(n5849), .IN2(n5850), .IN3(n5851), .IN4(n5852), .QN(
        n5829) );
  OA221X1 U5809 ( .IN1(n30945), .IN2(n11), .IN3(n30953), .IN4(n54), .IN5(n5853), .Q(n5852) );
  OA22X1 U5810 ( .IN1(n30961), .IN2(n97), .IN3(n30969), .IN4(n140), .Q(n5853)
         );
  OA221X1 U5811 ( .IN1(n30913), .IN2(n183), .IN3(n30921), .IN4(n226), .IN5(
        n5854), .Q(n5851) );
  OA22X1 U5812 ( .IN1(n30929), .IN2(n269), .IN3(n30937), .IN4(n312), .Q(n5854)
         );
  OA221X1 U5813 ( .IN1(n30881), .IN2(n355), .IN3(n30889), .IN4(n398), .IN5(
        n5855), .Q(n5850) );
  OA22X1 U5814 ( .IN1(n30897), .IN2(n441), .IN3(n30905), .IN4(n484), .Q(n5855)
         );
  OA221X1 U5815 ( .IN1(n30849), .IN2(n527), .IN3(n30857), .IN4(n570), .IN5(
        n5856), .Q(n5849) );
  OA22X1 U5816 ( .IN1(n30865), .IN2(n613), .IN3(n30873), .IN4(n656), .Q(n5856)
         );
  NAND4X0 U5817 ( .IN1(n5857), .IN2(n5858), .IN3(n5859), .IN4(n5860), .QN(
        n5828) );
  OA221X1 U5818 ( .IN1(n30817), .IN2(n11), .IN3(n30825), .IN4(n54), .IN5(n5861), .Q(n5860) );
  OA22X1 U5819 ( .IN1(n30833), .IN2(n97), .IN3(n30841), .IN4(n140), .Q(n5861)
         );
  OA221X1 U5820 ( .IN1(n30785), .IN2(n183), .IN3(n30793), .IN4(n226), .IN5(
        n5862), .Q(n5859) );
  OA22X1 U5821 ( .IN1(n30801), .IN2(n269), .IN3(n30809), .IN4(n312), .Q(n5862)
         );
  OA221X1 U5822 ( .IN1(n30753), .IN2(n355), .IN3(n30761), .IN4(n398), .IN5(
        n5863), .Q(n5858) );
  OA22X1 U5823 ( .IN1(n30769), .IN2(n441), .IN3(n30777), .IN4(n484), .Q(n5863)
         );
  OA221X1 U5824 ( .IN1(n30721), .IN2(n527), .IN3(n30729), .IN4(n570), .IN5(
        n5864), .Q(n5857) );
  OA22X1 U5825 ( .IN1(n30737), .IN2(n613), .IN3(n30745), .IN4(n656), .Q(n5864)
         );
  OR4X1 U5826 ( .IN1(n5865), .IN2(n5866), .IN3(n5867), .IN4(n5868), .Q(n2178)
         );
  AO221X1 U5827 ( .IN1(n2157), .IN2(n5869), .IN3(n2159), .IN4(n5870), .IN5(
        n5871), .Q(n5868) );
  AO22X1 U5828 ( .IN1(n2162), .IN2(n5872), .IN3(n2164), .IN4(n5873), .Q(n5871)
         );
  NAND4X0 U5829 ( .IN1(n5874), .IN2(n5875), .IN3(n5876), .IN4(n5877), .QN(
        n5873) );
  OA221X1 U5830 ( .IN1(n28648), .IN2(n11), .IN3(n28656), .IN4(n54), .IN5(n5878), .Q(n5877) );
  OA22X1 U5831 ( .IN1(n28664), .IN2(n97), .IN3(n28672), .IN4(n140), .Q(n5878)
         );
  OA221X1 U5832 ( .IN1(n28616), .IN2(n183), .IN3(n28624), .IN4(n226), .IN5(
        n5879), .Q(n5876) );
  OA22X1 U5833 ( .IN1(n28632), .IN2(n269), .IN3(n28640), .IN4(n312), .Q(n5879)
         );
  OA221X1 U5834 ( .IN1(n28584), .IN2(n355), .IN3(n28592), .IN4(n398), .IN5(
        n5880), .Q(n5875) );
  OA22X1 U5835 ( .IN1(n28600), .IN2(n441), .IN3(n28608), .IN4(n484), .Q(n5880)
         );
  OA221X1 U5836 ( .IN1(n28552), .IN2(n527), .IN3(n28560), .IN4(n570), .IN5(
        n5881), .Q(n5874) );
  OA22X1 U5837 ( .IN1(n28568), .IN2(n613), .IN3(n28576), .IN4(n656), .Q(n5881)
         );
  NAND4X0 U5838 ( .IN1(n5882), .IN2(n5883), .IN3(n5884), .IN4(n5885), .QN(
        n5872) );
  OA221X1 U5839 ( .IN1(n28520), .IN2(n11), .IN3(n28528), .IN4(n54), .IN5(n5886), .Q(n5885) );
  OA22X1 U5840 ( .IN1(n28536), .IN2(n97), .IN3(n28544), .IN4(n140), .Q(n5886)
         );
  OA221X1 U5841 ( .IN1(n28488), .IN2(n183), .IN3(n28496), .IN4(n226), .IN5(
        n5887), .Q(n5884) );
  OA22X1 U5842 ( .IN1(n28504), .IN2(n269), .IN3(n28512), .IN4(n312), .Q(n5887)
         );
  OA221X1 U5843 ( .IN1(n28456), .IN2(n355), .IN3(n28464), .IN4(n398), .IN5(
        n5888), .Q(n5883) );
  OA22X1 U5844 ( .IN1(n28472), .IN2(n441), .IN3(n28480), .IN4(n484), .Q(n5888)
         );
  OA221X1 U5845 ( .IN1(n28424), .IN2(n527), .IN3(n28432), .IN4(n570), .IN5(
        n5889), .Q(n5882) );
  OA22X1 U5846 ( .IN1(n28440), .IN2(n613), .IN3(n28448), .IN4(n656), .Q(n5889)
         );
  NAND4X0 U5847 ( .IN1(n5890), .IN2(n5891), .IN3(n5892), .IN4(n5893), .QN(
        n5870) );
  OA221X1 U5848 ( .IN1(n28392), .IN2(n11), .IN3(n28400), .IN4(n54), .IN5(n5894), .Q(n5893) );
  OA22X1 U5849 ( .IN1(n28408), .IN2(n97), .IN3(n28416), .IN4(n140), .Q(n5894)
         );
  OA221X1 U5850 ( .IN1(n28360), .IN2(n183), .IN3(n28368), .IN4(n226), .IN5(
        n5895), .Q(n5892) );
  OA22X1 U5851 ( .IN1(n28376), .IN2(n269), .IN3(n28384), .IN4(n312), .Q(n5895)
         );
  OA221X1 U5852 ( .IN1(n28328), .IN2(n355), .IN3(n28336), .IN4(n398), .IN5(
        n5896), .Q(n5891) );
  OA22X1 U5853 ( .IN1(n28344), .IN2(n441), .IN3(n28352), .IN4(n484), .Q(n5896)
         );
  OA221X1 U5854 ( .IN1(n28296), .IN2(n527), .IN3(n28304), .IN4(n570), .IN5(
        n5897), .Q(n5890) );
  OA22X1 U5855 ( .IN1(n28312), .IN2(n613), .IN3(n28320), .IN4(n656), .Q(n5897)
         );
  NAND4X0 U5856 ( .IN1(n5898), .IN2(n5899), .IN3(n5900), .IN4(n5901), .QN(
        n5869) );
  OA221X1 U5857 ( .IN1(n28264), .IN2(n11), .IN3(n28272), .IN4(n54), .IN5(n5902), .Q(n5901) );
  OA22X1 U5858 ( .IN1(n28280), .IN2(n97), .IN3(n28288), .IN4(n140), .Q(n5902)
         );
  OA221X1 U5859 ( .IN1(n28232), .IN2(n183), .IN3(n28240), .IN4(n226), .IN5(
        n5903), .Q(n5900) );
  OA22X1 U5860 ( .IN1(n28248), .IN2(n269), .IN3(n28256), .IN4(n312), .Q(n5903)
         );
  OA221X1 U5861 ( .IN1(n28200), .IN2(n355), .IN3(n28208), .IN4(n398), .IN5(
        n5904), .Q(n5899) );
  OA22X1 U5862 ( .IN1(n28216), .IN2(n441), .IN3(n28224), .IN4(n484), .Q(n5904)
         );
  OA221X1 U5863 ( .IN1(n28168), .IN2(n527), .IN3(n28176), .IN4(n570), .IN5(
        n5905), .Q(n5898) );
  OA22X1 U5864 ( .IN1(n28184), .IN2(n613), .IN3(n28192), .IN4(n656), .Q(n5905)
         );
  AO221X1 U5865 ( .IN1(n2246), .IN2(n5906), .IN3(n2248), .IN4(n5907), .IN5(
        n5908), .Q(n5867) );
  AO22X1 U5866 ( .IN1(n2251), .IN2(n5909), .IN3(n2253), .IN4(n5910), .Q(n5908)
         );
  NAND4X0 U5867 ( .IN1(n5911), .IN2(n5912), .IN3(n5913), .IN4(n5914), .QN(
        n5910) );
  OA221X1 U5868 ( .IN1(n28136), .IN2(n11), .IN3(n28144), .IN4(n54), .IN5(n5915), .Q(n5914) );
  OA22X1 U5869 ( .IN1(n28152), .IN2(n97), .IN3(n28160), .IN4(n140), .Q(n5915)
         );
  OA221X1 U5870 ( .IN1(n28104), .IN2(n183), .IN3(n28112), .IN4(n226), .IN5(
        n5916), .Q(n5913) );
  OA22X1 U5871 ( .IN1(n28120), .IN2(n269), .IN3(n28128), .IN4(n312), .Q(n5916)
         );
  OA221X1 U5872 ( .IN1(n28072), .IN2(n355), .IN3(n28080), .IN4(n398), .IN5(
        n5917), .Q(n5912) );
  OA22X1 U5873 ( .IN1(n28088), .IN2(n441), .IN3(n28096), .IN4(n484), .Q(n5917)
         );
  OA221X1 U5874 ( .IN1(n28040), .IN2(n527), .IN3(n28048), .IN4(n570), .IN5(
        n5918), .Q(n5911) );
  OA22X1 U5875 ( .IN1(n28056), .IN2(n613), .IN3(n28064), .IN4(n656), .Q(n5918)
         );
  NAND4X0 U5876 ( .IN1(n5919), .IN2(n5920), .IN3(n5921), .IN4(n5922), .QN(
        n5909) );
  OA221X1 U5877 ( .IN1(n28008), .IN2(n11), .IN3(n28016), .IN4(n54), .IN5(n5923), .Q(n5922) );
  OA22X1 U5878 ( .IN1(n28024), .IN2(n97), .IN3(n28032), .IN4(n140), .Q(n5923)
         );
  OA221X1 U5879 ( .IN1(n27976), .IN2(n183), .IN3(n27984), .IN4(n226), .IN5(
        n5924), .Q(n5921) );
  OA22X1 U5880 ( .IN1(n27992), .IN2(n269), .IN3(n28000), .IN4(n312), .Q(n5924)
         );
  OA221X1 U5881 ( .IN1(n27944), .IN2(n355), .IN3(n27952), .IN4(n398), .IN5(
        n5925), .Q(n5920) );
  OA22X1 U5882 ( .IN1(n27960), .IN2(n441), .IN3(n27968), .IN4(n484), .Q(n5925)
         );
  OA221X1 U5883 ( .IN1(n27912), .IN2(n527), .IN3(n27920), .IN4(n570), .IN5(
        n5926), .Q(n5919) );
  OA22X1 U5884 ( .IN1(n27928), .IN2(n613), .IN3(n27936), .IN4(n656), .Q(n5926)
         );
  NAND4X0 U5885 ( .IN1(n5927), .IN2(n5928), .IN3(n5929), .IN4(n5930), .QN(
        n5907) );
  OA221X1 U5886 ( .IN1(n27880), .IN2(n11), .IN3(n27888), .IN4(n54), .IN5(n5931), .Q(n5930) );
  OA22X1 U5887 ( .IN1(n27896), .IN2(n97), .IN3(n27904), .IN4(n140), .Q(n5931)
         );
  OA221X1 U5888 ( .IN1(n27848), .IN2(n183), .IN3(n27856), .IN4(n226), .IN5(
        n5932), .Q(n5929) );
  OA22X1 U5889 ( .IN1(n27864), .IN2(n269), .IN3(n27872), .IN4(n312), .Q(n5932)
         );
  OA221X1 U5890 ( .IN1(n27816), .IN2(n355), .IN3(n27824), .IN4(n398), .IN5(
        n5933), .Q(n5928) );
  OA22X1 U5891 ( .IN1(n27832), .IN2(n441), .IN3(n27840), .IN4(n484), .Q(n5933)
         );
  OA221X1 U5892 ( .IN1(n27784), .IN2(n527), .IN3(n27792), .IN4(n570), .IN5(
        n5934), .Q(n5927) );
  OA22X1 U5893 ( .IN1(n27800), .IN2(n613), .IN3(n27808), .IN4(n656), .Q(n5934)
         );
  NAND4X0 U5894 ( .IN1(n5935), .IN2(n5936), .IN3(n5937), .IN4(n5938), .QN(
        n5906) );
  OA221X1 U5895 ( .IN1(n27752), .IN2(n11), .IN3(n27760), .IN4(n54), .IN5(n5939), .Q(n5938) );
  OA22X1 U5896 ( .IN1(n27768), .IN2(n97), .IN3(n27776), .IN4(n140), .Q(n5939)
         );
  OA221X1 U5897 ( .IN1(n27720), .IN2(n183), .IN3(n27728), .IN4(n226), .IN5(
        n5940), .Q(n5937) );
  OA22X1 U5898 ( .IN1(n27736), .IN2(n269), .IN3(n27744), .IN4(n312), .Q(n5940)
         );
  OA221X1 U5899 ( .IN1(n27688), .IN2(n355), .IN3(n27696), .IN4(n398), .IN5(
        n5941), .Q(n5936) );
  OA22X1 U5900 ( .IN1(n27704), .IN2(n441), .IN3(n27712), .IN4(n484), .Q(n5941)
         );
  OA221X1 U5901 ( .IN1(n27656), .IN2(n527), .IN3(n27664), .IN4(n570), .IN5(
        n5942), .Q(n5935) );
  OA22X1 U5902 ( .IN1(n27672), .IN2(n613), .IN3(n27680), .IN4(n656), .Q(n5942)
         );
  AO221X1 U5903 ( .IN1(n2287), .IN2(n5943), .IN3(n2289), .IN4(n5944), .IN5(
        n5945), .Q(n5866) );
  AO22X1 U5904 ( .IN1(n2292), .IN2(n5946), .IN3(n2294), .IN4(n5947), .Q(n5945)
         );
  NAND4X0 U5905 ( .IN1(n5948), .IN2(n5949), .IN3(n5950), .IN4(n5951), .QN(
        n5947) );
  OA221X1 U5906 ( .IN1(n29672), .IN2(n10), .IN3(n29680), .IN4(n53), .IN5(n5952), .Q(n5951) );
  OA22X1 U5907 ( .IN1(n29688), .IN2(n96), .IN3(n29696), .IN4(n139), .Q(n5952)
         );
  OA221X1 U5908 ( .IN1(n29640), .IN2(n182), .IN3(n29648), .IN4(n225), .IN5(
        n5953), .Q(n5950) );
  OA22X1 U5909 ( .IN1(n29656), .IN2(n268), .IN3(n29664), .IN4(n311), .Q(n5953)
         );
  OA221X1 U5910 ( .IN1(n29608), .IN2(n354), .IN3(n29616), .IN4(n397), .IN5(
        n5954), .Q(n5949) );
  OA22X1 U5911 ( .IN1(n29624), .IN2(n440), .IN3(n29632), .IN4(n483), .Q(n5954)
         );
  OA221X1 U5912 ( .IN1(n29576), .IN2(n526), .IN3(n29584), .IN4(n569), .IN5(
        n5955), .Q(n5948) );
  OA22X1 U5913 ( .IN1(n29592), .IN2(n612), .IN3(n29600), .IN4(n655), .Q(n5955)
         );
  NAND4X0 U5914 ( .IN1(n5956), .IN2(n5957), .IN3(n5958), .IN4(n5959), .QN(
        n5946) );
  OA221X1 U5915 ( .IN1(n29544), .IN2(n10), .IN3(n29552), .IN4(n53), .IN5(n5960), .Q(n5959) );
  OA22X1 U5916 ( .IN1(n29560), .IN2(n96), .IN3(n29568), .IN4(n139), .Q(n5960)
         );
  OA221X1 U5917 ( .IN1(n29512), .IN2(n182), .IN3(n29520), .IN4(n225), .IN5(
        n5961), .Q(n5958) );
  OA22X1 U5918 ( .IN1(n29528), .IN2(n268), .IN3(n29536), .IN4(n311), .Q(n5961)
         );
  OA221X1 U5919 ( .IN1(n29480), .IN2(n354), .IN3(n29488), .IN4(n397), .IN5(
        n5962), .Q(n5957) );
  OA22X1 U5920 ( .IN1(n29496), .IN2(n440), .IN3(n29504), .IN4(n483), .Q(n5962)
         );
  OA221X1 U5921 ( .IN1(n29448), .IN2(n526), .IN3(n29456), .IN4(n569), .IN5(
        n5963), .Q(n5956) );
  OA22X1 U5922 ( .IN1(n29464), .IN2(n612), .IN3(n29472), .IN4(n655), .Q(n5963)
         );
  NAND4X0 U5923 ( .IN1(n5964), .IN2(n5965), .IN3(n5966), .IN4(n5967), .QN(
        n5944) );
  OA221X1 U5924 ( .IN1(n29416), .IN2(n10), .IN3(n29424), .IN4(n53), .IN5(n5968), .Q(n5967) );
  OA22X1 U5925 ( .IN1(n29432), .IN2(n96), .IN3(n29440), .IN4(n139), .Q(n5968)
         );
  OA221X1 U5926 ( .IN1(n29384), .IN2(n182), .IN3(n29392), .IN4(n225), .IN5(
        n5969), .Q(n5966) );
  OA22X1 U5927 ( .IN1(n29400), .IN2(n268), .IN3(n29408), .IN4(n311), .Q(n5969)
         );
  OA221X1 U5928 ( .IN1(n29352), .IN2(n354), .IN3(n29360), .IN4(n397), .IN5(
        n5970), .Q(n5965) );
  OA22X1 U5929 ( .IN1(n29368), .IN2(n440), .IN3(n29376), .IN4(n483), .Q(n5970)
         );
  OA221X1 U5930 ( .IN1(n29320), .IN2(n526), .IN3(n29328), .IN4(n569), .IN5(
        n5971), .Q(n5964) );
  OA22X1 U5931 ( .IN1(n29336), .IN2(n612), .IN3(n29344), .IN4(n655), .Q(n5971)
         );
  NAND4X0 U5932 ( .IN1(n5972), .IN2(n5973), .IN3(n5974), .IN4(n5975), .QN(
        n5943) );
  OA221X1 U5933 ( .IN1(n29288), .IN2(n10), .IN3(n29296), .IN4(n53), .IN5(n5976), .Q(n5975) );
  OA22X1 U5934 ( .IN1(n29304), .IN2(n96), .IN3(n29312), .IN4(n139), .Q(n5976)
         );
  OA221X1 U5935 ( .IN1(n29256), .IN2(n182), .IN3(n29264), .IN4(n225), .IN5(
        n5977), .Q(n5974) );
  OA22X1 U5936 ( .IN1(n29272), .IN2(n268), .IN3(n29280), .IN4(n311), .Q(n5977)
         );
  OA221X1 U5937 ( .IN1(n29224), .IN2(n354), .IN3(n29232), .IN4(n397), .IN5(
        n5978), .Q(n5973) );
  OA22X1 U5938 ( .IN1(n29240), .IN2(n440), .IN3(n29248), .IN4(n483), .Q(n5978)
         );
  OA221X1 U5939 ( .IN1(n29192), .IN2(n526), .IN3(n29200), .IN4(n569), .IN5(
        n5979), .Q(n5972) );
  OA22X1 U5940 ( .IN1(n29208), .IN2(n612), .IN3(n29216), .IN4(n655), .Q(n5979)
         );
  AO221X1 U5941 ( .IN1(n2328), .IN2(n5980), .IN3(n2330), .IN4(n5981), .IN5(
        n5982), .Q(n5865) );
  AO22X1 U5942 ( .IN1(n2333), .IN2(n5983), .IN3(n2335), .IN4(n5984), .Q(n5982)
         );
  NAND4X0 U5943 ( .IN1(n5985), .IN2(n5986), .IN3(n5987), .IN4(n5988), .QN(
        n5984) );
  OA221X1 U5944 ( .IN1(n29160), .IN2(n10), .IN3(n29168), .IN4(n53), .IN5(n5989), .Q(n5988) );
  OA22X1 U5945 ( .IN1(n29176), .IN2(n96), .IN3(n29184), .IN4(n139), .Q(n5989)
         );
  OA221X1 U5946 ( .IN1(n29128), .IN2(n182), .IN3(n29136), .IN4(n225), .IN5(
        n5990), .Q(n5987) );
  OA22X1 U5947 ( .IN1(n29144), .IN2(n268), .IN3(n29152), .IN4(n311), .Q(n5990)
         );
  OA221X1 U5948 ( .IN1(n29096), .IN2(n354), .IN3(n29104), .IN4(n397), .IN5(
        n5991), .Q(n5986) );
  OA22X1 U5949 ( .IN1(n29112), .IN2(n440), .IN3(n29120), .IN4(n483), .Q(n5991)
         );
  OA221X1 U5950 ( .IN1(n29064), .IN2(n526), .IN3(n29072), .IN4(n569), .IN5(
        n5992), .Q(n5985) );
  OA22X1 U5951 ( .IN1(n29080), .IN2(n612), .IN3(n29088), .IN4(n655), .Q(n5992)
         );
  NAND4X0 U5952 ( .IN1(n5993), .IN2(n5994), .IN3(n5995), .IN4(n5996), .QN(
        n5983) );
  OA221X1 U5953 ( .IN1(n29032), .IN2(n10), .IN3(n29040), .IN4(n53), .IN5(n5997), .Q(n5996) );
  OA22X1 U5954 ( .IN1(n29048), .IN2(n96), .IN3(n29056), .IN4(n139), .Q(n5997)
         );
  OA221X1 U5955 ( .IN1(n29000), .IN2(n182), .IN3(n29008), .IN4(n225), .IN5(
        n5998), .Q(n5995) );
  OA22X1 U5956 ( .IN1(n29016), .IN2(n268), .IN3(n29024), .IN4(n311), .Q(n5998)
         );
  OA221X1 U5957 ( .IN1(n28968), .IN2(n354), .IN3(n28976), .IN4(n397), .IN5(
        n5999), .Q(n5994) );
  OA22X1 U5958 ( .IN1(n28984), .IN2(n440), .IN3(n28992), .IN4(n483), .Q(n5999)
         );
  OA221X1 U5959 ( .IN1(n28936), .IN2(n526), .IN3(n28944), .IN4(n569), .IN5(
        n6000), .Q(n5993) );
  OA22X1 U5960 ( .IN1(n28952), .IN2(n612), .IN3(n28960), .IN4(n655), .Q(n6000)
         );
  NAND4X0 U5961 ( .IN1(n6001), .IN2(n6002), .IN3(n6003), .IN4(n6004), .QN(
        n5981) );
  OA221X1 U5962 ( .IN1(n28904), .IN2(n10), .IN3(n28912), .IN4(n53), .IN5(n6005), .Q(n6004) );
  OA22X1 U5963 ( .IN1(n28920), .IN2(n96), .IN3(n28928), .IN4(n139), .Q(n6005)
         );
  OA221X1 U5964 ( .IN1(n28872), .IN2(n182), .IN3(n28880), .IN4(n225), .IN5(
        n6006), .Q(n6003) );
  OA22X1 U5965 ( .IN1(n28888), .IN2(n268), .IN3(n28896), .IN4(n311), .Q(n6006)
         );
  OA221X1 U5966 ( .IN1(n28840), .IN2(n354), .IN3(n28848), .IN4(n397), .IN5(
        n6007), .Q(n6002) );
  OA22X1 U5967 ( .IN1(n28856), .IN2(n440), .IN3(n28864), .IN4(n483), .Q(n6007)
         );
  OA221X1 U5968 ( .IN1(n28808), .IN2(n526), .IN3(n28816), .IN4(n569), .IN5(
        n6008), .Q(n6001) );
  OA22X1 U5969 ( .IN1(n28824), .IN2(n612), .IN3(n28832), .IN4(n655), .Q(n6008)
         );
  NAND4X0 U5970 ( .IN1(n6009), .IN2(n6010), .IN3(n6011), .IN4(n6012), .QN(
        n5980) );
  OA221X1 U5971 ( .IN1(n28776), .IN2(n10), .IN3(n28784), .IN4(n53), .IN5(n6013), .Q(n6012) );
  OA22X1 U5972 ( .IN1(n28792), .IN2(n96), .IN3(n28800), .IN4(n139), .Q(n6013)
         );
  OA221X1 U5973 ( .IN1(n28744), .IN2(n182), .IN3(n28752), .IN4(n225), .IN5(
        n6014), .Q(n6011) );
  OA22X1 U5974 ( .IN1(n28760), .IN2(n268), .IN3(n28768), .IN4(n311), .Q(n6014)
         );
  OA221X1 U5975 ( .IN1(n28712), .IN2(n354), .IN3(n28720), .IN4(n397), .IN5(
        n6015), .Q(n6010) );
  OA22X1 U5976 ( .IN1(n28728), .IN2(n440), .IN3(n28736), .IN4(n483), .Q(n6015)
         );
  OA221X1 U5977 ( .IN1(n28680), .IN2(n526), .IN3(n28688), .IN4(n569), .IN5(
        n6016), .Q(n6009) );
  OA22X1 U5978 ( .IN1(n28696), .IN2(n612), .IN3(n28704), .IN4(n655), .Q(n6016)
         );
  OR4X1 U5979 ( .IN1(n6017), .IN2(n6018), .IN3(n6019), .IN4(n6020), .Q(n2177)
         );
  AO221X1 U5980 ( .IN1(n2157), .IN2(n6021), .IN3(n2159), .IN4(n6022), .IN5(
        n6023), .Q(n6020) );
  AO22X1 U5981 ( .IN1(n2162), .IN2(n6024), .IN3(n2164), .IN4(n6025), .Q(n6023)
         );
  NAND4X0 U5982 ( .IN1(n6026), .IN2(n6027), .IN3(n6028), .IN4(n6029), .QN(
        n6025) );
  OA221X1 U5983 ( .IN1(n28647), .IN2(n10), .IN3(n28655), .IN4(n53), .IN5(n6030), .Q(n6029) );
  OA22X1 U5984 ( .IN1(n28663), .IN2(n96), .IN3(n28671), .IN4(n139), .Q(n6030)
         );
  OA221X1 U5985 ( .IN1(n28615), .IN2(n182), .IN3(n28623), .IN4(n225), .IN5(
        n6031), .Q(n6028) );
  OA22X1 U5986 ( .IN1(n28631), .IN2(n268), .IN3(n28639), .IN4(n311), .Q(n6031)
         );
  OA221X1 U5987 ( .IN1(n28583), .IN2(n354), .IN3(n28591), .IN4(n397), .IN5(
        n6032), .Q(n6027) );
  OA22X1 U5988 ( .IN1(n28599), .IN2(n440), .IN3(n28607), .IN4(n483), .Q(n6032)
         );
  OA221X1 U5989 ( .IN1(n28551), .IN2(n526), .IN3(n28559), .IN4(n569), .IN5(
        n6033), .Q(n6026) );
  OA22X1 U5990 ( .IN1(n28567), .IN2(n612), .IN3(n28575), .IN4(n655), .Q(n6033)
         );
  NAND4X0 U5991 ( .IN1(n6034), .IN2(n6035), .IN3(n6036), .IN4(n6037), .QN(
        n6024) );
  OA221X1 U5992 ( .IN1(n28519), .IN2(n10), .IN3(n28527), .IN4(n53), .IN5(n6038), .Q(n6037) );
  OA22X1 U5993 ( .IN1(n28535), .IN2(n96), .IN3(n28543), .IN4(n139), .Q(n6038)
         );
  OA221X1 U5994 ( .IN1(n28487), .IN2(n182), .IN3(n28495), .IN4(n225), .IN5(
        n6039), .Q(n6036) );
  OA22X1 U5995 ( .IN1(n28503), .IN2(n268), .IN3(n28511), .IN4(n311), .Q(n6039)
         );
  OA221X1 U5996 ( .IN1(n28455), .IN2(n354), .IN3(n28463), .IN4(n397), .IN5(
        n6040), .Q(n6035) );
  OA22X1 U5997 ( .IN1(n28471), .IN2(n440), .IN3(n28479), .IN4(n483), .Q(n6040)
         );
  OA221X1 U5998 ( .IN1(n28423), .IN2(n526), .IN3(n28431), .IN4(n569), .IN5(
        n6041), .Q(n6034) );
  OA22X1 U5999 ( .IN1(n28439), .IN2(n612), .IN3(n28447), .IN4(n655), .Q(n6041)
         );
  NAND4X0 U6000 ( .IN1(n6042), .IN2(n6043), .IN3(n6044), .IN4(n6045), .QN(
        n6022) );
  OA221X1 U6001 ( .IN1(n28391), .IN2(n10), .IN3(n28399), .IN4(n53), .IN5(n6046), .Q(n6045) );
  OA22X1 U6002 ( .IN1(n28407), .IN2(n96), .IN3(n28415), .IN4(n139), .Q(n6046)
         );
  OA221X1 U6003 ( .IN1(n28359), .IN2(n182), .IN3(n28367), .IN4(n225), .IN5(
        n6047), .Q(n6044) );
  OA22X1 U6004 ( .IN1(n28375), .IN2(n268), .IN3(n28383), .IN4(n311), .Q(n6047)
         );
  OA221X1 U6005 ( .IN1(n28327), .IN2(n354), .IN3(n28335), .IN4(n397), .IN5(
        n6048), .Q(n6043) );
  OA22X1 U6006 ( .IN1(n28343), .IN2(n440), .IN3(n28351), .IN4(n483), .Q(n6048)
         );
  OA221X1 U6007 ( .IN1(n28295), .IN2(n526), .IN3(n28303), .IN4(n569), .IN5(
        n6049), .Q(n6042) );
  OA22X1 U6008 ( .IN1(n28311), .IN2(n612), .IN3(n28319), .IN4(n655), .Q(n6049)
         );
  NAND4X0 U6009 ( .IN1(n6050), .IN2(n6051), .IN3(n6052), .IN4(n6053), .QN(
        n6021) );
  OA221X1 U6010 ( .IN1(n28263), .IN2(n10), .IN3(n28271), .IN4(n53), .IN5(n6054), .Q(n6053) );
  OA22X1 U6011 ( .IN1(n28279), .IN2(n96), .IN3(n28287), .IN4(n139), .Q(n6054)
         );
  OA221X1 U6012 ( .IN1(n28231), .IN2(n182), .IN3(n28239), .IN4(n225), .IN5(
        n6055), .Q(n6052) );
  OA22X1 U6013 ( .IN1(n28247), .IN2(n268), .IN3(n28255), .IN4(n311), .Q(n6055)
         );
  OA221X1 U6014 ( .IN1(n28199), .IN2(n354), .IN3(n28207), .IN4(n397), .IN5(
        n6056), .Q(n6051) );
  OA22X1 U6015 ( .IN1(n28215), .IN2(n440), .IN3(n28223), .IN4(n483), .Q(n6056)
         );
  OA221X1 U6016 ( .IN1(n28167), .IN2(n526), .IN3(n28175), .IN4(n569), .IN5(
        n6057), .Q(n6050) );
  OA22X1 U6017 ( .IN1(n28183), .IN2(n612), .IN3(n28191), .IN4(n655), .Q(n6057)
         );
  AO221X1 U6018 ( .IN1(n2246), .IN2(n6058), .IN3(n2248), .IN4(n6059), .IN5(
        n6060), .Q(n6019) );
  AO22X1 U6019 ( .IN1(n2251), .IN2(n6061), .IN3(n2253), .IN4(n6062), .Q(n6060)
         );
  NAND4X0 U6020 ( .IN1(n6063), .IN2(n6064), .IN3(n6065), .IN4(n6066), .QN(
        n6062) );
  OA221X1 U6021 ( .IN1(n28135), .IN2(n9), .IN3(n28143), .IN4(n52), .IN5(n6067), 
        .Q(n6066) );
  OA22X1 U6022 ( .IN1(n28151), .IN2(n95), .IN3(n28159), .IN4(n138), .Q(n6067)
         );
  OA221X1 U6023 ( .IN1(n28103), .IN2(n181), .IN3(n28111), .IN4(n224), .IN5(
        n6068), .Q(n6065) );
  OA22X1 U6024 ( .IN1(n28119), .IN2(n267), .IN3(n28127), .IN4(n310), .Q(n6068)
         );
  OA221X1 U6025 ( .IN1(n28071), .IN2(n353), .IN3(n28079), .IN4(n396), .IN5(
        n6069), .Q(n6064) );
  OA22X1 U6026 ( .IN1(n28087), .IN2(n439), .IN3(n28095), .IN4(n482), .Q(n6069)
         );
  OA221X1 U6027 ( .IN1(n28039), .IN2(n525), .IN3(n28047), .IN4(n568), .IN5(
        n6070), .Q(n6063) );
  OA22X1 U6028 ( .IN1(n28055), .IN2(n611), .IN3(n28063), .IN4(n654), .Q(n6070)
         );
  NAND4X0 U6029 ( .IN1(n6071), .IN2(n6072), .IN3(n6073), .IN4(n6074), .QN(
        n6061) );
  OA221X1 U6030 ( .IN1(n28007), .IN2(n9), .IN3(n28015), .IN4(n52), .IN5(n6075), 
        .Q(n6074) );
  OA22X1 U6031 ( .IN1(n28023), .IN2(n95), .IN3(n28031), .IN4(n138), .Q(n6075)
         );
  OA221X1 U6032 ( .IN1(n27975), .IN2(n181), .IN3(n27983), .IN4(n224), .IN5(
        n6076), .Q(n6073) );
  OA22X1 U6033 ( .IN1(n27991), .IN2(n267), .IN3(n27999), .IN4(n310), .Q(n6076)
         );
  OA221X1 U6034 ( .IN1(n27943), .IN2(n353), .IN3(n27951), .IN4(n396), .IN5(
        n6077), .Q(n6072) );
  OA22X1 U6035 ( .IN1(n27959), .IN2(n439), .IN3(n27967), .IN4(n482), .Q(n6077)
         );
  OA221X1 U6036 ( .IN1(n27911), .IN2(n525), .IN3(n27919), .IN4(n568), .IN5(
        n6078), .Q(n6071) );
  OA22X1 U6037 ( .IN1(n27927), .IN2(n611), .IN3(n27935), .IN4(n654), .Q(n6078)
         );
  NAND4X0 U6038 ( .IN1(n6079), .IN2(n6080), .IN3(n6081), .IN4(n6082), .QN(
        n6059) );
  OA221X1 U6039 ( .IN1(n27879), .IN2(n9), .IN3(n27887), .IN4(n52), .IN5(n6083), 
        .Q(n6082) );
  OA22X1 U6040 ( .IN1(n27895), .IN2(n95), .IN3(n27903), .IN4(n138), .Q(n6083)
         );
  OA221X1 U6041 ( .IN1(n27847), .IN2(n181), .IN3(n27855), .IN4(n224), .IN5(
        n6084), .Q(n6081) );
  OA22X1 U6042 ( .IN1(n27863), .IN2(n267), .IN3(n27871), .IN4(n310), .Q(n6084)
         );
  OA221X1 U6043 ( .IN1(n27815), .IN2(n353), .IN3(n27823), .IN4(n396), .IN5(
        n6085), .Q(n6080) );
  OA22X1 U6044 ( .IN1(n27831), .IN2(n439), .IN3(n27839), .IN4(n482), .Q(n6085)
         );
  OA221X1 U6045 ( .IN1(n27783), .IN2(n525), .IN3(n27791), .IN4(n568), .IN5(
        n6086), .Q(n6079) );
  OA22X1 U6046 ( .IN1(n27799), .IN2(n611), .IN3(n27807), .IN4(n654), .Q(n6086)
         );
  NAND4X0 U6047 ( .IN1(n6087), .IN2(n6088), .IN3(n6089), .IN4(n6090), .QN(
        n6058) );
  OA221X1 U6048 ( .IN1(n27751), .IN2(n9), .IN3(n27759), .IN4(n52), .IN5(n6091), 
        .Q(n6090) );
  OA22X1 U6049 ( .IN1(n27767), .IN2(n95), .IN3(n27775), .IN4(n138), .Q(n6091)
         );
  OA221X1 U6050 ( .IN1(n27719), .IN2(n181), .IN3(n27727), .IN4(n224), .IN5(
        n6092), .Q(n6089) );
  OA22X1 U6051 ( .IN1(n27735), .IN2(n267), .IN3(n27743), .IN4(n310), .Q(n6092)
         );
  OA221X1 U6052 ( .IN1(n27687), .IN2(n353), .IN3(n27695), .IN4(n396), .IN5(
        n6093), .Q(n6088) );
  OA22X1 U6053 ( .IN1(n27703), .IN2(n439), .IN3(n27711), .IN4(n482), .Q(n6093)
         );
  OA221X1 U6054 ( .IN1(n27655), .IN2(n525), .IN3(n27663), .IN4(n568), .IN5(
        n6094), .Q(n6087) );
  OA22X1 U6055 ( .IN1(n27671), .IN2(n611), .IN3(n27679), .IN4(n654), .Q(n6094)
         );
  AO221X1 U6056 ( .IN1(n2287), .IN2(n6095), .IN3(n2289), .IN4(n6096), .IN5(
        n6097), .Q(n6018) );
  AO22X1 U6057 ( .IN1(n2292), .IN2(n6098), .IN3(n2294), .IN4(n6099), .Q(n6097)
         );
  NAND4X0 U6058 ( .IN1(n6100), .IN2(n6101), .IN3(n6102), .IN4(n6103), .QN(
        n6099) );
  OA221X1 U6059 ( .IN1(n29671), .IN2(n9), .IN3(n29679), .IN4(n52), .IN5(n6104), 
        .Q(n6103) );
  OA22X1 U6060 ( .IN1(n29687), .IN2(n95), .IN3(n29695), .IN4(n138), .Q(n6104)
         );
  OA221X1 U6061 ( .IN1(n29639), .IN2(n181), .IN3(n29647), .IN4(n224), .IN5(
        n6105), .Q(n6102) );
  OA22X1 U6062 ( .IN1(n29655), .IN2(n267), .IN3(n29663), .IN4(n310), .Q(n6105)
         );
  OA221X1 U6063 ( .IN1(n29607), .IN2(n353), .IN3(n29615), .IN4(n396), .IN5(
        n6106), .Q(n6101) );
  OA22X1 U6064 ( .IN1(n29623), .IN2(n439), .IN3(n29631), .IN4(n482), .Q(n6106)
         );
  OA221X1 U6065 ( .IN1(n29575), .IN2(n525), .IN3(n29583), .IN4(n568), .IN5(
        n6107), .Q(n6100) );
  OA22X1 U6066 ( .IN1(n29591), .IN2(n611), .IN3(n29599), .IN4(n654), .Q(n6107)
         );
  NAND4X0 U6067 ( .IN1(n6108), .IN2(n6109), .IN3(n6110), .IN4(n6111), .QN(
        n6098) );
  OA221X1 U6068 ( .IN1(n29543), .IN2(n9), .IN3(n29551), .IN4(n52), .IN5(n6112), 
        .Q(n6111) );
  OA22X1 U6069 ( .IN1(n29559), .IN2(n95), .IN3(n29567), .IN4(n138), .Q(n6112)
         );
  OA221X1 U6070 ( .IN1(n29511), .IN2(n181), .IN3(n29519), .IN4(n224), .IN5(
        n6113), .Q(n6110) );
  OA22X1 U6071 ( .IN1(n29527), .IN2(n267), .IN3(n29535), .IN4(n310), .Q(n6113)
         );
  OA221X1 U6072 ( .IN1(n29479), .IN2(n353), .IN3(n29487), .IN4(n396), .IN5(
        n6114), .Q(n6109) );
  OA22X1 U6073 ( .IN1(n29495), .IN2(n439), .IN3(n29503), .IN4(n482), .Q(n6114)
         );
  OA221X1 U6074 ( .IN1(n29447), .IN2(n525), .IN3(n29455), .IN4(n568), .IN5(
        n6115), .Q(n6108) );
  OA22X1 U6075 ( .IN1(n29463), .IN2(n611), .IN3(n29471), .IN4(n654), .Q(n6115)
         );
  NAND4X0 U6076 ( .IN1(n6116), .IN2(n6117), .IN3(n6118), .IN4(n6119), .QN(
        n6096) );
  OA221X1 U6077 ( .IN1(n29415), .IN2(n9), .IN3(n29423), .IN4(n52), .IN5(n6120), 
        .Q(n6119) );
  OA22X1 U6078 ( .IN1(n29431), .IN2(n95), .IN3(n29439), .IN4(n138), .Q(n6120)
         );
  OA221X1 U6079 ( .IN1(n29383), .IN2(n181), .IN3(n29391), .IN4(n224), .IN5(
        n6121), .Q(n6118) );
  OA22X1 U6080 ( .IN1(n29399), .IN2(n267), .IN3(n29407), .IN4(n310), .Q(n6121)
         );
  OA221X1 U6081 ( .IN1(n29351), .IN2(n353), .IN3(n29359), .IN4(n396), .IN5(
        n6122), .Q(n6117) );
  OA22X1 U6082 ( .IN1(n29367), .IN2(n439), .IN3(n29375), .IN4(n482), .Q(n6122)
         );
  OA221X1 U6083 ( .IN1(n29319), .IN2(n525), .IN3(n29327), .IN4(n568), .IN5(
        n6123), .Q(n6116) );
  OA22X1 U6084 ( .IN1(n29335), .IN2(n611), .IN3(n29343), .IN4(n654), .Q(n6123)
         );
  NAND4X0 U6085 ( .IN1(n6124), .IN2(n6125), .IN3(n6126), .IN4(n6127), .QN(
        n6095) );
  OA221X1 U6086 ( .IN1(n29287), .IN2(n9), .IN3(n29295), .IN4(n52), .IN5(n6128), 
        .Q(n6127) );
  OA22X1 U6087 ( .IN1(n29303), .IN2(n95), .IN3(n29311), .IN4(n138), .Q(n6128)
         );
  OA221X1 U6088 ( .IN1(n29255), .IN2(n181), .IN3(n29263), .IN4(n224), .IN5(
        n6129), .Q(n6126) );
  OA22X1 U6089 ( .IN1(n29271), .IN2(n267), .IN3(n29279), .IN4(n310), .Q(n6129)
         );
  OA221X1 U6090 ( .IN1(n29223), .IN2(n353), .IN3(n29231), .IN4(n396), .IN5(
        n6130), .Q(n6125) );
  OA22X1 U6091 ( .IN1(n29239), .IN2(n439), .IN3(n29247), .IN4(n482), .Q(n6130)
         );
  OA221X1 U6092 ( .IN1(n29191), .IN2(n525), .IN3(n29199), .IN4(n568), .IN5(
        n6131), .Q(n6124) );
  OA22X1 U6093 ( .IN1(n29207), .IN2(n611), .IN3(n29215), .IN4(n654), .Q(n6131)
         );
  AO221X1 U6094 ( .IN1(n2328), .IN2(n6132), .IN3(n2330), .IN4(n6133), .IN5(
        n6134), .Q(n6017) );
  AO22X1 U6095 ( .IN1(n2333), .IN2(n6135), .IN3(n2335), .IN4(n6136), .Q(n6134)
         );
  NAND4X0 U6096 ( .IN1(n6137), .IN2(n6138), .IN3(n6139), .IN4(n6140), .QN(
        n6136) );
  OA221X1 U6097 ( .IN1(n29159), .IN2(n9), .IN3(n29167), .IN4(n52), .IN5(n6141), 
        .Q(n6140) );
  OA22X1 U6098 ( .IN1(n29175), .IN2(n95), .IN3(n29183), .IN4(n138), .Q(n6141)
         );
  OA221X1 U6099 ( .IN1(n29127), .IN2(n181), .IN3(n29135), .IN4(n224), .IN5(
        n6142), .Q(n6139) );
  OA22X1 U6100 ( .IN1(n29143), .IN2(n267), .IN3(n29151), .IN4(n310), .Q(n6142)
         );
  OA221X1 U6101 ( .IN1(n29095), .IN2(n353), .IN3(n29103), .IN4(n396), .IN5(
        n6143), .Q(n6138) );
  OA22X1 U6102 ( .IN1(n29111), .IN2(n439), .IN3(n29119), .IN4(n482), .Q(n6143)
         );
  OA221X1 U6103 ( .IN1(n29063), .IN2(n525), .IN3(n29071), .IN4(n568), .IN5(
        n6144), .Q(n6137) );
  OA22X1 U6104 ( .IN1(n29079), .IN2(n611), .IN3(n29087), .IN4(n654), .Q(n6144)
         );
  NAND4X0 U6105 ( .IN1(n6145), .IN2(n6146), .IN3(n6147), .IN4(n6148), .QN(
        n6135) );
  OA221X1 U6106 ( .IN1(n29031), .IN2(n9), .IN3(n29039), .IN4(n52), .IN5(n6149), 
        .Q(n6148) );
  OA22X1 U6107 ( .IN1(n29047), .IN2(n95), .IN3(n29055), .IN4(n138), .Q(n6149)
         );
  OA221X1 U6108 ( .IN1(n28999), .IN2(n181), .IN3(n29007), .IN4(n224), .IN5(
        n6150), .Q(n6147) );
  OA22X1 U6109 ( .IN1(n29015), .IN2(n267), .IN3(n29023), .IN4(n310), .Q(n6150)
         );
  OA221X1 U6110 ( .IN1(n28967), .IN2(n353), .IN3(n28975), .IN4(n396), .IN5(
        n6151), .Q(n6146) );
  OA22X1 U6111 ( .IN1(n28983), .IN2(n439), .IN3(n28991), .IN4(n482), .Q(n6151)
         );
  OA221X1 U6112 ( .IN1(n28935), .IN2(n525), .IN3(n28943), .IN4(n568), .IN5(
        n6152), .Q(n6145) );
  OA22X1 U6113 ( .IN1(n28951), .IN2(n611), .IN3(n28959), .IN4(n654), .Q(n6152)
         );
  NAND4X0 U6114 ( .IN1(n6153), .IN2(n6154), .IN3(n6155), .IN4(n6156), .QN(
        n6133) );
  OA221X1 U6115 ( .IN1(n28903), .IN2(n9), .IN3(n28911), .IN4(n52), .IN5(n6157), 
        .Q(n6156) );
  OA22X1 U6116 ( .IN1(n28919), .IN2(n95), .IN3(n28927), .IN4(n138), .Q(n6157)
         );
  OA221X1 U6117 ( .IN1(n28871), .IN2(n181), .IN3(n28879), .IN4(n224), .IN5(
        n6158), .Q(n6155) );
  OA22X1 U6118 ( .IN1(n28887), .IN2(n267), .IN3(n28895), .IN4(n310), .Q(n6158)
         );
  OA221X1 U6119 ( .IN1(n28839), .IN2(n353), .IN3(n28847), .IN4(n396), .IN5(
        n6159), .Q(n6154) );
  OA22X1 U6120 ( .IN1(n28855), .IN2(n439), .IN3(n28863), .IN4(n482), .Q(n6159)
         );
  OA221X1 U6121 ( .IN1(n28807), .IN2(n525), .IN3(n28815), .IN4(n568), .IN5(
        n6160), .Q(n6153) );
  OA22X1 U6122 ( .IN1(n28823), .IN2(n611), .IN3(n28831), .IN4(n654), .Q(n6160)
         );
  NAND4X0 U6123 ( .IN1(n6161), .IN2(n6162), .IN3(n6163), .IN4(n6164), .QN(
        n6132) );
  OA221X1 U6124 ( .IN1(n28775), .IN2(n9), .IN3(n28783), .IN4(n52), .IN5(n6165), 
        .Q(n6164) );
  OA22X1 U6125 ( .IN1(n28791), .IN2(n95), .IN3(n28799), .IN4(n138), .Q(n6165)
         );
  OA221X1 U6126 ( .IN1(n28743), .IN2(n181), .IN3(n28751), .IN4(n224), .IN5(
        n6166), .Q(n6163) );
  OA22X1 U6127 ( .IN1(n28759), .IN2(n267), .IN3(n28767), .IN4(n310), .Q(n6166)
         );
  OA221X1 U6128 ( .IN1(n28711), .IN2(n353), .IN3(n28719), .IN4(n396), .IN5(
        n6167), .Q(n6162) );
  OA22X1 U6129 ( .IN1(n28727), .IN2(n439), .IN3(n28735), .IN4(n482), .Q(n6167)
         );
  OA221X1 U6130 ( .IN1(n28679), .IN2(n525), .IN3(n28687), .IN4(n568), .IN5(
        n6168), .Q(n6161) );
  OA22X1 U6131 ( .IN1(n28695), .IN2(n611), .IN3(n28703), .IN4(n654), .Q(n6168)
         );
  OR4X1 U6132 ( .IN1(n6169), .IN2(n6170), .IN3(n6171), .IN4(n6172), .Q(n2176)
         );
  AO221X1 U6133 ( .IN1(n2157), .IN2(n6173), .IN3(n2159), .IN4(n6174), .IN5(
        n6175), .Q(n6172) );
  AO22X1 U6134 ( .IN1(n2162), .IN2(n6176), .IN3(n2164), .IN4(n6177), .Q(n6175)
         );
  NAND4X0 U6135 ( .IN1(n6178), .IN2(n6179), .IN3(n6180), .IN4(n6181), .QN(
        n6177) );
  OA221X1 U6136 ( .IN1(n28646), .IN2(n8), .IN3(n28654), .IN4(n51), .IN5(n6182), 
        .Q(n6181) );
  OA22X1 U6137 ( .IN1(n28662), .IN2(n94), .IN3(n28670), .IN4(n137), .Q(n6182)
         );
  OA221X1 U6138 ( .IN1(n28614), .IN2(n180), .IN3(n28622), .IN4(n223), .IN5(
        n6183), .Q(n6180) );
  OA22X1 U6139 ( .IN1(n28630), .IN2(n266), .IN3(n28638), .IN4(n309), .Q(n6183)
         );
  OA221X1 U6140 ( .IN1(n28582), .IN2(n352), .IN3(n28590), .IN4(n395), .IN5(
        n6184), .Q(n6179) );
  OA22X1 U6141 ( .IN1(n28598), .IN2(n438), .IN3(n28606), .IN4(n481), .Q(n6184)
         );
  OA221X1 U6142 ( .IN1(n28550), .IN2(n524), .IN3(n28558), .IN4(n567), .IN5(
        n6185), .Q(n6178) );
  OA22X1 U6143 ( .IN1(n28566), .IN2(n610), .IN3(n28574), .IN4(n653), .Q(n6185)
         );
  NAND4X0 U6144 ( .IN1(n6186), .IN2(n6187), .IN3(n6188), .IN4(n6189), .QN(
        n6176) );
  OA221X1 U6145 ( .IN1(n28518), .IN2(n8), .IN3(n28526), .IN4(n51), .IN5(n6190), 
        .Q(n6189) );
  OA22X1 U6146 ( .IN1(n28534), .IN2(n94), .IN3(n28542), .IN4(n137), .Q(n6190)
         );
  OA221X1 U6147 ( .IN1(n28486), .IN2(n180), .IN3(n28494), .IN4(n223), .IN5(
        n6191), .Q(n6188) );
  OA22X1 U6148 ( .IN1(n28502), .IN2(n266), .IN3(n28510), .IN4(n309), .Q(n6191)
         );
  OA221X1 U6149 ( .IN1(n28454), .IN2(n352), .IN3(n28462), .IN4(n395), .IN5(
        n6192), .Q(n6187) );
  OA22X1 U6150 ( .IN1(n28470), .IN2(n438), .IN3(n28478), .IN4(n481), .Q(n6192)
         );
  OA221X1 U6151 ( .IN1(n28422), .IN2(n524), .IN3(n28430), .IN4(n567), .IN5(
        n6193), .Q(n6186) );
  OA22X1 U6152 ( .IN1(n28438), .IN2(n610), .IN3(n28446), .IN4(n653), .Q(n6193)
         );
  NAND4X0 U6153 ( .IN1(n6194), .IN2(n6195), .IN3(n6196), .IN4(n6197), .QN(
        n6174) );
  OA221X1 U6154 ( .IN1(n28390), .IN2(n8), .IN3(n28398), .IN4(n51), .IN5(n6198), 
        .Q(n6197) );
  OA22X1 U6155 ( .IN1(n28406), .IN2(n94), .IN3(n28414), .IN4(n137), .Q(n6198)
         );
  OA221X1 U6156 ( .IN1(n28358), .IN2(n180), .IN3(n28366), .IN4(n223), .IN5(
        n6199), .Q(n6196) );
  OA22X1 U6157 ( .IN1(n28374), .IN2(n266), .IN3(n28382), .IN4(n309), .Q(n6199)
         );
  OA221X1 U6158 ( .IN1(n28326), .IN2(n352), .IN3(n28334), .IN4(n395), .IN5(
        n6200), .Q(n6195) );
  OA22X1 U6159 ( .IN1(n28342), .IN2(n438), .IN3(n28350), .IN4(n481), .Q(n6200)
         );
  OA221X1 U6160 ( .IN1(n28294), .IN2(n524), .IN3(n28302), .IN4(n567), .IN5(
        n6201), .Q(n6194) );
  OA22X1 U6161 ( .IN1(n28310), .IN2(n610), .IN3(n28318), .IN4(n653), .Q(n6201)
         );
  NAND4X0 U6162 ( .IN1(n6202), .IN2(n6203), .IN3(n6204), .IN4(n6205), .QN(
        n6173) );
  OA221X1 U6163 ( .IN1(n28262), .IN2(n8), .IN3(n28270), .IN4(n51), .IN5(n6206), 
        .Q(n6205) );
  OA22X1 U6164 ( .IN1(n28278), .IN2(n94), .IN3(n28286), .IN4(n137), .Q(n6206)
         );
  OA221X1 U6165 ( .IN1(n28230), .IN2(n180), .IN3(n28238), .IN4(n223), .IN5(
        n6207), .Q(n6204) );
  OA22X1 U6166 ( .IN1(n28246), .IN2(n266), .IN3(n28254), .IN4(n309), .Q(n6207)
         );
  OA221X1 U6167 ( .IN1(n28198), .IN2(n352), .IN3(n28206), .IN4(n395), .IN5(
        n6208), .Q(n6203) );
  OA22X1 U6168 ( .IN1(n28214), .IN2(n438), .IN3(n28222), .IN4(n481), .Q(n6208)
         );
  OA221X1 U6169 ( .IN1(n28166), .IN2(n524), .IN3(n28174), .IN4(n567), .IN5(
        n6209), .Q(n6202) );
  OA22X1 U6170 ( .IN1(n28182), .IN2(n610), .IN3(n28190), .IN4(n653), .Q(n6209)
         );
  AO221X1 U6171 ( .IN1(n2246), .IN2(n6210), .IN3(n2248), .IN4(n6211), .IN5(
        n6212), .Q(n6171) );
  AO22X1 U6172 ( .IN1(n2251), .IN2(n6213), .IN3(n2253), .IN4(n6214), .Q(n6212)
         );
  NAND4X0 U6173 ( .IN1(n6215), .IN2(n6216), .IN3(n6217), .IN4(n6218), .QN(
        n6214) );
  OA221X1 U6174 ( .IN1(n28134), .IN2(n8), .IN3(n28142), .IN4(n51), .IN5(n6219), 
        .Q(n6218) );
  OA22X1 U6175 ( .IN1(n28150), .IN2(n94), .IN3(n28158), .IN4(n137), .Q(n6219)
         );
  OA221X1 U6176 ( .IN1(n28102), .IN2(n180), .IN3(n28110), .IN4(n223), .IN5(
        n6220), .Q(n6217) );
  OA22X1 U6177 ( .IN1(n28118), .IN2(n266), .IN3(n28126), .IN4(n309), .Q(n6220)
         );
  OA221X1 U6178 ( .IN1(n28070), .IN2(n352), .IN3(n28078), .IN4(n395), .IN5(
        n6221), .Q(n6216) );
  OA22X1 U6179 ( .IN1(n28086), .IN2(n438), .IN3(n28094), .IN4(n481), .Q(n6221)
         );
  OA221X1 U6180 ( .IN1(n28038), .IN2(n524), .IN3(n28046), .IN4(n567), .IN5(
        n6222), .Q(n6215) );
  OA22X1 U6181 ( .IN1(n28054), .IN2(n610), .IN3(n28062), .IN4(n653), .Q(n6222)
         );
  NAND4X0 U6182 ( .IN1(n6223), .IN2(n6224), .IN3(n6225), .IN4(n6226), .QN(
        n6213) );
  OA221X1 U6183 ( .IN1(n28006), .IN2(n8), .IN3(n28014), .IN4(n51), .IN5(n6227), 
        .Q(n6226) );
  OA22X1 U6184 ( .IN1(n28022), .IN2(n94), .IN3(n28030), .IN4(n137), .Q(n6227)
         );
  OA221X1 U6185 ( .IN1(n27974), .IN2(n180), .IN3(n27982), .IN4(n223), .IN5(
        n6228), .Q(n6225) );
  OA22X1 U6186 ( .IN1(n27990), .IN2(n266), .IN3(n27998), .IN4(n309), .Q(n6228)
         );
  OA221X1 U6187 ( .IN1(n27942), .IN2(n352), .IN3(n27950), .IN4(n395), .IN5(
        n6229), .Q(n6224) );
  OA22X1 U6188 ( .IN1(n27958), .IN2(n438), .IN3(n27966), .IN4(n481), .Q(n6229)
         );
  OA221X1 U6189 ( .IN1(n27910), .IN2(n524), .IN3(n27918), .IN4(n567), .IN5(
        n6230), .Q(n6223) );
  OA22X1 U6190 ( .IN1(n27926), .IN2(n610), .IN3(n27934), .IN4(n653), .Q(n6230)
         );
  NAND4X0 U6191 ( .IN1(n6231), .IN2(n6232), .IN3(n6233), .IN4(n6234), .QN(
        n6211) );
  OA221X1 U6192 ( .IN1(n27878), .IN2(n8), .IN3(n27886), .IN4(n51), .IN5(n6235), 
        .Q(n6234) );
  OA22X1 U6193 ( .IN1(n27894), .IN2(n94), .IN3(n27902), .IN4(n137), .Q(n6235)
         );
  OA221X1 U6194 ( .IN1(n27846), .IN2(n180), .IN3(n27854), .IN4(n223), .IN5(
        n6236), .Q(n6233) );
  OA22X1 U6195 ( .IN1(n27862), .IN2(n266), .IN3(n27870), .IN4(n309), .Q(n6236)
         );
  OA221X1 U6196 ( .IN1(n27814), .IN2(n352), .IN3(n27822), .IN4(n395), .IN5(
        n6237), .Q(n6232) );
  OA22X1 U6197 ( .IN1(n27830), .IN2(n438), .IN3(n27838), .IN4(n481), .Q(n6237)
         );
  OA221X1 U6198 ( .IN1(n27782), .IN2(n524), .IN3(n27790), .IN4(n567), .IN5(
        n6238), .Q(n6231) );
  OA22X1 U6199 ( .IN1(n27798), .IN2(n610), .IN3(n27806), .IN4(n653), .Q(n6238)
         );
  NAND4X0 U6200 ( .IN1(n6239), .IN2(n6240), .IN3(n6241), .IN4(n6242), .QN(
        n6210) );
  OA221X1 U6201 ( .IN1(n27750), .IN2(n8), .IN3(n27758), .IN4(n51), .IN5(n6243), 
        .Q(n6242) );
  OA22X1 U6202 ( .IN1(n27766), .IN2(n94), .IN3(n27774), .IN4(n137), .Q(n6243)
         );
  OA221X1 U6203 ( .IN1(n27718), .IN2(n180), .IN3(n27726), .IN4(n223), .IN5(
        n6244), .Q(n6241) );
  OA22X1 U6204 ( .IN1(n27734), .IN2(n266), .IN3(n27742), .IN4(n309), .Q(n6244)
         );
  OA221X1 U6205 ( .IN1(n27686), .IN2(n352), .IN3(n27694), .IN4(n395), .IN5(
        n6245), .Q(n6240) );
  OA22X1 U6206 ( .IN1(n27702), .IN2(n438), .IN3(n27710), .IN4(n481), .Q(n6245)
         );
  OA221X1 U6207 ( .IN1(n27654), .IN2(n524), .IN3(n27662), .IN4(n567), .IN5(
        n6246), .Q(n6239) );
  OA22X1 U6208 ( .IN1(n27670), .IN2(n610), .IN3(n27678), .IN4(n653), .Q(n6246)
         );
  AO221X1 U6209 ( .IN1(n2287), .IN2(n6247), .IN3(n2289), .IN4(n6248), .IN5(
        n6249), .Q(n6170) );
  AO22X1 U6210 ( .IN1(n2292), .IN2(n6250), .IN3(n2294), .IN4(n6251), .Q(n6249)
         );
  NAND4X0 U6211 ( .IN1(n6252), .IN2(n6253), .IN3(n6254), .IN4(n6255), .QN(
        n6251) );
  OA221X1 U6212 ( .IN1(n29670), .IN2(n8), .IN3(n29678), .IN4(n51), .IN5(n6256), 
        .Q(n6255) );
  OA22X1 U6213 ( .IN1(n29686), .IN2(n94), .IN3(n29694), .IN4(n137), .Q(n6256)
         );
  OA221X1 U6214 ( .IN1(n29638), .IN2(n180), .IN3(n29646), .IN4(n223), .IN5(
        n6257), .Q(n6254) );
  OA22X1 U6215 ( .IN1(n29654), .IN2(n266), .IN3(n29662), .IN4(n309), .Q(n6257)
         );
  OA221X1 U6216 ( .IN1(n29606), .IN2(n352), .IN3(n29614), .IN4(n395), .IN5(
        n6258), .Q(n6253) );
  OA22X1 U6217 ( .IN1(n29622), .IN2(n438), .IN3(n29630), .IN4(n481), .Q(n6258)
         );
  OA221X1 U6218 ( .IN1(n29574), .IN2(n524), .IN3(n29582), .IN4(n567), .IN5(
        n6259), .Q(n6252) );
  OA22X1 U6219 ( .IN1(n29590), .IN2(n610), .IN3(n29598), .IN4(n653), .Q(n6259)
         );
  NAND4X0 U6220 ( .IN1(n6260), .IN2(n6261), .IN3(n6262), .IN4(n6263), .QN(
        n6250) );
  OA221X1 U6221 ( .IN1(n29542), .IN2(n8), .IN3(n29550), .IN4(n51), .IN5(n6264), 
        .Q(n6263) );
  OA22X1 U6222 ( .IN1(n29558), .IN2(n94), .IN3(n29566), .IN4(n137), .Q(n6264)
         );
  OA221X1 U6223 ( .IN1(n29510), .IN2(n180), .IN3(n29518), .IN4(n223), .IN5(
        n6265), .Q(n6262) );
  OA22X1 U6224 ( .IN1(n29526), .IN2(n266), .IN3(n29534), .IN4(n309), .Q(n6265)
         );
  OA221X1 U6225 ( .IN1(n29478), .IN2(n352), .IN3(n29486), .IN4(n395), .IN5(
        n6266), .Q(n6261) );
  OA22X1 U6226 ( .IN1(n29494), .IN2(n438), .IN3(n29502), .IN4(n481), .Q(n6266)
         );
  OA221X1 U6227 ( .IN1(n29446), .IN2(n524), .IN3(n29454), .IN4(n567), .IN5(
        n6267), .Q(n6260) );
  OA22X1 U6228 ( .IN1(n29462), .IN2(n610), .IN3(n29470), .IN4(n653), .Q(n6267)
         );
  NAND4X0 U6229 ( .IN1(n6268), .IN2(n6269), .IN3(n6270), .IN4(n6271), .QN(
        n6248) );
  OA221X1 U6230 ( .IN1(n29414), .IN2(n8), .IN3(n29422), .IN4(n51), .IN5(n6272), 
        .Q(n6271) );
  OA22X1 U6231 ( .IN1(n29430), .IN2(n94), .IN3(n29438), .IN4(n137), .Q(n6272)
         );
  OA221X1 U6232 ( .IN1(n29382), .IN2(n180), .IN3(n29390), .IN4(n223), .IN5(
        n6273), .Q(n6270) );
  OA22X1 U6233 ( .IN1(n29398), .IN2(n266), .IN3(n29406), .IN4(n309), .Q(n6273)
         );
  OA221X1 U6234 ( .IN1(n29350), .IN2(n352), .IN3(n29358), .IN4(n395), .IN5(
        n6274), .Q(n6269) );
  OA22X1 U6235 ( .IN1(n29366), .IN2(n438), .IN3(n29374), .IN4(n481), .Q(n6274)
         );
  OA221X1 U6236 ( .IN1(n29318), .IN2(n524), .IN3(n29326), .IN4(n567), .IN5(
        n6275), .Q(n6268) );
  OA22X1 U6237 ( .IN1(n29334), .IN2(n610), .IN3(n29342), .IN4(n653), .Q(n6275)
         );
  NAND4X0 U6238 ( .IN1(n6276), .IN2(n6277), .IN3(n6278), .IN4(n6279), .QN(
        n6247) );
  OA221X1 U6239 ( .IN1(n29286), .IN2(n8), .IN3(n29294), .IN4(n51), .IN5(n6280), 
        .Q(n6279) );
  OA22X1 U6240 ( .IN1(n29302), .IN2(n94), .IN3(n29310), .IN4(n137), .Q(n6280)
         );
  OA221X1 U6241 ( .IN1(n29254), .IN2(n180), .IN3(n29262), .IN4(n223), .IN5(
        n6281), .Q(n6278) );
  OA22X1 U6242 ( .IN1(n29270), .IN2(n266), .IN3(n29278), .IN4(n309), .Q(n6281)
         );
  OA221X1 U6243 ( .IN1(n29222), .IN2(n352), .IN3(n29230), .IN4(n395), .IN5(
        n6282), .Q(n6277) );
  OA22X1 U6244 ( .IN1(n29238), .IN2(n438), .IN3(n29246), .IN4(n481), .Q(n6282)
         );
  OA221X1 U6245 ( .IN1(n29190), .IN2(n524), .IN3(n29198), .IN4(n567), .IN5(
        n6283), .Q(n6276) );
  OA22X1 U6246 ( .IN1(n29206), .IN2(n610), .IN3(n29214), .IN4(n653), .Q(n6283)
         );
  AO221X1 U6247 ( .IN1(n2328), .IN2(n6284), .IN3(n2330), .IN4(n6285), .IN5(
        n6286), .Q(n6169) );
  AO22X1 U6248 ( .IN1(n2333), .IN2(n6287), .IN3(n2335), .IN4(n6288), .Q(n6286)
         );
  NAND4X0 U6249 ( .IN1(n6289), .IN2(n6290), .IN3(n6291), .IN4(n6292), .QN(
        n6288) );
  OA221X1 U6250 ( .IN1(n29158), .IN2(n7), .IN3(n29166), .IN4(n50), .IN5(n6293), 
        .Q(n6292) );
  OA22X1 U6251 ( .IN1(n29174), .IN2(n93), .IN3(n29182), .IN4(n136), .Q(n6293)
         );
  OA221X1 U6252 ( .IN1(n29126), .IN2(n179), .IN3(n29134), .IN4(n222), .IN5(
        n6294), .Q(n6291) );
  OA22X1 U6253 ( .IN1(n29142), .IN2(n265), .IN3(n29150), .IN4(n308), .Q(n6294)
         );
  OA221X1 U6254 ( .IN1(n29094), .IN2(n351), .IN3(n29102), .IN4(n394), .IN5(
        n6295), .Q(n6290) );
  OA22X1 U6255 ( .IN1(n29110), .IN2(n437), .IN3(n29118), .IN4(n480), .Q(n6295)
         );
  OA221X1 U6256 ( .IN1(n29062), .IN2(n523), .IN3(n29070), .IN4(n566), .IN5(
        n6296), .Q(n6289) );
  OA22X1 U6257 ( .IN1(n29078), .IN2(n609), .IN3(n29086), .IN4(n652), .Q(n6296)
         );
  NAND4X0 U6258 ( .IN1(n6297), .IN2(n6298), .IN3(n6299), .IN4(n6300), .QN(
        n6287) );
  OA221X1 U6259 ( .IN1(n29030), .IN2(n7), .IN3(n29038), .IN4(n50), .IN5(n6301), 
        .Q(n6300) );
  OA22X1 U6260 ( .IN1(n29046), .IN2(n93), .IN3(n29054), .IN4(n136), .Q(n6301)
         );
  OA221X1 U6261 ( .IN1(n28998), .IN2(n179), .IN3(n29006), .IN4(n222), .IN5(
        n6302), .Q(n6299) );
  OA22X1 U6262 ( .IN1(n29014), .IN2(n265), .IN3(n29022), .IN4(n308), .Q(n6302)
         );
  OA221X1 U6263 ( .IN1(n28966), .IN2(n351), .IN3(n28974), .IN4(n394), .IN5(
        n6303), .Q(n6298) );
  OA22X1 U6264 ( .IN1(n28982), .IN2(n437), .IN3(n28990), .IN4(n480), .Q(n6303)
         );
  OA221X1 U6265 ( .IN1(n28934), .IN2(n523), .IN3(n28942), .IN4(n566), .IN5(
        n6304), .Q(n6297) );
  OA22X1 U6266 ( .IN1(n28950), .IN2(n609), .IN3(n28958), .IN4(n652), .Q(n6304)
         );
  NAND4X0 U6267 ( .IN1(n6305), .IN2(n6306), .IN3(n6307), .IN4(n6308), .QN(
        n6285) );
  OA221X1 U6268 ( .IN1(n28902), .IN2(n7), .IN3(n28910), .IN4(n50), .IN5(n6309), 
        .Q(n6308) );
  OA22X1 U6269 ( .IN1(n28918), .IN2(n93), .IN3(n28926), .IN4(n136), .Q(n6309)
         );
  OA221X1 U6270 ( .IN1(n28870), .IN2(n179), .IN3(n28878), .IN4(n222), .IN5(
        n6310), .Q(n6307) );
  OA22X1 U6271 ( .IN1(n28886), .IN2(n265), .IN3(n28894), .IN4(n308), .Q(n6310)
         );
  OA221X1 U6272 ( .IN1(n28838), .IN2(n351), .IN3(n28846), .IN4(n394), .IN5(
        n6311), .Q(n6306) );
  OA22X1 U6273 ( .IN1(n28854), .IN2(n437), .IN3(n28862), .IN4(n480), .Q(n6311)
         );
  OA221X1 U6274 ( .IN1(n28806), .IN2(n523), .IN3(n28814), .IN4(n566), .IN5(
        n6312), .Q(n6305) );
  OA22X1 U6275 ( .IN1(n28822), .IN2(n609), .IN3(n28830), .IN4(n652), .Q(n6312)
         );
  NAND4X0 U6276 ( .IN1(n6313), .IN2(n6314), .IN3(n6315), .IN4(n6316), .QN(
        n6284) );
  OA221X1 U6277 ( .IN1(n28774), .IN2(n7), .IN3(n28782), .IN4(n50), .IN5(n6317), 
        .Q(n6316) );
  OA22X1 U6278 ( .IN1(n28790), .IN2(n93), .IN3(n28798), .IN4(n136), .Q(n6317)
         );
  OA221X1 U6279 ( .IN1(n28742), .IN2(n179), .IN3(n28750), .IN4(n222), .IN5(
        n6318), .Q(n6315) );
  OA22X1 U6280 ( .IN1(n28758), .IN2(n265), .IN3(n28766), .IN4(n308), .Q(n6318)
         );
  OA221X1 U6281 ( .IN1(n28710), .IN2(n351), .IN3(n28718), .IN4(n394), .IN5(
        n6319), .Q(n6314) );
  OA22X1 U6282 ( .IN1(n28726), .IN2(n437), .IN3(n28734), .IN4(n480), .Q(n6319)
         );
  OA221X1 U6283 ( .IN1(n28678), .IN2(n523), .IN3(n28686), .IN4(n566), .IN5(
        n6320), .Q(n6313) );
  OA22X1 U6284 ( .IN1(n28694), .IN2(n609), .IN3(n28702), .IN4(n652), .Q(n6320)
         );
  OR4X1 U6285 ( .IN1(n6321), .IN2(n6322), .IN3(n6323), .IN4(n6324), .Q(n2175)
         );
  AO221X1 U6286 ( .IN1(n2157), .IN2(n6325), .IN3(n2159), .IN4(n6326), .IN5(
        n6327), .Q(n6324) );
  AO22X1 U6287 ( .IN1(n2162), .IN2(n6328), .IN3(n2164), .IN4(n6329), .Q(n6327)
         );
  NAND4X0 U6288 ( .IN1(n6330), .IN2(n6331), .IN3(n6332), .IN4(n6333), .QN(
        n6329) );
  OA221X1 U6289 ( .IN1(n28645), .IN2(n7), .IN3(n28653), .IN4(n50), .IN5(n6334), 
        .Q(n6333) );
  OA22X1 U6290 ( .IN1(n28661), .IN2(n93), .IN3(n28669), .IN4(n136), .Q(n6334)
         );
  OA221X1 U6291 ( .IN1(n28613), .IN2(n179), .IN3(n28621), .IN4(n222), .IN5(
        n6335), .Q(n6332) );
  OA22X1 U6292 ( .IN1(n28629), .IN2(n265), .IN3(n28637), .IN4(n308), .Q(n6335)
         );
  OA221X1 U6293 ( .IN1(n28581), .IN2(n351), .IN3(n28589), .IN4(n394), .IN5(
        n6336), .Q(n6331) );
  OA22X1 U6294 ( .IN1(n28597), .IN2(n437), .IN3(n28605), .IN4(n480), .Q(n6336)
         );
  OA221X1 U6295 ( .IN1(n28549), .IN2(n523), .IN3(n28557), .IN4(n566), .IN5(
        n6337), .Q(n6330) );
  OA22X1 U6296 ( .IN1(n28565), .IN2(n609), .IN3(n28573), .IN4(n652), .Q(n6337)
         );
  NAND4X0 U6297 ( .IN1(n6338), .IN2(n6339), .IN3(n6340), .IN4(n6341), .QN(
        n6328) );
  OA221X1 U6298 ( .IN1(n28517), .IN2(n7), .IN3(n28525), .IN4(n50), .IN5(n6342), 
        .Q(n6341) );
  OA22X1 U6299 ( .IN1(n28533), .IN2(n93), .IN3(n28541), .IN4(n136), .Q(n6342)
         );
  OA221X1 U6300 ( .IN1(n28485), .IN2(n179), .IN3(n28493), .IN4(n222), .IN5(
        n6343), .Q(n6340) );
  OA22X1 U6301 ( .IN1(n28501), .IN2(n265), .IN3(n28509), .IN4(n308), .Q(n6343)
         );
  OA221X1 U6302 ( .IN1(n28453), .IN2(n351), .IN3(n28461), .IN4(n394), .IN5(
        n6344), .Q(n6339) );
  OA22X1 U6303 ( .IN1(n28469), .IN2(n437), .IN3(n28477), .IN4(n480), .Q(n6344)
         );
  OA221X1 U6304 ( .IN1(n28421), .IN2(n523), .IN3(n28429), .IN4(n566), .IN5(
        n6345), .Q(n6338) );
  OA22X1 U6305 ( .IN1(n28437), .IN2(n609), .IN3(n28445), .IN4(n652), .Q(n6345)
         );
  NAND4X0 U6306 ( .IN1(n6346), .IN2(n6347), .IN3(n6348), .IN4(n6349), .QN(
        n6326) );
  OA221X1 U6307 ( .IN1(n28389), .IN2(n7), .IN3(n28397), .IN4(n50), .IN5(n6350), 
        .Q(n6349) );
  OA22X1 U6308 ( .IN1(n28405), .IN2(n93), .IN3(n28413), .IN4(n136), .Q(n6350)
         );
  OA221X1 U6309 ( .IN1(n28357), .IN2(n179), .IN3(n28365), .IN4(n222), .IN5(
        n6351), .Q(n6348) );
  OA22X1 U6310 ( .IN1(n28373), .IN2(n265), .IN3(n28381), .IN4(n308), .Q(n6351)
         );
  OA221X1 U6311 ( .IN1(n28325), .IN2(n351), .IN3(n28333), .IN4(n394), .IN5(
        n6352), .Q(n6347) );
  OA22X1 U6312 ( .IN1(n28341), .IN2(n437), .IN3(n28349), .IN4(n480), .Q(n6352)
         );
  OA221X1 U6313 ( .IN1(n28293), .IN2(n523), .IN3(n28301), .IN4(n566), .IN5(
        n6353), .Q(n6346) );
  OA22X1 U6314 ( .IN1(n28309), .IN2(n609), .IN3(n28317), .IN4(n652), .Q(n6353)
         );
  NAND4X0 U6315 ( .IN1(n6354), .IN2(n6355), .IN3(n6356), .IN4(n6357), .QN(
        n6325) );
  OA221X1 U6316 ( .IN1(n28261), .IN2(n7), .IN3(n28269), .IN4(n50), .IN5(n6358), 
        .Q(n6357) );
  OA22X1 U6317 ( .IN1(n28277), .IN2(n93), .IN3(n28285), .IN4(n136), .Q(n6358)
         );
  OA221X1 U6318 ( .IN1(n28229), .IN2(n179), .IN3(n28237), .IN4(n222), .IN5(
        n6359), .Q(n6356) );
  OA22X1 U6319 ( .IN1(n28245), .IN2(n265), .IN3(n28253), .IN4(n308), .Q(n6359)
         );
  OA221X1 U6320 ( .IN1(n28197), .IN2(n351), .IN3(n28205), .IN4(n394), .IN5(
        n6360), .Q(n6355) );
  OA22X1 U6321 ( .IN1(n28213), .IN2(n437), .IN3(n28221), .IN4(n480), .Q(n6360)
         );
  OA221X1 U6322 ( .IN1(n28165), .IN2(n523), .IN3(n28173), .IN4(n566), .IN5(
        n6361), .Q(n6354) );
  OA22X1 U6323 ( .IN1(n28181), .IN2(n609), .IN3(n28189), .IN4(n652), .Q(n6361)
         );
  AO221X1 U6324 ( .IN1(n2246), .IN2(n6362), .IN3(n2248), .IN4(n6363), .IN5(
        n6364), .Q(n6323) );
  AO22X1 U6325 ( .IN1(n2251), .IN2(n6365), .IN3(n2253), .IN4(n6366), .Q(n6364)
         );
  NAND4X0 U6326 ( .IN1(n6367), .IN2(n6368), .IN3(n6369), .IN4(n6370), .QN(
        n6366) );
  OA221X1 U6327 ( .IN1(n28133), .IN2(n7), .IN3(n28141), .IN4(n50), .IN5(n6371), 
        .Q(n6370) );
  OA22X1 U6328 ( .IN1(n28149), .IN2(n93), .IN3(n28157), .IN4(n136), .Q(n6371)
         );
  OA221X1 U6329 ( .IN1(n28101), .IN2(n179), .IN3(n28109), .IN4(n222), .IN5(
        n6372), .Q(n6369) );
  OA22X1 U6330 ( .IN1(n28117), .IN2(n265), .IN3(n28125), .IN4(n308), .Q(n6372)
         );
  OA221X1 U6331 ( .IN1(n28069), .IN2(n351), .IN3(n28077), .IN4(n394), .IN5(
        n6373), .Q(n6368) );
  OA22X1 U6332 ( .IN1(n28085), .IN2(n437), .IN3(n28093), .IN4(n480), .Q(n6373)
         );
  OA221X1 U6333 ( .IN1(n28037), .IN2(n523), .IN3(n28045), .IN4(n566), .IN5(
        n6374), .Q(n6367) );
  OA22X1 U6334 ( .IN1(n28053), .IN2(n609), .IN3(n28061), .IN4(n652), .Q(n6374)
         );
  NAND4X0 U6335 ( .IN1(n6375), .IN2(n6376), .IN3(n6377), .IN4(n6378), .QN(
        n6365) );
  OA221X1 U6336 ( .IN1(n28005), .IN2(n7), .IN3(n28013), .IN4(n50), .IN5(n6379), 
        .Q(n6378) );
  OA22X1 U6337 ( .IN1(n28021), .IN2(n93), .IN3(n28029), .IN4(n136), .Q(n6379)
         );
  OA221X1 U6338 ( .IN1(n27973), .IN2(n179), .IN3(n27981), .IN4(n222), .IN5(
        n6380), .Q(n6377) );
  OA22X1 U6339 ( .IN1(n27989), .IN2(n265), .IN3(n27997), .IN4(n308), .Q(n6380)
         );
  OA221X1 U6340 ( .IN1(n27941), .IN2(n351), .IN3(n27949), .IN4(n394), .IN5(
        n6381), .Q(n6376) );
  OA22X1 U6341 ( .IN1(n27957), .IN2(n437), .IN3(n27965), .IN4(n480), .Q(n6381)
         );
  OA221X1 U6342 ( .IN1(n27909), .IN2(n523), .IN3(n27917), .IN4(n566), .IN5(
        n6382), .Q(n6375) );
  OA22X1 U6343 ( .IN1(n27925), .IN2(n609), .IN3(n27933), .IN4(n652), .Q(n6382)
         );
  NAND4X0 U6344 ( .IN1(n6383), .IN2(n6384), .IN3(n6385), .IN4(n6386), .QN(
        n6363) );
  OA221X1 U6345 ( .IN1(n27877), .IN2(n7), .IN3(n27885), .IN4(n50), .IN5(n6387), 
        .Q(n6386) );
  OA22X1 U6346 ( .IN1(n27893), .IN2(n93), .IN3(n27901), .IN4(n136), .Q(n6387)
         );
  OA221X1 U6347 ( .IN1(n27845), .IN2(n179), .IN3(n27853), .IN4(n222), .IN5(
        n6388), .Q(n6385) );
  OA22X1 U6348 ( .IN1(n27861), .IN2(n265), .IN3(n27869), .IN4(n308), .Q(n6388)
         );
  OA221X1 U6349 ( .IN1(n27813), .IN2(n351), .IN3(n27821), .IN4(n394), .IN5(
        n6389), .Q(n6384) );
  OA22X1 U6350 ( .IN1(n27829), .IN2(n437), .IN3(n27837), .IN4(n480), .Q(n6389)
         );
  OA221X1 U6351 ( .IN1(n27781), .IN2(n523), .IN3(n27789), .IN4(n566), .IN5(
        n6390), .Q(n6383) );
  OA22X1 U6352 ( .IN1(n27797), .IN2(n609), .IN3(n27805), .IN4(n652), .Q(n6390)
         );
  NAND4X0 U6353 ( .IN1(n6391), .IN2(n6392), .IN3(n6393), .IN4(n6394), .QN(
        n6362) );
  OA221X1 U6354 ( .IN1(n27749), .IN2(n7), .IN3(n27757), .IN4(n50), .IN5(n6395), 
        .Q(n6394) );
  OA22X1 U6355 ( .IN1(n27765), .IN2(n93), .IN3(n27773), .IN4(n136), .Q(n6395)
         );
  OA221X1 U6356 ( .IN1(n27717), .IN2(n179), .IN3(n27725), .IN4(n222), .IN5(
        n6396), .Q(n6393) );
  OA22X1 U6357 ( .IN1(n27733), .IN2(n265), .IN3(n27741), .IN4(n308), .Q(n6396)
         );
  OA221X1 U6358 ( .IN1(n27685), .IN2(n351), .IN3(n27693), .IN4(n394), .IN5(
        n6397), .Q(n6392) );
  OA22X1 U6359 ( .IN1(n27701), .IN2(n437), .IN3(n27709), .IN4(n480), .Q(n6397)
         );
  OA221X1 U6360 ( .IN1(n27653), .IN2(n523), .IN3(n27661), .IN4(n566), .IN5(
        n6398), .Q(n6391) );
  OA22X1 U6361 ( .IN1(n27669), .IN2(n609), .IN3(n27677), .IN4(n652), .Q(n6398)
         );
  AO221X1 U6362 ( .IN1(n2287), .IN2(n6399), .IN3(n2289), .IN4(n6400), .IN5(
        n6401), .Q(n6322) );
  AO22X1 U6363 ( .IN1(n2292), .IN2(n6402), .IN3(n2294), .IN4(n6403), .Q(n6401)
         );
  NAND4X0 U6364 ( .IN1(n6404), .IN2(n6405), .IN3(n6406), .IN4(n6407), .QN(
        n6403) );
  OA221X1 U6365 ( .IN1(n29669), .IN2(n6), .IN3(n29677), .IN4(n49), .IN5(n6408), 
        .Q(n6407) );
  OA22X1 U6366 ( .IN1(n29685), .IN2(n92), .IN3(n29693), .IN4(n135), .Q(n6408)
         );
  OA221X1 U6367 ( .IN1(n29637), .IN2(n178), .IN3(n29645), .IN4(n221), .IN5(
        n6409), .Q(n6406) );
  OA22X1 U6368 ( .IN1(n29653), .IN2(n264), .IN3(n29661), .IN4(n307), .Q(n6409)
         );
  OA221X1 U6369 ( .IN1(n29605), .IN2(n350), .IN3(n29613), .IN4(n393), .IN5(
        n6410), .Q(n6405) );
  OA22X1 U6370 ( .IN1(n29621), .IN2(n436), .IN3(n29629), .IN4(n479), .Q(n6410)
         );
  OA221X1 U6371 ( .IN1(n29573), .IN2(n522), .IN3(n29581), .IN4(n565), .IN5(
        n6411), .Q(n6404) );
  OA22X1 U6372 ( .IN1(n29589), .IN2(n608), .IN3(n29597), .IN4(n651), .Q(n6411)
         );
  NAND4X0 U6373 ( .IN1(n6412), .IN2(n6413), .IN3(n6414), .IN4(n6415), .QN(
        n6402) );
  OA221X1 U6374 ( .IN1(n29541), .IN2(n6), .IN3(n29549), .IN4(n49), .IN5(n6416), 
        .Q(n6415) );
  OA22X1 U6375 ( .IN1(n29557), .IN2(n92), .IN3(n29565), .IN4(n135), .Q(n6416)
         );
  OA221X1 U6376 ( .IN1(n29509), .IN2(n178), .IN3(n29517), .IN4(n221), .IN5(
        n6417), .Q(n6414) );
  OA22X1 U6377 ( .IN1(n29525), .IN2(n264), .IN3(n29533), .IN4(n307), .Q(n6417)
         );
  OA221X1 U6378 ( .IN1(n29477), .IN2(n350), .IN3(n29485), .IN4(n393), .IN5(
        n6418), .Q(n6413) );
  OA22X1 U6379 ( .IN1(n29493), .IN2(n436), .IN3(n29501), .IN4(n479), .Q(n6418)
         );
  OA221X1 U6380 ( .IN1(n29445), .IN2(n522), .IN3(n29453), .IN4(n565), .IN5(
        n6419), .Q(n6412) );
  OA22X1 U6381 ( .IN1(n29461), .IN2(n608), .IN3(n29469), .IN4(n651), .Q(n6419)
         );
  NAND4X0 U6382 ( .IN1(n6420), .IN2(n6421), .IN3(n6422), .IN4(n6423), .QN(
        n6400) );
  OA221X1 U6383 ( .IN1(n29413), .IN2(n6), .IN3(n29421), .IN4(n49), .IN5(n6424), 
        .Q(n6423) );
  OA22X1 U6384 ( .IN1(n29429), .IN2(n92), .IN3(n29437), .IN4(n135), .Q(n6424)
         );
  OA221X1 U6385 ( .IN1(n29381), .IN2(n178), .IN3(n29389), .IN4(n221), .IN5(
        n6425), .Q(n6422) );
  OA22X1 U6386 ( .IN1(n29397), .IN2(n264), .IN3(n29405), .IN4(n307), .Q(n6425)
         );
  OA221X1 U6387 ( .IN1(n29349), .IN2(n350), .IN3(n29357), .IN4(n393), .IN5(
        n6426), .Q(n6421) );
  OA22X1 U6388 ( .IN1(n29365), .IN2(n436), .IN3(n29373), .IN4(n479), .Q(n6426)
         );
  OA221X1 U6389 ( .IN1(n29317), .IN2(n522), .IN3(n29325), .IN4(n565), .IN5(
        n6427), .Q(n6420) );
  OA22X1 U6390 ( .IN1(n29333), .IN2(n608), .IN3(n29341), .IN4(n651), .Q(n6427)
         );
  NAND4X0 U6391 ( .IN1(n6428), .IN2(n6429), .IN3(n6430), .IN4(n6431), .QN(
        n6399) );
  OA221X1 U6392 ( .IN1(n29285), .IN2(n6), .IN3(n29293), .IN4(n49), .IN5(n6432), 
        .Q(n6431) );
  OA22X1 U6393 ( .IN1(n29301), .IN2(n92), .IN3(n29309), .IN4(n135), .Q(n6432)
         );
  OA221X1 U6394 ( .IN1(n29253), .IN2(n178), .IN3(n29261), .IN4(n221), .IN5(
        n6433), .Q(n6430) );
  OA22X1 U6395 ( .IN1(n29269), .IN2(n264), .IN3(n29277), .IN4(n307), .Q(n6433)
         );
  OA221X1 U6396 ( .IN1(n29221), .IN2(n350), .IN3(n29229), .IN4(n393), .IN5(
        n6434), .Q(n6429) );
  OA22X1 U6397 ( .IN1(n29237), .IN2(n436), .IN3(n29245), .IN4(n479), .Q(n6434)
         );
  OA221X1 U6398 ( .IN1(n29189), .IN2(n522), .IN3(n29197), .IN4(n565), .IN5(
        n6435), .Q(n6428) );
  OA22X1 U6399 ( .IN1(n29205), .IN2(n608), .IN3(n29213), .IN4(n651), .Q(n6435)
         );
  AO221X1 U6400 ( .IN1(n2328), .IN2(n6436), .IN3(n2330), .IN4(n6437), .IN5(
        n6438), .Q(n6321) );
  AO22X1 U6401 ( .IN1(n2333), .IN2(n6439), .IN3(n2335), .IN4(n6440), .Q(n6438)
         );
  NAND4X0 U6402 ( .IN1(n6441), .IN2(n6442), .IN3(n6443), .IN4(n6444), .QN(
        n6440) );
  OA221X1 U6403 ( .IN1(n29157), .IN2(n6), .IN3(n29165), .IN4(n49), .IN5(n6445), 
        .Q(n6444) );
  OA22X1 U6404 ( .IN1(n29173), .IN2(n92), .IN3(n29181), .IN4(n135), .Q(n6445)
         );
  OA221X1 U6405 ( .IN1(n29125), .IN2(n178), .IN3(n29133), .IN4(n221), .IN5(
        n6446), .Q(n6443) );
  OA22X1 U6406 ( .IN1(n29141), .IN2(n264), .IN3(n29149), .IN4(n307), .Q(n6446)
         );
  OA221X1 U6407 ( .IN1(n29093), .IN2(n350), .IN3(n29101), .IN4(n393), .IN5(
        n6447), .Q(n6442) );
  OA22X1 U6408 ( .IN1(n29109), .IN2(n436), .IN3(n29117), .IN4(n479), .Q(n6447)
         );
  OA221X1 U6409 ( .IN1(n29061), .IN2(n522), .IN3(n29069), .IN4(n565), .IN5(
        n6448), .Q(n6441) );
  OA22X1 U6410 ( .IN1(n29077), .IN2(n608), .IN3(n29085), .IN4(n651), .Q(n6448)
         );
  NAND4X0 U6411 ( .IN1(n6449), .IN2(n6450), .IN3(n6451), .IN4(n6452), .QN(
        n6439) );
  OA221X1 U6412 ( .IN1(n29029), .IN2(n6), .IN3(n29037), .IN4(n49), .IN5(n6453), 
        .Q(n6452) );
  OA22X1 U6413 ( .IN1(n29045), .IN2(n92), .IN3(n29053), .IN4(n135), .Q(n6453)
         );
  OA221X1 U6414 ( .IN1(n28997), .IN2(n178), .IN3(n29005), .IN4(n221), .IN5(
        n6454), .Q(n6451) );
  OA22X1 U6415 ( .IN1(n29013), .IN2(n264), .IN3(n29021), .IN4(n307), .Q(n6454)
         );
  OA221X1 U6416 ( .IN1(n28965), .IN2(n350), .IN3(n28973), .IN4(n393), .IN5(
        n6455), .Q(n6450) );
  OA22X1 U6417 ( .IN1(n28981), .IN2(n436), .IN3(n28989), .IN4(n479), .Q(n6455)
         );
  OA221X1 U6418 ( .IN1(n28933), .IN2(n522), .IN3(n28941), .IN4(n565), .IN5(
        n6456), .Q(n6449) );
  OA22X1 U6419 ( .IN1(n28949), .IN2(n608), .IN3(n28957), .IN4(n651), .Q(n6456)
         );
  NAND4X0 U6420 ( .IN1(n6457), .IN2(n6458), .IN3(n6459), .IN4(n6460), .QN(
        n6437) );
  OA221X1 U6421 ( .IN1(n28901), .IN2(n6), .IN3(n28909), .IN4(n49), .IN5(n6461), 
        .Q(n6460) );
  OA22X1 U6422 ( .IN1(n28917), .IN2(n92), .IN3(n28925), .IN4(n135), .Q(n6461)
         );
  OA221X1 U6423 ( .IN1(n28869), .IN2(n178), .IN3(n28877), .IN4(n221), .IN5(
        n6462), .Q(n6459) );
  OA22X1 U6424 ( .IN1(n28885), .IN2(n264), .IN3(n28893), .IN4(n307), .Q(n6462)
         );
  OA221X1 U6425 ( .IN1(n28837), .IN2(n350), .IN3(n28845), .IN4(n393), .IN5(
        n6463), .Q(n6458) );
  OA22X1 U6426 ( .IN1(n28853), .IN2(n436), .IN3(n28861), .IN4(n479), .Q(n6463)
         );
  OA221X1 U6427 ( .IN1(n28805), .IN2(n522), .IN3(n28813), .IN4(n565), .IN5(
        n6464), .Q(n6457) );
  OA22X1 U6428 ( .IN1(n28821), .IN2(n608), .IN3(n28829), .IN4(n651), .Q(n6464)
         );
  NAND4X0 U6429 ( .IN1(n6465), .IN2(n6466), .IN3(n6467), .IN4(n6468), .QN(
        n6436) );
  OA221X1 U6430 ( .IN1(n28773), .IN2(n6), .IN3(n28781), .IN4(n49), .IN5(n6469), 
        .Q(n6468) );
  OA22X1 U6431 ( .IN1(n28789), .IN2(n92), .IN3(n28797), .IN4(n135), .Q(n6469)
         );
  OA221X1 U6432 ( .IN1(n28741), .IN2(n178), .IN3(n28749), .IN4(n221), .IN5(
        n6470), .Q(n6467) );
  OA22X1 U6433 ( .IN1(n28757), .IN2(n264), .IN3(n28765), .IN4(n307), .Q(n6470)
         );
  OA221X1 U6434 ( .IN1(n28709), .IN2(n350), .IN3(n28717), .IN4(n393), .IN5(
        n6471), .Q(n6466) );
  OA22X1 U6435 ( .IN1(n28725), .IN2(n436), .IN3(n28733), .IN4(n479), .Q(n6471)
         );
  OA221X1 U6436 ( .IN1(n28677), .IN2(n522), .IN3(n28685), .IN4(n565), .IN5(
        n6472), .Q(n6465) );
  OA22X1 U6437 ( .IN1(n28693), .IN2(n608), .IN3(n28701), .IN4(n651), .Q(n6472)
         );
  OR4X1 U6438 ( .IN1(n6473), .IN2(n6474), .IN3(n6475), .IN4(n6476), .Q(n2174)
         );
  AO221X1 U6439 ( .IN1(n2157), .IN2(n6477), .IN3(n2159), .IN4(n6478), .IN5(
        n6479), .Q(n6476) );
  AO22X1 U6440 ( .IN1(n2162), .IN2(n6480), .IN3(n2164), .IN4(n6481), .Q(n6479)
         );
  NAND4X0 U6441 ( .IN1(n6482), .IN2(n6483), .IN3(n6484), .IN4(n6485), .QN(
        n6481) );
  OA221X1 U6442 ( .IN1(n28644), .IN2(n6), .IN3(n28652), .IN4(n49), .IN5(n6486), 
        .Q(n6485) );
  OA22X1 U6443 ( .IN1(n28660), .IN2(n92), .IN3(n28668), .IN4(n135), .Q(n6486)
         );
  OA221X1 U6444 ( .IN1(n28612), .IN2(n178), .IN3(n28620), .IN4(n221), .IN5(
        n6487), .Q(n6484) );
  OA22X1 U6445 ( .IN1(n28628), .IN2(n264), .IN3(n28636), .IN4(n307), .Q(n6487)
         );
  OA221X1 U6446 ( .IN1(n28580), .IN2(n350), .IN3(n28588), .IN4(n393), .IN5(
        n6488), .Q(n6483) );
  OA22X1 U6447 ( .IN1(n28596), .IN2(n436), .IN3(n28604), .IN4(n479), .Q(n6488)
         );
  OA221X1 U6448 ( .IN1(n28548), .IN2(n522), .IN3(n28556), .IN4(n565), .IN5(
        n6489), .Q(n6482) );
  OA22X1 U6449 ( .IN1(n28564), .IN2(n608), .IN3(n28572), .IN4(n651), .Q(n6489)
         );
  NAND4X0 U6450 ( .IN1(n6490), .IN2(n6491), .IN3(n6492), .IN4(n6493), .QN(
        n6480) );
  OA221X1 U6451 ( .IN1(n28516), .IN2(n6), .IN3(n28524), .IN4(n49), .IN5(n6494), 
        .Q(n6493) );
  OA22X1 U6452 ( .IN1(n28532), .IN2(n92), .IN3(n28540), .IN4(n135), .Q(n6494)
         );
  OA221X1 U6453 ( .IN1(n28484), .IN2(n178), .IN3(n28492), .IN4(n221), .IN5(
        n6495), .Q(n6492) );
  OA22X1 U6454 ( .IN1(n28500), .IN2(n264), .IN3(n28508), .IN4(n307), .Q(n6495)
         );
  OA221X1 U6455 ( .IN1(n28452), .IN2(n350), .IN3(n28460), .IN4(n393), .IN5(
        n6496), .Q(n6491) );
  OA22X1 U6456 ( .IN1(n28468), .IN2(n436), .IN3(n28476), .IN4(n479), .Q(n6496)
         );
  OA221X1 U6457 ( .IN1(n28420), .IN2(n522), .IN3(n28428), .IN4(n565), .IN5(
        n6497), .Q(n6490) );
  OA22X1 U6458 ( .IN1(n28436), .IN2(n608), .IN3(n28444), .IN4(n651), .Q(n6497)
         );
  NAND4X0 U6459 ( .IN1(n6498), .IN2(n6499), .IN3(n6500), .IN4(n6501), .QN(
        n6478) );
  OA221X1 U6460 ( .IN1(n28388), .IN2(n6), .IN3(n28396), .IN4(n49), .IN5(n6502), 
        .Q(n6501) );
  OA22X1 U6461 ( .IN1(n28404), .IN2(n92), .IN3(n28412), .IN4(n135), .Q(n6502)
         );
  OA221X1 U6462 ( .IN1(n28356), .IN2(n178), .IN3(n28364), .IN4(n221), .IN5(
        n6503), .Q(n6500) );
  OA22X1 U6463 ( .IN1(n28372), .IN2(n264), .IN3(n28380), .IN4(n307), .Q(n6503)
         );
  OA221X1 U6464 ( .IN1(n28324), .IN2(n350), .IN3(n28332), .IN4(n393), .IN5(
        n6504), .Q(n6499) );
  OA22X1 U6465 ( .IN1(n28340), .IN2(n436), .IN3(n28348), .IN4(n479), .Q(n6504)
         );
  OA221X1 U6466 ( .IN1(n28292), .IN2(n522), .IN3(n28300), .IN4(n565), .IN5(
        n6505), .Q(n6498) );
  OA22X1 U6467 ( .IN1(n28308), .IN2(n608), .IN3(n28316), .IN4(n651), .Q(n6505)
         );
  NAND4X0 U6468 ( .IN1(n6506), .IN2(n6507), .IN3(n6508), .IN4(n6509), .QN(
        n6477) );
  OA221X1 U6469 ( .IN1(n28260), .IN2(n6), .IN3(n28268), .IN4(n49), .IN5(n6510), 
        .Q(n6509) );
  OA22X1 U6470 ( .IN1(n28276), .IN2(n92), .IN3(n28284), .IN4(n135), .Q(n6510)
         );
  OA221X1 U6471 ( .IN1(n28228), .IN2(n178), .IN3(n28236), .IN4(n221), .IN5(
        n6511), .Q(n6508) );
  OA22X1 U6472 ( .IN1(n28244), .IN2(n264), .IN3(n28252), .IN4(n307), .Q(n6511)
         );
  OA221X1 U6473 ( .IN1(n28196), .IN2(n350), .IN3(n28204), .IN4(n393), .IN5(
        n6512), .Q(n6507) );
  OA22X1 U6474 ( .IN1(n28212), .IN2(n436), .IN3(n28220), .IN4(n479), .Q(n6512)
         );
  OA221X1 U6475 ( .IN1(n28164), .IN2(n522), .IN3(n28172), .IN4(n565), .IN5(
        n6513), .Q(n6506) );
  OA22X1 U6476 ( .IN1(n28180), .IN2(n608), .IN3(n28188), .IN4(n651), .Q(n6513)
         );
  AO221X1 U6477 ( .IN1(n2246), .IN2(n6514), .IN3(n2248), .IN4(n6515), .IN5(
        n6516), .Q(n6475) );
  AO22X1 U6478 ( .IN1(n2251), .IN2(n6517), .IN3(n2253), .IN4(n6518), .Q(n6516)
         );
  NAND4X0 U6479 ( .IN1(n6519), .IN2(n6520), .IN3(n6521), .IN4(n6522), .QN(
        n6518) );
  OA221X1 U6480 ( .IN1(n28132), .IN2(n5), .IN3(n28140), .IN4(n48), .IN5(n6523), 
        .Q(n6522) );
  OA22X1 U6481 ( .IN1(n28148), .IN2(n91), .IN3(n28156), .IN4(n134), .Q(n6523)
         );
  OA221X1 U6482 ( .IN1(n28100), .IN2(n177), .IN3(n28108), .IN4(n220), .IN5(
        n6524), .Q(n6521) );
  OA22X1 U6483 ( .IN1(n28116), .IN2(n263), .IN3(n28124), .IN4(n306), .Q(n6524)
         );
  OA221X1 U6484 ( .IN1(n28068), .IN2(n349), .IN3(n28076), .IN4(n392), .IN5(
        n6525), .Q(n6520) );
  OA22X1 U6485 ( .IN1(n28084), .IN2(n435), .IN3(n28092), .IN4(n478), .Q(n6525)
         );
  OA221X1 U6486 ( .IN1(n28036), .IN2(n521), .IN3(n28044), .IN4(n564), .IN5(
        n6526), .Q(n6519) );
  OA22X1 U6487 ( .IN1(n28052), .IN2(n607), .IN3(n28060), .IN4(n650), .Q(n6526)
         );
  NAND4X0 U6488 ( .IN1(n6527), .IN2(n6528), .IN3(n6529), .IN4(n6530), .QN(
        n6517) );
  OA221X1 U6489 ( .IN1(n28004), .IN2(n5), .IN3(n28012), .IN4(n48), .IN5(n6531), 
        .Q(n6530) );
  OA22X1 U6490 ( .IN1(n28020), .IN2(n91), .IN3(n28028), .IN4(n134), .Q(n6531)
         );
  OA221X1 U6491 ( .IN1(n27972), .IN2(n177), .IN3(n27980), .IN4(n220), .IN5(
        n6532), .Q(n6529) );
  OA22X1 U6492 ( .IN1(n27988), .IN2(n263), .IN3(n27996), .IN4(n306), .Q(n6532)
         );
  OA221X1 U6493 ( .IN1(n27940), .IN2(n349), .IN3(n27948), .IN4(n392), .IN5(
        n6533), .Q(n6528) );
  OA22X1 U6494 ( .IN1(n27956), .IN2(n435), .IN3(n27964), .IN4(n478), .Q(n6533)
         );
  OA221X1 U6495 ( .IN1(n27908), .IN2(n521), .IN3(n27916), .IN4(n564), .IN5(
        n6534), .Q(n6527) );
  OA22X1 U6496 ( .IN1(n27924), .IN2(n607), .IN3(n27932), .IN4(n650), .Q(n6534)
         );
  NAND4X0 U6497 ( .IN1(n6535), .IN2(n6536), .IN3(n6537), .IN4(n6538), .QN(
        n6515) );
  OA221X1 U6498 ( .IN1(n27876), .IN2(n5), .IN3(n27884), .IN4(n48), .IN5(n6539), 
        .Q(n6538) );
  OA22X1 U6499 ( .IN1(n27892), .IN2(n91), .IN3(n27900), .IN4(n134), .Q(n6539)
         );
  OA221X1 U6500 ( .IN1(n27844), .IN2(n177), .IN3(n27852), .IN4(n220), .IN5(
        n6540), .Q(n6537) );
  OA22X1 U6501 ( .IN1(n27860), .IN2(n263), .IN3(n27868), .IN4(n306), .Q(n6540)
         );
  OA221X1 U6502 ( .IN1(n27812), .IN2(n349), .IN3(n27820), .IN4(n392), .IN5(
        n6541), .Q(n6536) );
  OA22X1 U6503 ( .IN1(n27828), .IN2(n435), .IN3(n27836), .IN4(n478), .Q(n6541)
         );
  OA221X1 U6504 ( .IN1(n27780), .IN2(n521), .IN3(n27788), .IN4(n564), .IN5(
        n6542), .Q(n6535) );
  OA22X1 U6505 ( .IN1(n27796), .IN2(n607), .IN3(n27804), .IN4(n650), .Q(n6542)
         );
  NAND4X0 U6506 ( .IN1(n6543), .IN2(n6544), .IN3(n6545), .IN4(n6546), .QN(
        n6514) );
  OA221X1 U6507 ( .IN1(n27748), .IN2(n5), .IN3(n27756), .IN4(n48), .IN5(n6547), 
        .Q(n6546) );
  OA22X1 U6508 ( .IN1(n27764), .IN2(n91), .IN3(n27772), .IN4(n134), .Q(n6547)
         );
  OA221X1 U6509 ( .IN1(n27716), .IN2(n177), .IN3(n27724), .IN4(n220), .IN5(
        n6548), .Q(n6545) );
  OA22X1 U6510 ( .IN1(n27732), .IN2(n263), .IN3(n27740), .IN4(n306), .Q(n6548)
         );
  OA221X1 U6511 ( .IN1(n27684), .IN2(n349), .IN3(n27692), .IN4(n392), .IN5(
        n6549), .Q(n6544) );
  OA22X1 U6512 ( .IN1(n27700), .IN2(n435), .IN3(n27708), .IN4(n478), .Q(n6549)
         );
  OA221X1 U6513 ( .IN1(n27652), .IN2(n521), .IN3(n27660), .IN4(n564), .IN5(
        n6550), .Q(n6543) );
  OA22X1 U6514 ( .IN1(n27668), .IN2(n607), .IN3(n27676), .IN4(n650), .Q(n6550)
         );
  AO221X1 U6515 ( .IN1(n2287), .IN2(n6551), .IN3(n2289), .IN4(n6552), .IN5(
        n6553), .Q(n6474) );
  AO22X1 U6516 ( .IN1(n2292), .IN2(n6554), .IN3(n2294), .IN4(n6555), .Q(n6553)
         );
  NAND4X0 U6517 ( .IN1(n6556), .IN2(n6557), .IN3(n6558), .IN4(n6559), .QN(
        n6555) );
  OA221X1 U6518 ( .IN1(n29668), .IN2(n5), .IN3(n29676), .IN4(n48), .IN5(n6560), 
        .Q(n6559) );
  OA22X1 U6519 ( .IN1(n29684), .IN2(n91), .IN3(n29692), .IN4(n134), .Q(n6560)
         );
  OA221X1 U6520 ( .IN1(n29636), .IN2(n177), .IN3(n29644), .IN4(n220), .IN5(
        n6561), .Q(n6558) );
  OA22X1 U6521 ( .IN1(n29652), .IN2(n263), .IN3(n29660), .IN4(n306), .Q(n6561)
         );
  OA221X1 U6522 ( .IN1(n29604), .IN2(n349), .IN3(n29612), .IN4(n392), .IN5(
        n6562), .Q(n6557) );
  OA22X1 U6523 ( .IN1(n29620), .IN2(n435), .IN3(n29628), .IN4(n478), .Q(n6562)
         );
  OA221X1 U6524 ( .IN1(n29572), .IN2(n521), .IN3(n29580), .IN4(n564), .IN5(
        n6563), .Q(n6556) );
  OA22X1 U6525 ( .IN1(n29588), .IN2(n607), .IN3(n29596), .IN4(n650), .Q(n6563)
         );
  NAND4X0 U6526 ( .IN1(n6564), .IN2(n6565), .IN3(n6566), .IN4(n6567), .QN(
        n6554) );
  OA221X1 U6527 ( .IN1(n29540), .IN2(n5), .IN3(n29548), .IN4(n48), .IN5(n6568), 
        .Q(n6567) );
  OA22X1 U6528 ( .IN1(n29556), .IN2(n91), .IN3(n29564), .IN4(n134), .Q(n6568)
         );
  OA221X1 U6529 ( .IN1(n29508), .IN2(n177), .IN3(n29516), .IN4(n220), .IN5(
        n6569), .Q(n6566) );
  OA22X1 U6530 ( .IN1(n29524), .IN2(n263), .IN3(n29532), .IN4(n306), .Q(n6569)
         );
  OA221X1 U6531 ( .IN1(n29476), .IN2(n349), .IN3(n29484), .IN4(n392), .IN5(
        n6570), .Q(n6565) );
  OA22X1 U6532 ( .IN1(n29492), .IN2(n435), .IN3(n29500), .IN4(n478), .Q(n6570)
         );
  OA221X1 U6533 ( .IN1(n29444), .IN2(n521), .IN3(n29452), .IN4(n564), .IN5(
        n6571), .Q(n6564) );
  OA22X1 U6534 ( .IN1(n29460), .IN2(n607), .IN3(n29468), .IN4(n650), .Q(n6571)
         );
  NAND4X0 U6535 ( .IN1(n6572), .IN2(n6573), .IN3(n6574), .IN4(n6575), .QN(
        n6552) );
  OA221X1 U6536 ( .IN1(n29412), .IN2(n5), .IN3(n29420), .IN4(n48), .IN5(n6576), 
        .Q(n6575) );
  OA22X1 U6537 ( .IN1(n29428), .IN2(n91), .IN3(n29436), .IN4(n134), .Q(n6576)
         );
  OA221X1 U6538 ( .IN1(n29380), .IN2(n177), .IN3(n29388), .IN4(n220), .IN5(
        n6577), .Q(n6574) );
  OA22X1 U6539 ( .IN1(n29396), .IN2(n263), .IN3(n29404), .IN4(n306), .Q(n6577)
         );
  OA221X1 U6540 ( .IN1(n29348), .IN2(n349), .IN3(n29356), .IN4(n392), .IN5(
        n6578), .Q(n6573) );
  OA22X1 U6541 ( .IN1(n29364), .IN2(n435), .IN3(n29372), .IN4(n478), .Q(n6578)
         );
  OA221X1 U6542 ( .IN1(n29316), .IN2(n521), .IN3(n29324), .IN4(n564), .IN5(
        n6579), .Q(n6572) );
  OA22X1 U6543 ( .IN1(n29332), .IN2(n607), .IN3(n29340), .IN4(n650), .Q(n6579)
         );
  NAND4X0 U6544 ( .IN1(n6580), .IN2(n6581), .IN3(n6582), .IN4(n6583), .QN(
        n6551) );
  OA221X1 U6545 ( .IN1(n29284), .IN2(n5), .IN3(n29292), .IN4(n48), .IN5(n6584), 
        .Q(n6583) );
  OA22X1 U6546 ( .IN1(n29300), .IN2(n91), .IN3(n29308), .IN4(n134), .Q(n6584)
         );
  OA221X1 U6547 ( .IN1(n29252), .IN2(n177), .IN3(n29260), .IN4(n220), .IN5(
        n6585), .Q(n6582) );
  OA22X1 U6548 ( .IN1(n29268), .IN2(n263), .IN3(n29276), .IN4(n306), .Q(n6585)
         );
  OA221X1 U6549 ( .IN1(n29220), .IN2(n349), .IN3(n29228), .IN4(n392), .IN5(
        n6586), .Q(n6581) );
  OA22X1 U6550 ( .IN1(n29236), .IN2(n435), .IN3(n29244), .IN4(n478), .Q(n6586)
         );
  OA221X1 U6551 ( .IN1(n29188), .IN2(n521), .IN3(n29196), .IN4(n564), .IN5(
        n6587), .Q(n6580) );
  OA22X1 U6552 ( .IN1(n29204), .IN2(n607), .IN3(n29212), .IN4(n650), .Q(n6587)
         );
  AO221X1 U6553 ( .IN1(n2328), .IN2(n6588), .IN3(n2330), .IN4(n6589), .IN5(
        n6590), .Q(n6473) );
  AO22X1 U6554 ( .IN1(n2333), .IN2(n6591), .IN3(n2335), .IN4(n6592), .Q(n6590)
         );
  NAND4X0 U6555 ( .IN1(n6593), .IN2(n6594), .IN3(n6595), .IN4(n6596), .QN(
        n6592) );
  OA221X1 U6556 ( .IN1(n29156), .IN2(n5), .IN3(n29164), .IN4(n48), .IN5(n6597), 
        .Q(n6596) );
  OA22X1 U6557 ( .IN1(n29172), .IN2(n91), .IN3(n29180), .IN4(n134), .Q(n6597)
         );
  OA221X1 U6558 ( .IN1(n29124), .IN2(n177), .IN3(n29132), .IN4(n220), .IN5(
        n6598), .Q(n6595) );
  OA22X1 U6559 ( .IN1(n29140), .IN2(n263), .IN3(n29148), .IN4(n306), .Q(n6598)
         );
  OA221X1 U6560 ( .IN1(n29092), .IN2(n349), .IN3(n29100), .IN4(n392), .IN5(
        n6599), .Q(n6594) );
  OA22X1 U6561 ( .IN1(n29108), .IN2(n435), .IN3(n29116), .IN4(n478), .Q(n6599)
         );
  OA221X1 U6562 ( .IN1(n29060), .IN2(n521), .IN3(n29068), .IN4(n564), .IN5(
        n6600), .Q(n6593) );
  OA22X1 U6563 ( .IN1(n29076), .IN2(n607), .IN3(n29084), .IN4(n650), .Q(n6600)
         );
  NAND4X0 U6564 ( .IN1(n6601), .IN2(n6602), .IN3(n6603), .IN4(n6604), .QN(
        n6591) );
  OA221X1 U6565 ( .IN1(n29028), .IN2(n5), .IN3(n29036), .IN4(n48), .IN5(n6605), 
        .Q(n6604) );
  OA22X1 U6566 ( .IN1(n29044), .IN2(n91), .IN3(n29052), .IN4(n134), .Q(n6605)
         );
  OA221X1 U6567 ( .IN1(n28996), .IN2(n177), .IN3(n29004), .IN4(n220), .IN5(
        n6606), .Q(n6603) );
  OA22X1 U6568 ( .IN1(n29012), .IN2(n263), .IN3(n29020), .IN4(n306), .Q(n6606)
         );
  OA221X1 U6569 ( .IN1(n28964), .IN2(n349), .IN3(n28972), .IN4(n392), .IN5(
        n6607), .Q(n6602) );
  OA22X1 U6570 ( .IN1(n28980), .IN2(n435), .IN3(n28988), .IN4(n478), .Q(n6607)
         );
  OA221X1 U6571 ( .IN1(n28932), .IN2(n521), .IN3(n28940), .IN4(n564), .IN5(
        n6608), .Q(n6601) );
  OA22X1 U6572 ( .IN1(n28948), .IN2(n607), .IN3(n28956), .IN4(n650), .Q(n6608)
         );
  NAND4X0 U6573 ( .IN1(n6609), .IN2(n6610), .IN3(n6611), .IN4(n6612), .QN(
        n6589) );
  OA221X1 U6574 ( .IN1(n28900), .IN2(n5), .IN3(n28908), .IN4(n48), .IN5(n6613), 
        .Q(n6612) );
  OA22X1 U6575 ( .IN1(n28916), .IN2(n91), .IN3(n28924), .IN4(n134), .Q(n6613)
         );
  OA221X1 U6576 ( .IN1(n28868), .IN2(n177), .IN3(n28876), .IN4(n220), .IN5(
        n6614), .Q(n6611) );
  OA22X1 U6577 ( .IN1(n28884), .IN2(n263), .IN3(n28892), .IN4(n306), .Q(n6614)
         );
  OA221X1 U6578 ( .IN1(n28836), .IN2(n349), .IN3(n28844), .IN4(n392), .IN5(
        n6615), .Q(n6610) );
  OA22X1 U6579 ( .IN1(n28852), .IN2(n435), .IN3(n28860), .IN4(n478), .Q(n6615)
         );
  OA221X1 U6580 ( .IN1(n28804), .IN2(n521), .IN3(n28812), .IN4(n564), .IN5(
        n6616), .Q(n6609) );
  OA22X1 U6581 ( .IN1(n28820), .IN2(n607), .IN3(n28828), .IN4(n650), .Q(n6616)
         );
  NAND4X0 U6582 ( .IN1(n6617), .IN2(n6618), .IN3(n6619), .IN4(n6620), .QN(
        n6588) );
  OA221X1 U6583 ( .IN1(n28772), .IN2(n5), .IN3(n28780), .IN4(n48), .IN5(n6621), 
        .Q(n6620) );
  OA22X1 U6584 ( .IN1(n28788), .IN2(n91), .IN3(n28796), .IN4(n134), .Q(n6621)
         );
  OA221X1 U6585 ( .IN1(n28740), .IN2(n177), .IN3(n28748), .IN4(n220), .IN5(
        n6622), .Q(n6619) );
  OA22X1 U6586 ( .IN1(n28756), .IN2(n263), .IN3(n28764), .IN4(n306), .Q(n6622)
         );
  OA221X1 U6587 ( .IN1(n28708), .IN2(n349), .IN3(n28716), .IN4(n392), .IN5(
        n6623), .Q(n6618) );
  OA22X1 U6588 ( .IN1(n28724), .IN2(n435), .IN3(n28732), .IN4(n478), .Q(n6623)
         );
  OA221X1 U6589 ( .IN1(n28676), .IN2(n521), .IN3(n28684), .IN4(n564), .IN5(
        n6624), .Q(n6617) );
  OA22X1 U6590 ( .IN1(n28692), .IN2(n607), .IN3(n28700), .IN4(n650), .Q(n6624)
         );
  OR4X1 U6591 ( .IN1(n6625), .IN2(n6626), .IN3(n6627), .IN4(n6628), .Q(n2173)
         );
  AO221X1 U6592 ( .IN1(n2157), .IN2(n6629), .IN3(n2159), .IN4(n6630), .IN5(
        n6631), .Q(n6628) );
  AO22X1 U6593 ( .IN1(n2162), .IN2(n6632), .IN3(n2164), .IN4(n6633), .Q(n6631)
         );
  NAND4X0 U6594 ( .IN1(n6634), .IN2(n6635), .IN3(n6636), .IN4(n6637), .QN(
        n6633) );
  OA221X1 U6595 ( .IN1(n28643), .IN2(n4), .IN3(n28651), .IN4(n47), .IN5(n6638), 
        .Q(n6637) );
  OA22X1 U6596 ( .IN1(n28659), .IN2(n90), .IN3(n28667), .IN4(n133), .Q(n6638)
         );
  OA221X1 U6597 ( .IN1(n28611), .IN2(n176), .IN3(n28619), .IN4(n219), .IN5(
        n6639), .Q(n6636) );
  OA22X1 U6598 ( .IN1(n28627), .IN2(n262), .IN3(n28635), .IN4(n305), .Q(n6639)
         );
  OA221X1 U6599 ( .IN1(n28579), .IN2(n348), .IN3(n28587), .IN4(n391), .IN5(
        n6640), .Q(n6635) );
  OA22X1 U6600 ( .IN1(n28595), .IN2(n434), .IN3(n28603), .IN4(n477), .Q(n6640)
         );
  OA221X1 U6601 ( .IN1(n28547), .IN2(n520), .IN3(n28555), .IN4(n563), .IN5(
        n6641), .Q(n6634) );
  OA22X1 U6602 ( .IN1(n28563), .IN2(n606), .IN3(n28571), .IN4(n649), .Q(n6641)
         );
  NAND4X0 U6603 ( .IN1(n6642), .IN2(n6643), .IN3(n6644), .IN4(n6645), .QN(
        n6632) );
  OA221X1 U6604 ( .IN1(n28515), .IN2(n4), .IN3(n28523), .IN4(n47), .IN5(n6646), 
        .Q(n6645) );
  OA22X1 U6605 ( .IN1(n28531), .IN2(n90), .IN3(n28539), .IN4(n133), .Q(n6646)
         );
  OA221X1 U6606 ( .IN1(n28483), .IN2(n176), .IN3(n28491), .IN4(n219), .IN5(
        n6647), .Q(n6644) );
  OA22X1 U6607 ( .IN1(n28499), .IN2(n262), .IN3(n28507), .IN4(n305), .Q(n6647)
         );
  OA221X1 U6608 ( .IN1(n28451), .IN2(n348), .IN3(n28459), .IN4(n391), .IN5(
        n6648), .Q(n6643) );
  OA22X1 U6609 ( .IN1(n28467), .IN2(n434), .IN3(n28475), .IN4(n477), .Q(n6648)
         );
  OA221X1 U6610 ( .IN1(n28419), .IN2(n520), .IN3(n28427), .IN4(n563), .IN5(
        n6649), .Q(n6642) );
  OA22X1 U6611 ( .IN1(n28435), .IN2(n606), .IN3(n28443), .IN4(n649), .Q(n6649)
         );
  NAND4X0 U6612 ( .IN1(n6650), .IN2(n6651), .IN3(n6652), .IN4(n6653), .QN(
        n6630) );
  OA221X1 U6613 ( .IN1(n28387), .IN2(n4), .IN3(n28395), .IN4(n47), .IN5(n6654), 
        .Q(n6653) );
  OA22X1 U6614 ( .IN1(n28403), .IN2(n90), .IN3(n28411), .IN4(n133), .Q(n6654)
         );
  OA221X1 U6615 ( .IN1(n28355), .IN2(n176), .IN3(n28363), .IN4(n219), .IN5(
        n6655), .Q(n6652) );
  OA22X1 U6616 ( .IN1(n28371), .IN2(n262), .IN3(n28379), .IN4(n305), .Q(n6655)
         );
  OA221X1 U6617 ( .IN1(n28323), .IN2(n348), .IN3(n28331), .IN4(n391), .IN5(
        n6656), .Q(n6651) );
  OA22X1 U6618 ( .IN1(n28339), .IN2(n434), .IN3(n28347), .IN4(n477), .Q(n6656)
         );
  OA221X1 U6619 ( .IN1(n28291), .IN2(n520), .IN3(n28299), .IN4(n563), .IN5(
        n6657), .Q(n6650) );
  OA22X1 U6620 ( .IN1(n28307), .IN2(n606), .IN3(n28315), .IN4(n649), .Q(n6657)
         );
  NAND4X0 U6621 ( .IN1(n6658), .IN2(n6659), .IN3(n6660), .IN4(n6661), .QN(
        n6629) );
  OA221X1 U6622 ( .IN1(n28259), .IN2(n4), .IN3(n28267), .IN4(n47), .IN5(n6662), 
        .Q(n6661) );
  OA22X1 U6623 ( .IN1(n28275), .IN2(n90), .IN3(n28283), .IN4(n133), .Q(n6662)
         );
  OA221X1 U6624 ( .IN1(n28227), .IN2(n176), .IN3(n28235), .IN4(n219), .IN5(
        n6663), .Q(n6660) );
  OA22X1 U6625 ( .IN1(n28243), .IN2(n262), .IN3(n28251), .IN4(n305), .Q(n6663)
         );
  OA221X1 U6626 ( .IN1(n28195), .IN2(n348), .IN3(n28203), .IN4(n391), .IN5(
        n6664), .Q(n6659) );
  OA22X1 U6627 ( .IN1(n28211), .IN2(n434), .IN3(n28219), .IN4(n477), .Q(n6664)
         );
  OA221X1 U6628 ( .IN1(n28163), .IN2(n520), .IN3(n28171), .IN4(n563), .IN5(
        n6665), .Q(n6658) );
  OA22X1 U6629 ( .IN1(n28179), .IN2(n606), .IN3(n28187), .IN4(n649), .Q(n6665)
         );
  AO221X1 U6630 ( .IN1(n2246), .IN2(n6666), .IN3(n2248), .IN4(n6667), .IN5(
        n6668), .Q(n6627) );
  AO22X1 U6631 ( .IN1(n2251), .IN2(n6669), .IN3(n2253), .IN4(n6670), .Q(n6668)
         );
  NAND4X0 U6632 ( .IN1(n6671), .IN2(n6672), .IN3(n6673), .IN4(n6674), .QN(
        n6670) );
  OA221X1 U6633 ( .IN1(n28131), .IN2(n4), .IN3(n28139), .IN4(n47), .IN5(n6675), 
        .Q(n6674) );
  OA22X1 U6634 ( .IN1(n28147), .IN2(n90), .IN3(n28155), .IN4(n133), .Q(n6675)
         );
  OA221X1 U6635 ( .IN1(n28099), .IN2(n176), .IN3(n28107), .IN4(n219), .IN5(
        n6676), .Q(n6673) );
  OA22X1 U6636 ( .IN1(n28115), .IN2(n262), .IN3(n28123), .IN4(n305), .Q(n6676)
         );
  OA221X1 U6637 ( .IN1(n28067), .IN2(n348), .IN3(n28075), .IN4(n391), .IN5(
        n6677), .Q(n6672) );
  OA22X1 U6638 ( .IN1(n28083), .IN2(n434), .IN3(n28091), .IN4(n477), .Q(n6677)
         );
  OA221X1 U6639 ( .IN1(n28035), .IN2(n520), .IN3(n28043), .IN4(n563), .IN5(
        n6678), .Q(n6671) );
  OA22X1 U6640 ( .IN1(n28051), .IN2(n606), .IN3(n28059), .IN4(n649), .Q(n6678)
         );
  NAND4X0 U6641 ( .IN1(n6679), .IN2(n6680), .IN3(n6681), .IN4(n6682), .QN(
        n6669) );
  OA221X1 U6642 ( .IN1(n28003), .IN2(n4), .IN3(n28011), .IN4(n47), .IN5(n6683), 
        .Q(n6682) );
  OA22X1 U6643 ( .IN1(n28019), .IN2(n90), .IN3(n28027), .IN4(n133), .Q(n6683)
         );
  OA221X1 U6644 ( .IN1(n27971), .IN2(n176), .IN3(n27979), .IN4(n219), .IN5(
        n6684), .Q(n6681) );
  OA22X1 U6645 ( .IN1(n27987), .IN2(n262), .IN3(n27995), .IN4(n305), .Q(n6684)
         );
  OA221X1 U6646 ( .IN1(n27939), .IN2(n348), .IN3(n27947), .IN4(n391), .IN5(
        n6685), .Q(n6680) );
  OA22X1 U6647 ( .IN1(n27955), .IN2(n434), .IN3(n27963), .IN4(n477), .Q(n6685)
         );
  OA221X1 U6648 ( .IN1(n27907), .IN2(n520), .IN3(n27915), .IN4(n563), .IN5(
        n6686), .Q(n6679) );
  OA22X1 U6649 ( .IN1(n27923), .IN2(n606), .IN3(n27931), .IN4(n649), .Q(n6686)
         );
  NAND4X0 U6650 ( .IN1(n6687), .IN2(n6688), .IN3(n6689), .IN4(n6690), .QN(
        n6667) );
  OA221X1 U6651 ( .IN1(n27875), .IN2(n4), .IN3(n27883), .IN4(n47), .IN5(n6691), 
        .Q(n6690) );
  OA22X1 U6652 ( .IN1(n27891), .IN2(n90), .IN3(n27899), .IN4(n133), .Q(n6691)
         );
  OA221X1 U6653 ( .IN1(n27843), .IN2(n176), .IN3(n27851), .IN4(n219), .IN5(
        n6692), .Q(n6689) );
  OA22X1 U6654 ( .IN1(n27859), .IN2(n262), .IN3(n27867), .IN4(n305), .Q(n6692)
         );
  OA221X1 U6655 ( .IN1(n27811), .IN2(n348), .IN3(n27819), .IN4(n391), .IN5(
        n6693), .Q(n6688) );
  OA22X1 U6656 ( .IN1(n27827), .IN2(n434), .IN3(n27835), .IN4(n477), .Q(n6693)
         );
  OA221X1 U6657 ( .IN1(n27779), .IN2(n520), .IN3(n27787), .IN4(n563), .IN5(
        n6694), .Q(n6687) );
  OA22X1 U6658 ( .IN1(n27795), .IN2(n606), .IN3(n27803), .IN4(n649), .Q(n6694)
         );
  NAND4X0 U6659 ( .IN1(n6695), .IN2(n6696), .IN3(n6697), .IN4(n6698), .QN(
        n6666) );
  OA221X1 U6660 ( .IN1(n27747), .IN2(n4), .IN3(n27755), .IN4(n47), .IN5(n6699), 
        .Q(n6698) );
  OA22X1 U6661 ( .IN1(n27763), .IN2(n90), .IN3(n27771), .IN4(n133), .Q(n6699)
         );
  OA221X1 U6662 ( .IN1(n27715), .IN2(n176), .IN3(n27723), .IN4(n219), .IN5(
        n6700), .Q(n6697) );
  OA22X1 U6663 ( .IN1(n27731), .IN2(n262), .IN3(n27739), .IN4(n305), .Q(n6700)
         );
  OA221X1 U6664 ( .IN1(n27683), .IN2(n348), .IN3(n27691), .IN4(n391), .IN5(
        n6701), .Q(n6696) );
  OA22X1 U6665 ( .IN1(n27699), .IN2(n434), .IN3(n27707), .IN4(n477), .Q(n6701)
         );
  OA221X1 U6666 ( .IN1(n27651), .IN2(n520), .IN3(n27659), .IN4(n563), .IN5(
        n6702), .Q(n6695) );
  OA22X1 U6667 ( .IN1(n27667), .IN2(n606), .IN3(n27675), .IN4(n649), .Q(n6702)
         );
  AO221X1 U6668 ( .IN1(n2287), .IN2(n6703), .IN3(n2289), .IN4(n6704), .IN5(
        n6705), .Q(n6626) );
  AO22X1 U6669 ( .IN1(n2292), .IN2(n6706), .IN3(n2294), .IN4(n6707), .Q(n6705)
         );
  NAND4X0 U6670 ( .IN1(n6708), .IN2(n6709), .IN3(n6710), .IN4(n6711), .QN(
        n6707) );
  OA221X1 U6671 ( .IN1(n29667), .IN2(n4), .IN3(n29675), .IN4(n47), .IN5(n6712), 
        .Q(n6711) );
  OA22X1 U6672 ( .IN1(n29683), .IN2(n90), .IN3(n29691), .IN4(n133), .Q(n6712)
         );
  OA221X1 U6673 ( .IN1(n29635), .IN2(n176), .IN3(n29643), .IN4(n219), .IN5(
        n6713), .Q(n6710) );
  OA22X1 U6674 ( .IN1(n29651), .IN2(n262), .IN3(n29659), .IN4(n305), .Q(n6713)
         );
  OA221X1 U6675 ( .IN1(n29603), .IN2(n348), .IN3(n29611), .IN4(n391), .IN5(
        n6714), .Q(n6709) );
  OA22X1 U6676 ( .IN1(n29619), .IN2(n434), .IN3(n29627), .IN4(n477), .Q(n6714)
         );
  OA221X1 U6677 ( .IN1(n29571), .IN2(n520), .IN3(n29579), .IN4(n563), .IN5(
        n6715), .Q(n6708) );
  OA22X1 U6678 ( .IN1(n29587), .IN2(n606), .IN3(n29595), .IN4(n649), .Q(n6715)
         );
  NAND4X0 U6679 ( .IN1(n6716), .IN2(n6717), .IN3(n6718), .IN4(n6719), .QN(
        n6706) );
  OA221X1 U6680 ( .IN1(n29539), .IN2(n4), .IN3(n29547), .IN4(n47), .IN5(n6720), 
        .Q(n6719) );
  OA22X1 U6681 ( .IN1(n29555), .IN2(n90), .IN3(n29563), .IN4(n133), .Q(n6720)
         );
  OA221X1 U6682 ( .IN1(n29507), .IN2(n176), .IN3(n29515), .IN4(n219), .IN5(
        n6721), .Q(n6718) );
  OA22X1 U6683 ( .IN1(n29523), .IN2(n262), .IN3(n29531), .IN4(n305), .Q(n6721)
         );
  OA221X1 U6684 ( .IN1(n29475), .IN2(n348), .IN3(n29483), .IN4(n391), .IN5(
        n6722), .Q(n6717) );
  OA22X1 U6685 ( .IN1(n29491), .IN2(n434), .IN3(n29499), .IN4(n477), .Q(n6722)
         );
  OA221X1 U6686 ( .IN1(n29443), .IN2(n520), .IN3(n29451), .IN4(n563), .IN5(
        n6723), .Q(n6716) );
  OA22X1 U6687 ( .IN1(n29459), .IN2(n606), .IN3(n29467), .IN4(n649), .Q(n6723)
         );
  NAND4X0 U6688 ( .IN1(n6724), .IN2(n6725), .IN3(n6726), .IN4(n6727), .QN(
        n6704) );
  OA221X1 U6689 ( .IN1(n29411), .IN2(n4), .IN3(n29419), .IN4(n47), .IN5(n6728), 
        .Q(n6727) );
  OA22X1 U6690 ( .IN1(n29427), .IN2(n90), .IN3(n29435), .IN4(n133), .Q(n6728)
         );
  OA221X1 U6691 ( .IN1(n29379), .IN2(n176), .IN3(n29387), .IN4(n219), .IN5(
        n6729), .Q(n6726) );
  OA22X1 U6692 ( .IN1(n29395), .IN2(n262), .IN3(n29403), .IN4(n305), .Q(n6729)
         );
  OA221X1 U6693 ( .IN1(n29347), .IN2(n348), .IN3(n29355), .IN4(n391), .IN5(
        n6730), .Q(n6725) );
  OA22X1 U6694 ( .IN1(n29363), .IN2(n434), .IN3(n29371), .IN4(n477), .Q(n6730)
         );
  OA221X1 U6695 ( .IN1(n29315), .IN2(n520), .IN3(n29323), .IN4(n563), .IN5(
        n6731), .Q(n6724) );
  OA22X1 U6696 ( .IN1(n29331), .IN2(n606), .IN3(n29339), .IN4(n649), .Q(n6731)
         );
  NAND4X0 U6697 ( .IN1(n6732), .IN2(n6733), .IN3(n6734), .IN4(n6735), .QN(
        n6703) );
  OA221X1 U6698 ( .IN1(n29283), .IN2(n4), .IN3(n29291), .IN4(n47), .IN5(n6736), 
        .Q(n6735) );
  OA22X1 U6699 ( .IN1(n29299), .IN2(n90), .IN3(n29307), .IN4(n133), .Q(n6736)
         );
  OA221X1 U6700 ( .IN1(n29251), .IN2(n176), .IN3(n29259), .IN4(n219), .IN5(
        n6737), .Q(n6734) );
  OA22X1 U6701 ( .IN1(n29267), .IN2(n262), .IN3(n29275), .IN4(n305), .Q(n6737)
         );
  OA221X1 U6702 ( .IN1(n29219), .IN2(n348), .IN3(n29227), .IN4(n391), .IN5(
        n6738), .Q(n6733) );
  OA22X1 U6703 ( .IN1(n29235), .IN2(n434), .IN3(n29243), .IN4(n477), .Q(n6738)
         );
  OA221X1 U6704 ( .IN1(n29187), .IN2(n520), .IN3(n29195), .IN4(n563), .IN5(
        n6739), .Q(n6732) );
  OA22X1 U6705 ( .IN1(n29203), .IN2(n606), .IN3(n29211), .IN4(n649), .Q(n6739)
         );
  AO221X1 U6706 ( .IN1(n2328), .IN2(n6740), .IN3(n2330), .IN4(n6741), .IN5(
        n6742), .Q(n6625) );
  AO22X1 U6707 ( .IN1(n2333), .IN2(n6743), .IN3(n2335), .IN4(n6744), .Q(n6742)
         );
  NAND4X0 U6708 ( .IN1(n6745), .IN2(n6746), .IN3(n6747), .IN4(n6748), .QN(
        n6744) );
  OA221X1 U6709 ( .IN1(n29155), .IN2(n3), .IN3(n29163), .IN4(n46), .IN5(n6749), 
        .Q(n6748) );
  OA22X1 U6710 ( .IN1(n29171), .IN2(n89), .IN3(n29179), .IN4(n132), .Q(n6749)
         );
  OA221X1 U6711 ( .IN1(n29123), .IN2(n175), .IN3(n29131), .IN4(n218), .IN5(
        n6750), .Q(n6747) );
  OA22X1 U6712 ( .IN1(n29139), .IN2(n261), .IN3(n29147), .IN4(n304), .Q(n6750)
         );
  OA221X1 U6713 ( .IN1(n29091), .IN2(n347), .IN3(n29099), .IN4(n390), .IN5(
        n6751), .Q(n6746) );
  OA22X1 U6714 ( .IN1(n29107), .IN2(n433), .IN3(n29115), .IN4(n476), .Q(n6751)
         );
  OA221X1 U6715 ( .IN1(n29059), .IN2(n519), .IN3(n29067), .IN4(n562), .IN5(
        n6752), .Q(n6745) );
  OA22X1 U6716 ( .IN1(n29075), .IN2(n605), .IN3(n29083), .IN4(n648), .Q(n6752)
         );
  NAND4X0 U6717 ( .IN1(n6753), .IN2(n6754), .IN3(n6755), .IN4(n6756), .QN(
        n6743) );
  OA221X1 U6718 ( .IN1(n29027), .IN2(n3), .IN3(n29035), .IN4(n46), .IN5(n6757), 
        .Q(n6756) );
  OA22X1 U6719 ( .IN1(n29043), .IN2(n89), .IN3(n29051), .IN4(n132), .Q(n6757)
         );
  OA221X1 U6720 ( .IN1(n28995), .IN2(n175), .IN3(n29003), .IN4(n218), .IN5(
        n6758), .Q(n6755) );
  OA22X1 U6721 ( .IN1(n29011), .IN2(n261), .IN3(n29019), .IN4(n304), .Q(n6758)
         );
  OA221X1 U6722 ( .IN1(n28963), .IN2(n347), .IN3(n28971), .IN4(n390), .IN5(
        n6759), .Q(n6754) );
  OA22X1 U6723 ( .IN1(n28979), .IN2(n433), .IN3(n28987), .IN4(n476), .Q(n6759)
         );
  OA221X1 U6724 ( .IN1(n28931), .IN2(n519), .IN3(n28939), .IN4(n562), .IN5(
        n6760), .Q(n6753) );
  OA22X1 U6725 ( .IN1(n28947), .IN2(n605), .IN3(n28955), .IN4(n648), .Q(n6760)
         );
  NAND4X0 U6726 ( .IN1(n6761), .IN2(n6762), .IN3(n6763), .IN4(n6764), .QN(
        n6741) );
  OA221X1 U6727 ( .IN1(n28899), .IN2(n3), .IN3(n28907), .IN4(n46), .IN5(n6765), 
        .Q(n6764) );
  OA22X1 U6728 ( .IN1(n28915), .IN2(n89), .IN3(n28923), .IN4(n132), .Q(n6765)
         );
  OA221X1 U6729 ( .IN1(n28867), .IN2(n175), .IN3(n28875), .IN4(n218), .IN5(
        n6766), .Q(n6763) );
  OA22X1 U6730 ( .IN1(n28883), .IN2(n261), .IN3(n28891), .IN4(n304), .Q(n6766)
         );
  OA221X1 U6731 ( .IN1(n28835), .IN2(n347), .IN3(n28843), .IN4(n390), .IN5(
        n6767), .Q(n6762) );
  OA22X1 U6732 ( .IN1(n28851), .IN2(n433), .IN3(n28859), .IN4(n476), .Q(n6767)
         );
  OA221X1 U6733 ( .IN1(n28803), .IN2(n519), .IN3(n28811), .IN4(n562), .IN5(
        n6768), .Q(n6761) );
  OA22X1 U6734 ( .IN1(n28819), .IN2(n605), .IN3(n28827), .IN4(n648), .Q(n6768)
         );
  NAND4X0 U6735 ( .IN1(n6769), .IN2(n6770), .IN3(n6771), .IN4(n6772), .QN(
        n6740) );
  OA221X1 U6736 ( .IN1(n28771), .IN2(n3), .IN3(n28779), .IN4(n46), .IN5(n6773), 
        .Q(n6772) );
  OA22X1 U6737 ( .IN1(n28787), .IN2(n89), .IN3(n28795), .IN4(n132), .Q(n6773)
         );
  OA221X1 U6738 ( .IN1(n28739), .IN2(n175), .IN3(n28747), .IN4(n218), .IN5(
        n6774), .Q(n6771) );
  OA22X1 U6739 ( .IN1(n28755), .IN2(n261), .IN3(n28763), .IN4(n304), .Q(n6774)
         );
  OA221X1 U6740 ( .IN1(n28707), .IN2(n347), .IN3(n28715), .IN4(n390), .IN5(
        n6775), .Q(n6770) );
  OA22X1 U6741 ( .IN1(n28723), .IN2(n433), .IN3(n28731), .IN4(n476), .Q(n6775)
         );
  OA221X1 U6742 ( .IN1(n28675), .IN2(n519), .IN3(n28683), .IN4(n562), .IN5(
        n6776), .Q(n6769) );
  OA22X1 U6743 ( .IN1(n28691), .IN2(n605), .IN3(n28699), .IN4(n648), .Q(n6776)
         );
  OR4X1 U6744 ( .IN1(n6777), .IN2(n6778), .IN3(n6779), .IN4(n6780), .Q(n2172)
         );
  AO221X1 U6745 ( .IN1(n2157), .IN2(n6781), .IN3(n2159), .IN4(n6782), .IN5(
        n6783), .Q(n6780) );
  AO22X1 U6746 ( .IN1(n2162), .IN2(n6784), .IN3(n2164), .IN4(n6785), .Q(n6783)
         );
  NAND4X0 U6747 ( .IN1(n6786), .IN2(n6787), .IN3(n6788), .IN4(n6789), .QN(
        n6785) );
  OA221X1 U6748 ( .IN1(n28642), .IN2(n3), .IN3(n28650), .IN4(n46), .IN5(n6790), 
        .Q(n6789) );
  OA22X1 U6749 ( .IN1(n28658), .IN2(n89), .IN3(n28666), .IN4(n132), .Q(n6790)
         );
  OA221X1 U6750 ( .IN1(n28610), .IN2(n175), .IN3(n28618), .IN4(n218), .IN5(
        n6791), .Q(n6788) );
  OA22X1 U6751 ( .IN1(n28626), .IN2(n261), .IN3(n28634), .IN4(n304), .Q(n6791)
         );
  OA221X1 U6752 ( .IN1(n28578), .IN2(n347), .IN3(n28586), .IN4(n390), .IN5(
        n6792), .Q(n6787) );
  OA22X1 U6753 ( .IN1(n28594), .IN2(n433), .IN3(n28602), .IN4(n476), .Q(n6792)
         );
  OA221X1 U6754 ( .IN1(n28546), .IN2(n519), .IN3(n28554), .IN4(n562), .IN5(
        n6793), .Q(n6786) );
  OA22X1 U6755 ( .IN1(n28562), .IN2(n605), .IN3(n28570), .IN4(n648), .Q(n6793)
         );
  NAND4X0 U6756 ( .IN1(n6794), .IN2(n6795), .IN3(n6796), .IN4(n6797), .QN(
        n6784) );
  OA221X1 U6757 ( .IN1(n28514), .IN2(n3), .IN3(n28522), .IN4(n46), .IN5(n6798), 
        .Q(n6797) );
  OA22X1 U6758 ( .IN1(n28530), .IN2(n89), .IN3(n28538), .IN4(n132), .Q(n6798)
         );
  OA221X1 U6759 ( .IN1(n28482), .IN2(n175), .IN3(n28490), .IN4(n218), .IN5(
        n6799), .Q(n6796) );
  OA22X1 U6760 ( .IN1(n28498), .IN2(n261), .IN3(n28506), .IN4(n304), .Q(n6799)
         );
  OA221X1 U6761 ( .IN1(n28450), .IN2(n347), .IN3(n28458), .IN4(n390), .IN5(
        n6800), .Q(n6795) );
  OA22X1 U6762 ( .IN1(n28466), .IN2(n433), .IN3(n28474), .IN4(n476), .Q(n6800)
         );
  OA221X1 U6763 ( .IN1(n28418), .IN2(n519), .IN3(n28426), .IN4(n562), .IN5(
        n6801), .Q(n6794) );
  OA22X1 U6764 ( .IN1(n28434), .IN2(n605), .IN3(n28442), .IN4(n648), .Q(n6801)
         );
  NAND4X0 U6765 ( .IN1(n6802), .IN2(n6803), .IN3(n6804), .IN4(n6805), .QN(
        n6782) );
  OA221X1 U6766 ( .IN1(n28386), .IN2(n3), .IN3(n28394), .IN4(n46), .IN5(n6806), 
        .Q(n6805) );
  OA22X1 U6767 ( .IN1(n28402), .IN2(n89), .IN3(n28410), .IN4(n132), .Q(n6806)
         );
  OA221X1 U6768 ( .IN1(n28354), .IN2(n175), .IN3(n28362), .IN4(n218), .IN5(
        n6807), .Q(n6804) );
  OA22X1 U6769 ( .IN1(n28370), .IN2(n261), .IN3(n28378), .IN4(n304), .Q(n6807)
         );
  OA221X1 U6770 ( .IN1(n28322), .IN2(n347), .IN3(n28330), .IN4(n390), .IN5(
        n6808), .Q(n6803) );
  OA22X1 U6771 ( .IN1(n28338), .IN2(n433), .IN3(n28346), .IN4(n476), .Q(n6808)
         );
  OA221X1 U6772 ( .IN1(n28290), .IN2(n519), .IN3(n28298), .IN4(n562), .IN5(
        n6809), .Q(n6802) );
  OA22X1 U6773 ( .IN1(n28306), .IN2(n605), .IN3(n28314), .IN4(n648), .Q(n6809)
         );
  NAND4X0 U6774 ( .IN1(n6810), .IN2(n6811), .IN3(n6812), .IN4(n6813), .QN(
        n6781) );
  OA221X1 U6775 ( .IN1(n28258), .IN2(n3), .IN3(n28266), .IN4(n46), .IN5(n6814), 
        .Q(n6813) );
  OA22X1 U6776 ( .IN1(n28274), .IN2(n89), .IN3(n28282), .IN4(n132), .Q(n6814)
         );
  OA221X1 U6777 ( .IN1(n28226), .IN2(n175), .IN3(n28234), .IN4(n218), .IN5(
        n6815), .Q(n6812) );
  OA22X1 U6778 ( .IN1(n28242), .IN2(n261), .IN3(n28250), .IN4(n304), .Q(n6815)
         );
  OA221X1 U6779 ( .IN1(n28194), .IN2(n347), .IN3(n28202), .IN4(n390), .IN5(
        n6816), .Q(n6811) );
  OA22X1 U6780 ( .IN1(n28210), .IN2(n433), .IN3(n28218), .IN4(n476), .Q(n6816)
         );
  OA221X1 U6781 ( .IN1(n28162), .IN2(n519), .IN3(n28170), .IN4(n562), .IN5(
        n6817), .Q(n6810) );
  OA22X1 U6782 ( .IN1(n28178), .IN2(n605), .IN3(n28186), .IN4(n648), .Q(n6817)
         );
  AO221X1 U6783 ( .IN1(n2246), .IN2(n6818), .IN3(n2248), .IN4(n6819), .IN5(
        n6820), .Q(n6779) );
  AO22X1 U6784 ( .IN1(n2251), .IN2(n6821), .IN3(n2253), .IN4(n6822), .Q(n6820)
         );
  NAND4X0 U6785 ( .IN1(n6823), .IN2(n6824), .IN3(n6825), .IN4(n6826), .QN(
        n6822) );
  OA221X1 U6786 ( .IN1(n28130), .IN2(n3), .IN3(n28138), .IN4(n46), .IN5(n6827), 
        .Q(n6826) );
  OA22X1 U6787 ( .IN1(n28146), .IN2(n89), .IN3(n28154), .IN4(n132), .Q(n6827)
         );
  OA221X1 U6788 ( .IN1(n28098), .IN2(n175), .IN3(n28106), .IN4(n218), .IN5(
        n6828), .Q(n6825) );
  OA22X1 U6789 ( .IN1(n28114), .IN2(n261), .IN3(n28122), .IN4(n304), .Q(n6828)
         );
  OA221X1 U6790 ( .IN1(n28066), .IN2(n347), .IN3(n28074), .IN4(n390), .IN5(
        n6829), .Q(n6824) );
  OA22X1 U6791 ( .IN1(n28082), .IN2(n433), .IN3(n28090), .IN4(n476), .Q(n6829)
         );
  OA221X1 U6792 ( .IN1(n28034), .IN2(n519), .IN3(n28042), .IN4(n562), .IN5(
        n6830), .Q(n6823) );
  OA22X1 U6793 ( .IN1(n28050), .IN2(n605), .IN3(n28058), .IN4(n648), .Q(n6830)
         );
  NAND4X0 U6794 ( .IN1(n6831), .IN2(n6832), .IN3(n6833), .IN4(n6834), .QN(
        n6821) );
  OA221X1 U6795 ( .IN1(n28002), .IN2(n3), .IN3(n28010), .IN4(n46), .IN5(n6835), 
        .Q(n6834) );
  OA22X1 U6796 ( .IN1(n28018), .IN2(n89), .IN3(n28026), .IN4(n132), .Q(n6835)
         );
  OA221X1 U6797 ( .IN1(n27970), .IN2(n175), .IN3(n27978), .IN4(n218), .IN5(
        n6836), .Q(n6833) );
  OA22X1 U6798 ( .IN1(n27986), .IN2(n261), .IN3(n27994), .IN4(n304), .Q(n6836)
         );
  OA221X1 U6799 ( .IN1(n27938), .IN2(n347), .IN3(n27946), .IN4(n390), .IN5(
        n6837), .Q(n6832) );
  OA22X1 U6800 ( .IN1(n27954), .IN2(n433), .IN3(n27962), .IN4(n476), .Q(n6837)
         );
  OA221X1 U6801 ( .IN1(n27906), .IN2(n519), .IN3(n27914), .IN4(n562), .IN5(
        n6838), .Q(n6831) );
  OA22X1 U6802 ( .IN1(n27922), .IN2(n605), .IN3(n27930), .IN4(n648), .Q(n6838)
         );
  NAND4X0 U6803 ( .IN1(n6839), .IN2(n6840), .IN3(n6841), .IN4(n6842), .QN(
        n6819) );
  OA221X1 U6804 ( .IN1(n27874), .IN2(n3), .IN3(n27882), .IN4(n46), .IN5(n6843), 
        .Q(n6842) );
  OA22X1 U6805 ( .IN1(n27890), .IN2(n89), .IN3(n27898), .IN4(n132), .Q(n6843)
         );
  OA221X1 U6806 ( .IN1(n27842), .IN2(n175), .IN3(n27850), .IN4(n218), .IN5(
        n6844), .Q(n6841) );
  OA22X1 U6807 ( .IN1(n27858), .IN2(n261), .IN3(n27866), .IN4(n304), .Q(n6844)
         );
  OA221X1 U6808 ( .IN1(n27810), .IN2(n347), .IN3(n27818), .IN4(n390), .IN5(
        n6845), .Q(n6840) );
  OA22X1 U6809 ( .IN1(n27826), .IN2(n433), .IN3(n27834), .IN4(n476), .Q(n6845)
         );
  OA221X1 U6810 ( .IN1(n27778), .IN2(n519), .IN3(n27786), .IN4(n562), .IN5(
        n6846), .Q(n6839) );
  OA22X1 U6811 ( .IN1(n27794), .IN2(n605), .IN3(n27802), .IN4(n648), .Q(n6846)
         );
  NAND4X0 U6812 ( .IN1(n6847), .IN2(n6848), .IN3(n6849), .IN4(n6850), .QN(
        n6818) );
  OA221X1 U6813 ( .IN1(n27746), .IN2(n3), .IN3(n27754), .IN4(n46), .IN5(n6851), 
        .Q(n6850) );
  OA22X1 U6814 ( .IN1(n27762), .IN2(n89), .IN3(n27770), .IN4(n132), .Q(n6851)
         );
  OA221X1 U6815 ( .IN1(n27714), .IN2(n175), .IN3(n27722), .IN4(n218), .IN5(
        n6852), .Q(n6849) );
  OA22X1 U6816 ( .IN1(n27730), .IN2(n261), .IN3(n27738), .IN4(n304), .Q(n6852)
         );
  OA221X1 U6817 ( .IN1(n27682), .IN2(n347), .IN3(n27690), .IN4(n390), .IN5(
        n6853), .Q(n6848) );
  OA22X1 U6818 ( .IN1(n27698), .IN2(n433), .IN3(n27706), .IN4(n476), .Q(n6853)
         );
  OA221X1 U6819 ( .IN1(n27650), .IN2(n519), .IN3(n27658), .IN4(n562), .IN5(
        n6854), .Q(n6847) );
  OA22X1 U6820 ( .IN1(n27666), .IN2(n605), .IN3(n27674), .IN4(n648), .Q(n6854)
         );
  AO221X1 U6821 ( .IN1(n2287), .IN2(n6855), .IN3(n2289), .IN4(n6856), .IN5(
        n6857), .Q(n6778) );
  AO22X1 U6822 ( .IN1(n2292), .IN2(n6858), .IN3(n2294), .IN4(n6859), .Q(n6857)
         );
  NAND4X0 U6823 ( .IN1(n6860), .IN2(n6861), .IN3(n6862), .IN4(n6863), .QN(
        n6859) );
  OA221X1 U6824 ( .IN1(n29666), .IN2(n2), .IN3(n29674), .IN4(n45), .IN5(n6864), 
        .Q(n6863) );
  OA22X1 U6825 ( .IN1(n29682), .IN2(n88), .IN3(n29690), .IN4(n131), .Q(n6864)
         );
  OA221X1 U6826 ( .IN1(n29634), .IN2(n174), .IN3(n29642), .IN4(n217), .IN5(
        n6865), .Q(n6862) );
  OA22X1 U6827 ( .IN1(n29650), .IN2(n260), .IN3(n29658), .IN4(n303), .Q(n6865)
         );
  OA221X1 U6828 ( .IN1(n29602), .IN2(n346), .IN3(n29610), .IN4(n389), .IN5(
        n6866), .Q(n6861) );
  OA22X1 U6829 ( .IN1(n29618), .IN2(n432), .IN3(n29626), .IN4(n475), .Q(n6866)
         );
  OA221X1 U6830 ( .IN1(n29570), .IN2(n518), .IN3(n29578), .IN4(n561), .IN5(
        n6867), .Q(n6860) );
  OA22X1 U6831 ( .IN1(n29586), .IN2(n604), .IN3(n29594), .IN4(n647), .Q(n6867)
         );
  NAND4X0 U6832 ( .IN1(n6868), .IN2(n6869), .IN3(n6870), .IN4(n6871), .QN(
        n6858) );
  OA221X1 U6833 ( .IN1(n29538), .IN2(n2), .IN3(n29546), .IN4(n45), .IN5(n6872), 
        .Q(n6871) );
  OA22X1 U6834 ( .IN1(n29554), .IN2(n88), .IN3(n29562), .IN4(n131), .Q(n6872)
         );
  OA221X1 U6835 ( .IN1(n29506), .IN2(n174), .IN3(n29514), .IN4(n217), .IN5(
        n6873), .Q(n6870) );
  OA22X1 U6836 ( .IN1(n29522), .IN2(n260), .IN3(n29530), .IN4(n303), .Q(n6873)
         );
  OA221X1 U6837 ( .IN1(n29474), .IN2(n346), .IN3(n29482), .IN4(n389), .IN5(
        n6874), .Q(n6869) );
  OA22X1 U6838 ( .IN1(n29490), .IN2(n432), .IN3(n29498), .IN4(n475), .Q(n6874)
         );
  OA221X1 U6839 ( .IN1(n29442), .IN2(n518), .IN3(n29450), .IN4(n561), .IN5(
        n6875), .Q(n6868) );
  OA22X1 U6840 ( .IN1(n29458), .IN2(n604), .IN3(n29466), .IN4(n647), .Q(n6875)
         );
  NAND4X0 U6841 ( .IN1(n6876), .IN2(n6877), .IN3(n6878), .IN4(n6879), .QN(
        n6856) );
  OA221X1 U6842 ( .IN1(n29410), .IN2(n2), .IN3(n29418), .IN4(n45), .IN5(n6880), 
        .Q(n6879) );
  OA22X1 U6843 ( .IN1(n29426), .IN2(n88), .IN3(n29434), .IN4(n131), .Q(n6880)
         );
  OA221X1 U6844 ( .IN1(n29378), .IN2(n174), .IN3(n29386), .IN4(n217), .IN5(
        n6881), .Q(n6878) );
  OA22X1 U6845 ( .IN1(n29394), .IN2(n260), .IN3(n29402), .IN4(n303), .Q(n6881)
         );
  OA221X1 U6846 ( .IN1(n29346), .IN2(n346), .IN3(n29354), .IN4(n389), .IN5(
        n6882), .Q(n6877) );
  OA22X1 U6847 ( .IN1(n29362), .IN2(n432), .IN3(n29370), .IN4(n475), .Q(n6882)
         );
  OA221X1 U6848 ( .IN1(n29314), .IN2(n518), .IN3(n29322), .IN4(n561), .IN5(
        n6883), .Q(n6876) );
  OA22X1 U6849 ( .IN1(n29330), .IN2(n604), .IN3(n29338), .IN4(n647), .Q(n6883)
         );
  NAND4X0 U6850 ( .IN1(n6884), .IN2(n6885), .IN3(n6886), .IN4(n6887), .QN(
        n6855) );
  OA221X1 U6851 ( .IN1(n29282), .IN2(n2), .IN3(n29290), .IN4(n45), .IN5(n6888), 
        .Q(n6887) );
  OA22X1 U6852 ( .IN1(n29298), .IN2(n88), .IN3(n29306), .IN4(n131), .Q(n6888)
         );
  OA221X1 U6853 ( .IN1(n29250), .IN2(n174), .IN3(n29258), .IN4(n217), .IN5(
        n6889), .Q(n6886) );
  OA22X1 U6854 ( .IN1(n29266), .IN2(n260), .IN3(n29274), .IN4(n303), .Q(n6889)
         );
  OA221X1 U6855 ( .IN1(n29218), .IN2(n346), .IN3(n29226), .IN4(n389), .IN5(
        n6890), .Q(n6885) );
  OA22X1 U6856 ( .IN1(n29234), .IN2(n432), .IN3(n29242), .IN4(n475), .Q(n6890)
         );
  OA221X1 U6857 ( .IN1(n29186), .IN2(n518), .IN3(n29194), .IN4(n561), .IN5(
        n6891), .Q(n6884) );
  OA22X1 U6858 ( .IN1(n29202), .IN2(n604), .IN3(n29210), .IN4(n647), .Q(n6891)
         );
  AO221X1 U6859 ( .IN1(n2328), .IN2(n6892), .IN3(n2330), .IN4(n6893), .IN5(
        n6894), .Q(n6777) );
  AO22X1 U6860 ( .IN1(n2333), .IN2(n6895), .IN3(n2335), .IN4(n6896), .Q(n6894)
         );
  NAND4X0 U6861 ( .IN1(n6897), .IN2(n6898), .IN3(n6899), .IN4(n6900), .QN(
        n6896) );
  OA221X1 U6862 ( .IN1(n29154), .IN2(n2), .IN3(n29162), .IN4(n45), .IN5(n6901), 
        .Q(n6900) );
  OA22X1 U6863 ( .IN1(n29170), .IN2(n88), .IN3(n29178), .IN4(n131), .Q(n6901)
         );
  OA221X1 U6864 ( .IN1(n29122), .IN2(n174), .IN3(n29130), .IN4(n217), .IN5(
        n6902), .Q(n6899) );
  OA22X1 U6865 ( .IN1(n29138), .IN2(n260), .IN3(n29146), .IN4(n303), .Q(n6902)
         );
  OA221X1 U6866 ( .IN1(n29090), .IN2(n346), .IN3(n29098), .IN4(n389), .IN5(
        n6903), .Q(n6898) );
  OA22X1 U6867 ( .IN1(n29106), .IN2(n432), .IN3(n29114), .IN4(n475), .Q(n6903)
         );
  OA221X1 U6868 ( .IN1(n29058), .IN2(n518), .IN3(n29066), .IN4(n561), .IN5(
        n6904), .Q(n6897) );
  OA22X1 U6869 ( .IN1(n29074), .IN2(n604), .IN3(n29082), .IN4(n647), .Q(n6904)
         );
  NAND4X0 U6870 ( .IN1(n6905), .IN2(n6906), .IN3(n6907), .IN4(n6908), .QN(
        n6895) );
  OA221X1 U6871 ( .IN1(n29026), .IN2(n2), .IN3(n29034), .IN4(n45), .IN5(n6909), 
        .Q(n6908) );
  OA22X1 U6872 ( .IN1(n29042), .IN2(n88), .IN3(n29050), .IN4(n131), .Q(n6909)
         );
  OA221X1 U6873 ( .IN1(n28994), .IN2(n174), .IN3(n29002), .IN4(n217), .IN5(
        n6910), .Q(n6907) );
  OA22X1 U6874 ( .IN1(n29010), .IN2(n260), .IN3(n29018), .IN4(n303), .Q(n6910)
         );
  OA221X1 U6875 ( .IN1(n28962), .IN2(n346), .IN3(n28970), .IN4(n389), .IN5(
        n6911), .Q(n6906) );
  OA22X1 U6876 ( .IN1(n28978), .IN2(n432), .IN3(n28986), .IN4(n475), .Q(n6911)
         );
  OA221X1 U6877 ( .IN1(n28930), .IN2(n518), .IN3(n28938), .IN4(n561), .IN5(
        n6912), .Q(n6905) );
  OA22X1 U6878 ( .IN1(n28946), .IN2(n604), .IN3(n28954), .IN4(n647), .Q(n6912)
         );
  NAND4X0 U6879 ( .IN1(n6913), .IN2(n6914), .IN3(n6915), .IN4(n6916), .QN(
        n6893) );
  OA221X1 U6880 ( .IN1(n28898), .IN2(n2), .IN3(n28906), .IN4(n45), .IN5(n6917), 
        .Q(n6916) );
  OA22X1 U6881 ( .IN1(n28914), .IN2(n88), .IN3(n28922), .IN4(n131), .Q(n6917)
         );
  OA221X1 U6882 ( .IN1(n28866), .IN2(n174), .IN3(n28874), .IN4(n217), .IN5(
        n6918), .Q(n6915) );
  OA22X1 U6883 ( .IN1(n28882), .IN2(n260), .IN3(n28890), .IN4(n303), .Q(n6918)
         );
  OA221X1 U6884 ( .IN1(n28834), .IN2(n346), .IN3(n28842), .IN4(n389), .IN5(
        n6919), .Q(n6914) );
  OA22X1 U6885 ( .IN1(n28850), .IN2(n432), .IN3(n28858), .IN4(n475), .Q(n6919)
         );
  OA221X1 U6886 ( .IN1(n28802), .IN2(n518), .IN3(n28810), .IN4(n561), .IN5(
        n6920), .Q(n6913) );
  OA22X1 U6887 ( .IN1(n28818), .IN2(n604), .IN3(n28826), .IN4(n647), .Q(n6920)
         );
  NAND4X0 U6888 ( .IN1(n6921), .IN2(n6922), .IN3(n6923), .IN4(n6924), .QN(
        n6892) );
  OA221X1 U6889 ( .IN1(n28770), .IN2(n2), .IN3(n28778), .IN4(n45), .IN5(n6925), 
        .Q(n6924) );
  OA22X1 U6890 ( .IN1(n28786), .IN2(n88), .IN3(n28794), .IN4(n131), .Q(n6925)
         );
  OA221X1 U6891 ( .IN1(n28738), .IN2(n174), .IN3(n28746), .IN4(n217), .IN5(
        n6926), .Q(n6923) );
  OA22X1 U6892 ( .IN1(n28754), .IN2(n260), .IN3(n28762), .IN4(n303), .Q(n6926)
         );
  OA221X1 U6893 ( .IN1(n28706), .IN2(n346), .IN3(n28714), .IN4(n389), .IN5(
        n6927), .Q(n6922) );
  OA22X1 U6894 ( .IN1(n28722), .IN2(n432), .IN3(n28730), .IN4(n475), .Q(n6927)
         );
  OA221X1 U6895 ( .IN1(n28674), .IN2(n518), .IN3(n28682), .IN4(n561), .IN5(
        n6928), .Q(n6921) );
  OA22X1 U6896 ( .IN1(n28690), .IN2(n604), .IN3(n28698), .IN4(n647), .Q(n6928)
         );
  OR4X1 U6897 ( .IN1(n6929), .IN2(n6930), .IN3(n6931), .IN4(n6932), .Q(n2171)
         );
  AO221X1 U6898 ( .IN1(n2157), .IN2(n6933), .IN3(n2159), .IN4(n6934), .IN5(
        n6935), .Q(n6932) );
  AO22X1 U6899 ( .IN1(n2162), .IN2(n6936), .IN3(n2164), .IN4(n6937), .Q(n6935)
         );
  NAND4X0 U6900 ( .IN1(n6938), .IN2(n6939), .IN3(n6940), .IN4(n6941), .QN(
        n6937) );
  OA221X1 U6901 ( .IN1(n28641), .IN2(n2), .IN3(n28649), .IN4(n45), .IN5(n6942), 
        .Q(n6941) );
  OA22X1 U6902 ( .IN1(n28657), .IN2(n88), .IN3(n28665), .IN4(n131), .Q(n6942)
         );
  OA221X1 U6903 ( .IN1(n28609), .IN2(n174), .IN3(n28617), .IN4(n217), .IN5(
        n6943), .Q(n6940) );
  OA22X1 U6904 ( .IN1(n28625), .IN2(n260), .IN3(n28633), .IN4(n303), .Q(n6943)
         );
  OA221X1 U6905 ( .IN1(n28577), .IN2(n346), .IN3(n28585), .IN4(n389), .IN5(
        n6944), .Q(n6939) );
  OA22X1 U6906 ( .IN1(n28593), .IN2(n432), .IN3(n28601), .IN4(n475), .Q(n6944)
         );
  OA221X1 U6907 ( .IN1(n28545), .IN2(n518), .IN3(n28553), .IN4(n561), .IN5(
        n6945), .Q(n6938) );
  OA22X1 U6908 ( .IN1(n28561), .IN2(n604), .IN3(n28569), .IN4(n647), .Q(n6945)
         );
  AND3X1 U6909 ( .IN1(n6946), .IN2(n6947), .IN3(n6948), .Q(n2164) );
  NAND4X0 U6910 ( .IN1(n6949), .IN2(n6950), .IN3(n6951), .IN4(n6952), .QN(
        n6936) );
  OA221X1 U6911 ( .IN1(n28513), .IN2(n2), .IN3(n28521), .IN4(n45), .IN5(n6953), 
        .Q(n6952) );
  OA22X1 U6912 ( .IN1(n28529), .IN2(n88), .IN3(n28537), .IN4(n131), .Q(n6953)
         );
  OA221X1 U6913 ( .IN1(n28481), .IN2(n174), .IN3(n28489), .IN4(n217), .IN5(
        n6954), .Q(n6951) );
  OA22X1 U6914 ( .IN1(n28497), .IN2(n260), .IN3(n28505), .IN4(n303), .Q(n6954)
         );
  OA221X1 U6915 ( .IN1(n28449), .IN2(n346), .IN3(n28457), .IN4(n389), .IN5(
        n6955), .Q(n6950) );
  OA22X1 U6916 ( .IN1(n28465), .IN2(n432), .IN3(n28473), .IN4(n475), .Q(n6955)
         );
  OA221X1 U6917 ( .IN1(n28417), .IN2(n518), .IN3(n28425), .IN4(n561), .IN5(
        n6956), .Q(n6949) );
  OA22X1 U6918 ( .IN1(n28433), .IN2(n604), .IN3(n28441), .IN4(n647), .Q(n6956)
         );
  AND3X1 U6919 ( .IN1(n6957), .IN2(n6947), .IN3(n6948), .Q(n2162) );
  NAND4X0 U6920 ( .IN1(n6958), .IN2(n6959), .IN3(n6960), .IN4(n6961), .QN(
        n6934) );
  OA221X1 U6921 ( .IN1(n28385), .IN2(n2), .IN3(n28393), .IN4(n45), .IN5(n6962), 
        .Q(n6961) );
  OA22X1 U6922 ( .IN1(n28401), .IN2(n88), .IN3(n28409), .IN4(n131), .Q(n6962)
         );
  OA221X1 U6923 ( .IN1(n28353), .IN2(n174), .IN3(n28361), .IN4(n217), .IN5(
        n6963), .Q(n6960) );
  OA22X1 U6924 ( .IN1(n28369), .IN2(n260), .IN3(n28377), .IN4(n303), .Q(n6963)
         );
  OA221X1 U6925 ( .IN1(n28321), .IN2(n346), .IN3(n28329), .IN4(n389), .IN5(
        n6964), .Q(n6959) );
  OA22X1 U6926 ( .IN1(n28337), .IN2(n432), .IN3(n28345), .IN4(n475), .Q(n6964)
         );
  OA221X1 U6927 ( .IN1(n28289), .IN2(n518), .IN3(n28297), .IN4(n561), .IN5(
        n6965), .Q(n6958) );
  OA22X1 U6928 ( .IN1(n28305), .IN2(n604), .IN3(n28313), .IN4(n647), .Q(n6965)
         );
  AND2X1 U6929 ( .IN1(n6966), .IN2(n6946), .Q(n2159) );
  NAND4X0 U6930 ( .IN1(n6967), .IN2(n6968), .IN3(n6969), .IN4(n6970), .QN(
        n6933) );
  OA221X1 U6931 ( .IN1(n28257), .IN2(n2), .IN3(n28265), .IN4(n45), .IN5(n6971), 
        .Q(n6970) );
  OA22X1 U6932 ( .IN1(n28273), .IN2(n88), .IN3(n28281), .IN4(n131), .Q(n6971)
         );
  OA221X1 U6933 ( .IN1(n28225), .IN2(n174), .IN3(n28233), .IN4(n217), .IN5(
        n6972), .Q(n6969) );
  OA22X1 U6934 ( .IN1(n28241), .IN2(n260), .IN3(n28249), .IN4(n303), .Q(n6972)
         );
  OA221X1 U6935 ( .IN1(n28193), .IN2(n346), .IN3(n28201), .IN4(n389), .IN5(
        n6973), .Q(n6968) );
  OA22X1 U6936 ( .IN1(n28209), .IN2(n432), .IN3(n28217), .IN4(n475), .Q(n6973)
         );
  OA221X1 U6937 ( .IN1(n28161), .IN2(n518), .IN3(n28169), .IN4(n561), .IN5(
        n6974), .Q(n6967) );
  OA22X1 U6938 ( .IN1(n28177), .IN2(n604), .IN3(n28185), .IN4(n647), .Q(n6974)
         );
  AND2X1 U6939 ( .IN1(n6966), .IN2(n6957), .Q(n2157) );
  AO221X1 U6940 ( .IN1(n2246), .IN2(n6975), .IN3(n2248), .IN4(n6976), .IN5(
        n6977), .Q(n6931) );
  AO22X1 U6941 ( .IN1(n2251), .IN2(n6978), .IN3(n2253), .IN4(n6979), .Q(n6977)
         );
  NAND4X0 U6942 ( .IN1(n6980), .IN2(n6981), .IN3(n6982), .IN4(n6983), .QN(
        n6979) );
  OA221X1 U6943 ( .IN1(n28129), .IN2(n1), .IN3(n28137), .IN4(n44), .IN5(n6984), 
        .Q(n6983) );
  OA22X1 U6944 ( .IN1(n28145), .IN2(n87), .IN3(n28153), .IN4(n130), .Q(n6984)
         );
  OA221X1 U6945 ( .IN1(n28097), .IN2(n173), .IN3(n28105), .IN4(n216), .IN5(
        n6985), .Q(n6982) );
  OA22X1 U6946 ( .IN1(n28113), .IN2(n259), .IN3(n28121), .IN4(n302), .Q(n6985)
         );
  OA221X1 U6947 ( .IN1(n28065), .IN2(n345), .IN3(n28073), .IN4(n388), .IN5(
        n6986), .Q(n6981) );
  OA22X1 U6948 ( .IN1(n28081), .IN2(n431), .IN3(n28089), .IN4(n474), .Q(n6986)
         );
  OA221X1 U6949 ( .IN1(n28033), .IN2(n517), .IN3(n28041), .IN4(n560), .IN5(
        n6987), .Q(n6980) );
  OA22X1 U6950 ( .IN1(n28049), .IN2(n603), .IN3(n28057), .IN4(n646), .Q(n6987)
         );
  AND3X1 U6951 ( .IN1(n6988), .IN2(n6947), .IN3(n6946), .Q(n2253) );
  NAND4X0 U6952 ( .IN1(n6989), .IN2(n6990), .IN3(n6991), .IN4(n6992), .QN(
        n6978) );
  OA221X1 U6953 ( .IN1(n28001), .IN2(n1), .IN3(n28009), .IN4(n44), .IN5(n6993), 
        .Q(n6992) );
  OA22X1 U6954 ( .IN1(n28017), .IN2(n87), .IN3(n28025), .IN4(n130), .Q(n6993)
         );
  OA221X1 U6955 ( .IN1(n27969), .IN2(n173), .IN3(n27977), .IN4(n216), .IN5(
        n6994), .Q(n6991) );
  OA22X1 U6956 ( .IN1(n27985), .IN2(n259), .IN3(n27993), .IN4(n302), .Q(n6994)
         );
  OA221X1 U6957 ( .IN1(n27937), .IN2(n345), .IN3(n27945), .IN4(n388), .IN5(
        n6995), .Q(n6990) );
  OA22X1 U6958 ( .IN1(n27953), .IN2(n431), .IN3(n27961), .IN4(n474), .Q(n6995)
         );
  OA221X1 U6959 ( .IN1(n27905), .IN2(n517), .IN3(n27913), .IN4(n560), .IN5(
        n6996), .Q(n6989) );
  OA22X1 U6960 ( .IN1(n27921), .IN2(n603), .IN3(n27929), .IN4(n646), .Q(n6996)
         );
  AND3X1 U6961 ( .IN1(n6988), .IN2(n6947), .IN3(n6957), .Q(n2251) );
  NAND4X0 U6962 ( .IN1(n6997), .IN2(n6998), .IN3(n6999), .IN4(n7000), .QN(
        n6976) );
  OA221X1 U6963 ( .IN1(n27873), .IN2(n1), .IN3(n27881), .IN4(n44), .IN5(n7001), 
        .Q(n7000) );
  OA22X1 U6964 ( .IN1(n27889), .IN2(n87), .IN3(n27897), .IN4(n130), .Q(n7001)
         );
  OA221X1 U6965 ( .IN1(n27841), .IN2(n173), .IN3(n27849), .IN4(n216), .IN5(
        n7002), .Q(n6999) );
  OA22X1 U6966 ( .IN1(n27857), .IN2(n259), .IN3(n27865), .IN4(n302), .Q(n7002)
         );
  OA221X1 U6967 ( .IN1(n27809), .IN2(n345), .IN3(n27817), .IN4(n388), .IN5(
        n7003), .Q(n6998) );
  OA22X1 U6968 ( .IN1(n27825), .IN2(n431), .IN3(n27833), .IN4(n474), .Q(n7003)
         );
  OA221X1 U6969 ( .IN1(n27777), .IN2(n517), .IN3(n27785), .IN4(n560), .IN5(
        n7004), .Q(n6997) );
  OA22X1 U6970 ( .IN1(n27793), .IN2(n603), .IN3(n27801), .IN4(n646), .Q(n7004)
         );
  AND3X1 U6971 ( .IN1(n6946), .IN2(n6947), .IN3(n7005), .Q(n2248) );
  NOR2X0 U6972 ( .IN1(N58), .IN2(n31745), .QN(n6946) );
  NAND4X0 U6973 ( .IN1(n7006), .IN2(n7007), .IN3(n7008), .IN4(n7009), .QN(
        n6975) );
  OA221X1 U6974 ( .IN1(n27745), .IN2(n1), .IN3(n27753), .IN4(n44), .IN5(n7010), 
        .Q(n7009) );
  OA22X1 U6975 ( .IN1(n27761), .IN2(n87), .IN3(n27769), .IN4(n130), .Q(n7010)
         );
  OA221X1 U6976 ( .IN1(n27713), .IN2(n173), .IN3(n27721), .IN4(n216), .IN5(
        n7011), .Q(n7008) );
  OA22X1 U6977 ( .IN1(n27729), .IN2(n259), .IN3(n27737), .IN4(n302), .Q(n7011)
         );
  OA221X1 U6978 ( .IN1(n27681), .IN2(n345), .IN3(n27689), .IN4(n388), .IN5(
        n7012), .Q(n7007) );
  OA22X1 U6979 ( .IN1(n27697), .IN2(n431), .IN3(n27705), .IN4(n474), .Q(n7012)
         );
  OA221X1 U6980 ( .IN1(n27649), .IN2(n517), .IN3(n27657), .IN4(n560), .IN5(
        n7013), .Q(n7006) );
  OA22X1 U6981 ( .IN1(n27665), .IN2(n603), .IN3(n27673), .IN4(n646), .Q(n7013)
         );
  AND3X1 U6982 ( .IN1(n6957), .IN2(n6947), .IN3(n7005), .Q(n2246) );
  NOR2X0 U6983 ( .IN1(n31745), .IN2(n31748), .QN(n6957) );
  AO221X1 U6984 ( .IN1(n2287), .IN2(n7014), .IN3(n2289), .IN4(n7015), .IN5(
        n7016), .Q(n6930) );
  AO22X1 U6985 ( .IN1(n2292), .IN2(n7017), .IN3(n2294), .IN4(n7018), .Q(n7016)
         );
  NAND4X0 U6986 ( .IN1(n7019), .IN2(n7020), .IN3(n7021), .IN4(n7022), .QN(
        n7018) );
  OA221X1 U6987 ( .IN1(n29665), .IN2(n1), .IN3(n29673), .IN4(n44), .IN5(n7023), 
        .Q(n7022) );
  OA22X1 U6988 ( .IN1(n29681), .IN2(n87), .IN3(n29689), .IN4(n130), .Q(n7023)
         );
  OA221X1 U6989 ( .IN1(n29633), .IN2(n173), .IN3(n29641), .IN4(n216), .IN5(
        n7024), .Q(n7021) );
  OA22X1 U6990 ( .IN1(n29649), .IN2(n259), .IN3(n29657), .IN4(n302), .Q(n7024)
         );
  OA221X1 U6991 ( .IN1(n29601), .IN2(n345), .IN3(n29609), .IN4(n388), .IN5(
        n7025), .Q(n7020) );
  OA22X1 U6992 ( .IN1(n29617), .IN2(n431), .IN3(n29625), .IN4(n474), .Q(n7025)
         );
  OA221X1 U6993 ( .IN1(n29569), .IN2(n517), .IN3(n29577), .IN4(n560), .IN5(
        n7026), .Q(n7019) );
  OA22X1 U6994 ( .IN1(n29585), .IN2(n603), .IN3(n29593), .IN4(n646), .Q(n7026)
         );
  AND3X1 U6995 ( .IN1(n6948), .IN2(n6947), .IN3(n7027), .Q(n2294) );
  NAND4X0 U6996 ( .IN1(n7028), .IN2(n7029), .IN3(n7030), .IN4(n7031), .QN(
        n7017) );
  OA221X1 U6997 ( .IN1(n29537), .IN2(n1), .IN3(n29545), .IN4(n44), .IN5(n7032), 
        .Q(n7031) );
  OA22X1 U6998 ( .IN1(n29553), .IN2(n87), .IN3(n29561), .IN4(n130), .Q(n7032)
         );
  OA221X1 U6999 ( .IN1(n29505), .IN2(n173), .IN3(n29513), .IN4(n216), .IN5(
        n7033), .Q(n7030) );
  OA22X1 U7000 ( .IN1(n29521), .IN2(n259), .IN3(n29529), .IN4(n302), .Q(n7033)
         );
  OA221X1 U7001 ( .IN1(n29473), .IN2(n345), .IN3(n29481), .IN4(n388), .IN5(
        n7034), .Q(n7029) );
  OA22X1 U7002 ( .IN1(n29489), .IN2(n431), .IN3(n29497), .IN4(n474), .Q(n7034)
         );
  OA221X1 U7003 ( .IN1(n29441), .IN2(n517), .IN3(n29449), .IN4(n560), .IN5(
        n7035), .Q(n7028) );
  OA22X1 U7004 ( .IN1(n29457), .IN2(n603), .IN3(n29465), .IN4(n646), .Q(n7035)
         );
  AND3X1 U7005 ( .IN1(n6948), .IN2(n6947), .IN3(n7036), .Q(n2292) );
  NOR2X0 U7006 ( .IN1(N60), .IN2(N59), .QN(n6948) );
  NAND4X0 U7007 ( .IN1(n7037), .IN2(n7038), .IN3(n7039), .IN4(n7040), .QN(
        n7015) );
  OA221X1 U7008 ( .IN1(n29409), .IN2(n1), .IN3(n29417), .IN4(n44), .IN5(n7041), 
        .Q(n7040) );
  OA22X1 U7009 ( .IN1(n29425), .IN2(n87), .IN3(n29433), .IN4(n130), .Q(n7041)
         );
  OA221X1 U7010 ( .IN1(n29377), .IN2(n173), .IN3(n29385), .IN4(n216), .IN5(
        n7042), .Q(n7039) );
  OA22X1 U7011 ( .IN1(n29393), .IN2(n259), .IN3(n29401), .IN4(n302), .Q(n7042)
         );
  OA221X1 U7012 ( .IN1(n29345), .IN2(n345), .IN3(n29353), .IN4(n388), .IN5(
        n7043), .Q(n7038) );
  OA22X1 U7013 ( .IN1(n29361), .IN2(n431), .IN3(n29369), .IN4(n474), .Q(n7043)
         );
  OA221X1 U7014 ( .IN1(n29313), .IN2(n517), .IN3(n29321), .IN4(n560), .IN5(
        n7044), .Q(n7037) );
  OA22X1 U7015 ( .IN1(n29329), .IN2(n603), .IN3(n29337), .IN4(n646), .Q(n7044)
         );
  AND2X1 U7016 ( .IN1(n7027), .IN2(n6966), .Q(n2289) );
  NAND4X0 U7017 ( .IN1(n7045), .IN2(n7046), .IN3(n7047), .IN4(n7048), .QN(
        n7014) );
  OA221X1 U7018 ( .IN1(n29281), .IN2(n1), .IN3(n29289), .IN4(n44), .IN5(n7049), 
        .Q(n7048) );
  OA22X1 U7019 ( .IN1(n29297), .IN2(n87), .IN3(n29305), .IN4(n130), .Q(n7049)
         );
  OA221X1 U7020 ( .IN1(n29249), .IN2(n173), .IN3(n29257), .IN4(n216), .IN5(
        n7050), .Q(n7047) );
  OA22X1 U7021 ( .IN1(n29265), .IN2(n259), .IN3(n29273), .IN4(n302), .Q(n7050)
         );
  OA221X1 U7022 ( .IN1(n29217), .IN2(n345), .IN3(n29225), .IN4(n388), .IN5(
        n7051), .Q(n7046) );
  OA22X1 U7023 ( .IN1(n29233), .IN2(n431), .IN3(n29241), .IN4(n474), .Q(n7051)
         );
  OA221X1 U7024 ( .IN1(n29185), .IN2(n517), .IN3(n29193), .IN4(n560), .IN5(
        n7052), .Q(n7045) );
  OA22X1 U7025 ( .IN1(n29201), .IN2(n603), .IN3(n29209), .IN4(n646), .Q(n7052)
         );
  AND2X1 U7026 ( .IN1(n7036), .IN2(n6966), .Q(n2287) );
  AND3X1 U7027 ( .IN1(N59), .IN2(n6947), .IN3(n31746), .Q(n6966) );
  AO221X1 U7028 ( .IN1(n2328), .IN2(n7053), .IN3(n2330), .IN4(n7054), .IN5(
        n7055), .Q(n6929) );
  AO22X1 U7029 ( .IN1(n2333), .IN2(n7056), .IN3(n2335), .IN4(n7057), .Q(n7055)
         );
  NAND4X0 U7030 ( .IN1(n7058), .IN2(n7059), .IN3(n7060), .IN4(n7061), .QN(
        n7057) );
  OA221X1 U7031 ( .IN1(n29153), .IN2(n1), .IN3(n29161), .IN4(n44), .IN5(n7062), 
        .Q(n7061) );
  OA22X1 U7032 ( .IN1(n29169), .IN2(n87), .IN3(n29177), .IN4(n130), .Q(n7062)
         );
  OA221X1 U7033 ( .IN1(n29121), .IN2(n173), .IN3(n29129), .IN4(n216), .IN5(
        n7063), .Q(n7060) );
  OA22X1 U7034 ( .IN1(n29137), .IN2(n259), .IN3(n29145), .IN4(n302), .Q(n7063)
         );
  OA221X1 U7035 ( .IN1(n29089), .IN2(n345), .IN3(n29097), .IN4(n388), .IN5(
        n7064), .Q(n7059) );
  OA22X1 U7036 ( .IN1(n29105), .IN2(n431), .IN3(n29113), .IN4(n474), .Q(n7064)
         );
  OA221X1 U7037 ( .IN1(n29057), .IN2(n517), .IN3(n29065), .IN4(n560), .IN5(
        n7065), .Q(n7058) );
  OA22X1 U7038 ( .IN1(n29073), .IN2(n603), .IN3(n29081), .IN4(n646), .Q(n7065)
         );
  AND3X1 U7039 ( .IN1(n6988), .IN2(n6947), .IN3(n7027), .Q(n2335) );
  NAND4X0 U7040 ( .IN1(n7066), .IN2(n7067), .IN3(n7068), .IN4(n7069), .QN(
        n7056) );
  OA221X1 U7041 ( .IN1(n29025), .IN2(n1), .IN3(n29033), .IN4(n44), .IN5(n7070), 
        .Q(n7069) );
  OA22X1 U7042 ( .IN1(n29041), .IN2(n87), .IN3(n29049), .IN4(n130), .Q(n7070)
         );
  OA221X1 U7043 ( .IN1(n28993), .IN2(n173), .IN3(n29001), .IN4(n216), .IN5(
        n7071), .Q(n7068) );
  OA22X1 U7044 ( .IN1(n29009), .IN2(n259), .IN3(n29017), .IN4(n302), .Q(n7071)
         );
  OA221X1 U7045 ( .IN1(n28961), .IN2(n345), .IN3(n28969), .IN4(n388), .IN5(
        n7072), .Q(n7067) );
  OA22X1 U7046 ( .IN1(n28977), .IN2(n431), .IN3(n28985), .IN4(n474), .Q(n7072)
         );
  OA221X1 U7047 ( .IN1(n28929), .IN2(n517), .IN3(n28937), .IN4(n560), .IN5(
        n7073), .Q(n7066) );
  OA22X1 U7048 ( .IN1(n28945), .IN2(n603), .IN3(n28953), .IN4(n646), .Q(n7073)
         );
  AND3X1 U7049 ( .IN1(n6988), .IN2(n6947), .IN3(n7036), .Q(n2333) );
  NOR2X0 U7050 ( .IN1(N59), .IN2(n31746), .QN(n6988) );
  NAND4X0 U7051 ( .IN1(n7074), .IN2(n7075), .IN3(n7076), .IN4(n7077), .QN(
        n7054) );
  OA221X1 U7052 ( .IN1(n28897), .IN2(n1), .IN3(n28905), .IN4(n44), .IN5(n7078), 
        .Q(n7077) );
  OA22X1 U7053 ( .IN1(n28913), .IN2(n87), .IN3(n28921), .IN4(n130), .Q(n7078)
         );
  OA221X1 U7054 ( .IN1(n28865), .IN2(n173), .IN3(n28873), .IN4(n216), .IN5(
        n7079), .Q(n7076) );
  OA22X1 U7055 ( .IN1(n28881), .IN2(n259), .IN3(n28889), .IN4(n302), .Q(n7079)
         );
  OA221X1 U7056 ( .IN1(n28833), .IN2(n345), .IN3(n28841), .IN4(n388), .IN5(
        n7080), .Q(n7075) );
  OA22X1 U7057 ( .IN1(n28849), .IN2(n431), .IN3(n28857), .IN4(n474), .Q(n7080)
         );
  OA221X1 U7058 ( .IN1(n28801), .IN2(n517), .IN3(n28809), .IN4(n560), .IN5(
        n7081), .Q(n7074) );
  OA22X1 U7059 ( .IN1(n28817), .IN2(n603), .IN3(n28825), .IN4(n646), .Q(n7081)
         );
  AND3X1 U7060 ( .IN1(n7005), .IN2(n6947), .IN3(n7027), .Q(n2330) );
  NOR2X0 U7061 ( .IN1(N61), .IN2(N58), .QN(n7027) );
  NAND4X0 U7062 ( .IN1(n7082), .IN2(n7083), .IN3(n7084), .IN4(n7085), .QN(
        n7053) );
  OA221X1 U7063 ( .IN1(n28769), .IN2(n1), .IN3(n28777), .IN4(n44), .IN5(n7086), 
        .Q(n7085) );
  OA22X1 U7064 ( .IN1(n28785), .IN2(n87), .IN3(n28793), .IN4(n130), .Q(n7086)
         );
  NAND2X0 U7065 ( .IN1(n7087), .IN2(n7088), .QN(n2206) );
  NAND2X0 U7066 ( .IN1(n7088), .IN2(n7089), .QN(n2205) );
  NAND2X0 U7067 ( .IN1(n7090), .IN2(n7087), .QN(n2194) );
  NAND2X0 U7068 ( .IN1(n7090), .IN2(n7089), .QN(n2170) );
  OA221X1 U7069 ( .IN1(n28737), .IN2(n173), .IN3(n28745), .IN4(n216), .IN5(
        n7091), .Q(n7084) );
  OA22X1 U7070 ( .IN1(n28753), .IN2(n259), .IN3(n28761), .IN4(n302), .Q(n7091)
         );
  NAND2X0 U7071 ( .IN1(n7092), .IN2(n7087), .QN(n2211) );
  NAND2X0 U7072 ( .IN1(n7092), .IN2(n7089), .QN(n2210) );
  NAND2X0 U7073 ( .IN1(n7093), .IN2(n7087), .QN(n2208) );
  NOR2X0 U7074 ( .IN1(N54), .IN2(N57), .QN(n7087) );
  NAND2X0 U7075 ( .IN1(n7093), .IN2(n7089), .QN(n2207) );
  NOR2X0 U7076 ( .IN1(N57), .IN2(n31750), .QN(n7089) );
  OA221X1 U7077 ( .IN1(n28705), .IN2(n345), .IN3(n28713), .IN4(n388), .IN5(
        n7094), .Q(n7083) );
  OA22X1 U7078 ( .IN1(n28721), .IN2(n431), .IN3(n28729), .IN4(n474), .Q(n7094)
         );
  NAND2X0 U7079 ( .IN1(n7095), .IN2(n7088), .QN(n2216) );
  NAND2X0 U7080 ( .IN1(n7096), .IN2(n7088), .QN(n2215) );
  NOR2X0 U7081 ( .IN1(N55), .IN2(N56), .QN(n7088) );
  NAND2X0 U7082 ( .IN1(n7095), .IN2(n7090), .QN(n2213) );
  NAND2X0 U7083 ( .IN1(n7096), .IN2(n7090), .QN(n2212) );
  NOR2X0 U7084 ( .IN1(N56), .IN2(n21497), .QN(n7090) );
  OA221X1 U7085 ( .IN1(n28673), .IN2(n517), .IN3(n28681), .IN4(n560), .IN5(
        n7097), .Q(n7082) );
  OA22X1 U7086 ( .IN1(n28689), .IN2(n603), .IN3(n28697), .IN4(n646), .Q(n7097)
         );
  NAND2X0 U7087 ( .IN1(n7095), .IN2(n7092), .QN(n2221) );
  NAND2X0 U7088 ( .IN1(n7096), .IN2(n7092), .QN(n2220) );
  NOR2X0 U7089 ( .IN1(N55), .IN2(n21496), .QN(n7092) );
  NAND2X0 U7090 ( .IN1(n7095), .IN2(n7093), .QN(n2218) );
  NOR2X0 U7091 ( .IN1(N54), .IN2(n31749), .QN(n7095) );
  NAND2X0 U7092 ( .IN1(n7096), .IN2(n7093), .QN(n2217) );
  NOR2X0 U7093 ( .IN1(n21497), .IN2(n21496), .QN(n7093) );
  NOR2X0 U7094 ( .IN1(n31750), .IN2(n31749), .QN(n7096) );
  AND3X1 U7095 ( .IN1(n7005), .IN2(n6947), .IN3(n7036), .Q(n2328) );
  NOR2X0 U7096 ( .IN1(N61), .IN2(n31748), .QN(n7036) );
  INVX0 U7097 ( .INP(rst), .ZN(n6947) );
  NOR2X0 U7098 ( .IN1(n31746), .IN2(n31747), .QN(n7005) );
  AO21X1 U7099 ( .IN1(oe), .IN2(ce), .IN3(test_se), .Q(n21510) );
  MUX21X1 U7100 ( .IN1(\mem0[255][7] ), .IN2(n843), .S(n7098), .Q(n18603) );
  MUX21X1 U7101 ( .IN1(\mem0[255][6] ), .IN2(n821), .S(n7098), .Q(n18602) );
  MUX21X1 U7102 ( .IN1(\mem0[255][5] ), .IN2(n799), .S(n7098), .Q(n18601) );
  MUX21X1 U7103 ( .IN1(\mem0[255][4] ), .IN2(n777), .S(n7098), .Q(n18600) );
  MUX21X1 U7104 ( .IN1(\mem0[255][3] ), .IN2(n755), .S(n7098), .Q(n18599) );
  MUX21X1 U7105 ( .IN1(\mem0[255][2] ), .IN2(n733), .S(n7098), .Q(n18598) );
  MUX21X1 U7106 ( .IN1(\mem0[255][1] ), .IN2(n711), .S(n7098), .Q(n18597) );
  MUX21X1 U7107 ( .IN1(\mem0[255][0] ), .IN2(n689), .S(n7098), .Q(n18596) );
  AND2X1 U7108 ( .IN1(n7099), .IN2(n7100), .Q(n7098) );
  MUX21X1 U7109 ( .IN1(\mem0[254][7] ), .IN2(n843), .S(n7101), .Q(n18595) );
  MUX21X1 U7110 ( .IN1(\mem0[254][6] ), .IN2(n821), .S(n7101), .Q(n18594) );
  MUX21X1 U7111 ( .IN1(\mem0[254][5] ), .IN2(n799), .S(n7101), .Q(n18593) );
  MUX21X1 U7112 ( .IN1(\mem0[254][4] ), .IN2(n777), .S(n7101), .Q(n18592) );
  MUX21X1 U7113 ( .IN1(\mem0[254][3] ), .IN2(n755), .S(n7101), .Q(n18591) );
  MUX21X1 U7114 ( .IN1(\mem0[254][2] ), .IN2(n733), .S(n7101), .Q(n18590) );
  MUX21X1 U7115 ( .IN1(\mem0[254][1] ), .IN2(n711), .S(n7101), .Q(n18589) );
  MUX21X1 U7116 ( .IN1(\mem0[254][0] ), .IN2(n689), .S(n7101), .Q(n18588) );
  AND2X1 U7117 ( .IN1(n7102), .IN2(n7100), .Q(n7101) );
  MUX21X1 U7118 ( .IN1(\mem0[253][7] ), .IN2(n843), .S(n7103), .Q(n18587) );
  MUX21X1 U7119 ( .IN1(\mem0[253][6] ), .IN2(n821), .S(n7103), .Q(n18586) );
  MUX21X1 U7120 ( .IN1(\mem0[253][5] ), .IN2(n799), .S(n7103), .Q(n18585) );
  MUX21X1 U7121 ( .IN1(\mem0[253][4] ), .IN2(n777), .S(n7103), .Q(n18584) );
  MUX21X1 U7122 ( .IN1(\mem0[253][3] ), .IN2(n755), .S(n7103), .Q(n18583) );
  MUX21X1 U7123 ( .IN1(\mem0[253][2] ), .IN2(n733), .S(n7103), .Q(n18582) );
  MUX21X1 U7124 ( .IN1(\mem0[253][1] ), .IN2(n711), .S(n7103), .Q(n18581) );
  MUX21X1 U7125 ( .IN1(\mem0[253][0] ), .IN2(n689), .S(n7103), .Q(n18580) );
  AND2X1 U7126 ( .IN1(n7104), .IN2(n7100), .Q(n7103) );
  MUX21X1 U7127 ( .IN1(\mem0[252][7] ), .IN2(n843), .S(n7105), .Q(n18579) );
  MUX21X1 U7128 ( .IN1(\mem0[252][6] ), .IN2(n821), .S(n7105), .Q(n18578) );
  MUX21X1 U7129 ( .IN1(\mem0[252][5] ), .IN2(n799), .S(n7105), .Q(n18577) );
  MUX21X1 U7130 ( .IN1(\mem0[252][4] ), .IN2(n777), .S(n7105), .Q(n18576) );
  MUX21X1 U7131 ( .IN1(\mem0[252][3] ), .IN2(n755), .S(n7105), .Q(n18575) );
  MUX21X1 U7132 ( .IN1(\mem0[252][2] ), .IN2(n733), .S(n7105), .Q(n18574) );
  MUX21X1 U7133 ( .IN1(\mem0[252][1] ), .IN2(n711), .S(n7105), .Q(n18573) );
  MUX21X1 U7134 ( .IN1(\mem0[252][0] ), .IN2(n689), .S(n7105), .Q(n18572) );
  AND2X1 U7135 ( .IN1(n7106), .IN2(n7100), .Q(n7105) );
  MUX21X1 U7136 ( .IN1(\mem0[251][7] ), .IN2(n843), .S(n7107), .Q(n18571) );
  MUX21X1 U7137 ( .IN1(\mem0[251][6] ), .IN2(n821), .S(n7107), .Q(n18570) );
  MUX21X1 U7138 ( .IN1(\mem0[251][5] ), .IN2(n799), .S(n7107), .Q(n18569) );
  MUX21X1 U7139 ( .IN1(\mem0[251][4] ), .IN2(n777), .S(n7107), .Q(n18568) );
  MUX21X1 U7140 ( .IN1(\mem0[251][3] ), .IN2(n755), .S(n7107), .Q(n18567) );
  MUX21X1 U7141 ( .IN1(\mem0[251][2] ), .IN2(n733), .S(n7107), .Q(n18566) );
  MUX21X1 U7142 ( .IN1(\mem0[251][1] ), .IN2(n711), .S(n7107), .Q(n18565) );
  MUX21X1 U7143 ( .IN1(\mem0[251][0] ), .IN2(n689), .S(n7107), .Q(n18564) );
  AND2X1 U7144 ( .IN1(n7108), .IN2(n7100), .Q(n7107) );
  MUX21X1 U7145 ( .IN1(\mem0[250][7] ), .IN2(n843), .S(n7109), .Q(n18563) );
  MUX21X1 U7146 ( .IN1(\mem0[250][6] ), .IN2(n821), .S(n7109), .Q(n18562) );
  MUX21X1 U7147 ( .IN1(\mem0[250][5] ), .IN2(n799), .S(n7109), .Q(n18561) );
  MUX21X1 U7148 ( .IN1(\mem0[250][4] ), .IN2(n777), .S(n7109), .Q(n18560) );
  MUX21X1 U7149 ( .IN1(\mem0[250][3] ), .IN2(n755), .S(n7109), .Q(n18559) );
  MUX21X1 U7150 ( .IN1(\mem0[250][2] ), .IN2(n733), .S(n7109), .Q(n18558) );
  MUX21X1 U7151 ( .IN1(\mem0[250][1] ), .IN2(n711), .S(n7109), .Q(n18557) );
  MUX21X1 U7152 ( .IN1(\mem0[250][0] ), .IN2(n689), .S(n7109), .Q(n18556) );
  AND2X1 U7153 ( .IN1(n7110), .IN2(n7100), .Q(n7109) );
  MUX21X1 U7154 ( .IN1(\mem0[249][7] ), .IN2(n843), .S(n7111), .Q(n18555) );
  MUX21X1 U7155 ( .IN1(\mem0[249][6] ), .IN2(n821), .S(n7111), .Q(n18554) );
  MUX21X1 U7156 ( .IN1(\mem0[249][5] ), .IN2(n799), .S(n7111), .Q(n18553) );
  MUX21X1 U7157 ( .IN1(\mem0[249][4] ), .IN2(n777), .S(n7111), .Q(n18552) );
  MUX21X1 U7158 ( .IN1(\mem0[249][3] ), .IN2(n755), .S(n7111), .Q(n18551) );
  MUX21X1 U7159 ( .IN1(\mem0[249][2] ), .IN2(n733), .S(n7111), .Q(n18550) );
  MUX21X1 U7160 ( .IN1(\mem0[249][1] ), .IN2(n711), .S(n7111), .Q(n18549) );
  MUX21X1 U7161 ( .IN1(\mem0[249][0] ), .IN2(n689), .S(n7111), .Q(n18548) );
  AND2X1 U7162 ( .IN1(n7112), .IN2(n7100), .Q(n7111) );
  MUX21X1 U7163 ( .IN1(\mem0[248][7] ), .IN2(n843), .S(n7113), .Q(n18547) );
  MUX21X1 U7164 ( .IN1(\mem0[248][6] ), .IN2(n821), .S(n7113), .Q(n18546) );
  MUX21X1 U7165 ( .IN1(\mem0[248][5] ), .IN2(n799), .S(n7113), .Q(n18545) );
  MUX21X1 U7166 ( .IN1(\mem0[248][4] ), .IN2(n777), .S(n7113), .Q(n18544) );
  MUX21X1 U7167 ( .IN1(\mem0[248][3] ), .IN2(n755), .S(n7113), .Q(n18543) );
  MUX21X1 U7168 ( .IN1(\mem0[248][2] ), .IN2(n733), .S(n7113), .Q(n18542) );
  MUX21X1 U7169 ( .IN1(\mem0[248][1] ), .IN2(n711), .S(n7113), .Q(n18541) );
  MUX21X1 U7170 ( .IN1(\mem0[248][0] ), .IN2(n689), .S(n7113), .Q(n18540) );
  AND2X1 U7171 ( .IN1(n7114), .IN2(n7100), .Q(n7113) );
  MUX21X1 U7172 ( .IN1(\mem0[247][7] ), .IN2(n843), .S(n7115), .Q(n18539) );
  MUX21X1 U7173 ( .IN1(\mem0[247][6] ), .IN2(n821), .S(n7115), .Q(n18538) );
  MUX21X1 U7174 ( .IN1(\mem0[247][5] ), .IN2(n799), .S(n7115), .Q(n18537) );
  MUX21X1 U7175 ( .IN1(\mem0[247][4] ), .IN2(n777), .S(n7115), .Q(n18536) );
  MUX21X1 U7176 ( .IN1(\mem0[247][3] ), .IN2(n755), .S(n7115), .Q(n18535) );
  MUX21X1 U7177 ( .IN1(\mem0[247][2] ), .IN2(n733), .S(n7115), .Q(n18534) );
  MUX21X1 U7178 ( .IN1(\mem0[247][1] ), .IN2(n711), .S(n7115), .Q(n18533) );
  MUX21X1 U7179 ( .IN1(\mem0[247][0] ), .IN2(n689), .S(n7115), .Q(n18532) );
  AND2X1 U7180 ( .IN1(n7116), .IN2(n7100), .Q(n7115) );
  MUX21X1 U7181 ( .IN1(\mem0[246][7] ), .IN2(n843), .S(n7117), .Q(n18531) );
  MUX21X1 U7182 ( .IN1(\mem0[246][6] ), .IN2(n821), .S(n7117), .Q(n18530) );
  MUX21X1 U7183 ( .IN1(\mem0[246][5] ), .IN2(n799), .S(n7117), .Q(n18529) );
  MUX21X1 U7184 ( .IN1(\mem0[246][4] ), .IN2(n777), .S(n7117), .Q(n18528) );
  MUX21X1 U7185 ( .IN1(\mem0[246][3] ), .IN2(n755), .S(n7117), .Q(n18527) );
  MUX21X1 U7186 ( .IN1(\mem0[246][2] ), .IN2(n733), .S(n7117), .Q(n18526) );
  MUX21X1 U7187 ( .IN1(\mem0[246][1] ), .IN2(n711), .S(n7117), .Q(n18525) );
  MUX21X1 U7188 ( .IN1(\mem0[246][0] ), .IN2(n689), .S(n7117), .Q(n18524) );
  AND2X1 U7189 ( .IN1(n7118), .IN2(n7100), .Q(n7117) );
  MUX21X1 U7190 ( .IN1(\mem0[245][7] ), .IN2(n843), .S(n7119), .Q(n18523) );
  MUX21X1 U7191 ( .IN1(\mem0[245][6] ), .IN2(n821), .S(n7119), .Q(n18522) );
  MUX21X1 U7192 ( .IN1(\mem0[245][5] ), .IN2(n799), .S(n7119), .Q(n18521) );
  MUX21X1 U7193 ( .IN1(\mem0[245][4] ), .IN2(n777), .S(n7119), .Q(n18520) );
  MUX21X1 U7194 ( .IN1(\mem0[245][3] ), .IN2(n755), .S(n7119), .Q(n18519) );
  MUX21X1 U7195 ( .IN1(\mem0[245][2] ), .IN2(n733), .S(n7119), .Q(n18518) );
  MUX21X1 U7196 ( .IN1(\mem0[245][1] ), .IN2(n711), .S(n7119), .Q(n18517) );
  MUX21X1 U7197 ( .IN1(\mem0[245][0] ), .IN2(n689), .S(n7119), .Q(n18516) );
  AND2X1 U7198 ( .IN1(n7120), .IN2(n7100), .Q(n7119) );
  MUX21X1 U7199 ( .IN1(\mem0[244][7] ), .IN2(n843), .S(n7121), .Q(n18515) );
  MUX21X1 U7200 ( .IN1(\mem0[244][6] ), .IN2(n821), .S(n7121), .Q(n18514) );
  MUX21X1 U7201 ( .IN1(\mem0[244][5] ), .IN2(n799), .S(n7121), .Q(n18513) );
  MUX21X1 U7202 ( .IN1(\mem0[244][4] ), .IN2(n777), .S(n7121), .Q(n18512) );
  MUX21X1 U7203 ( .IN1(\mem0[244][3] ), .IN2(n755), .S(n7121), .Q(n18511) );
  MUX21X1 U7204 ( .IN1(\mem0[244][2] ), .IN2(n733), .S(n7121), .Q(n18510) );
  MUX21X1 U7205 ( .IN1(\mem0[244][1] ), .IN2(n711), .S(n7121), .Q(n18509) );
  MUX21X1 U7206 ( .IN1(\mem0[244][0] ), .IN2(n689), .S(n7121), .Q(n18508) );
  AND2X1 U7207 ( .IN1(n7122), .IN2(n7100), .Q(n7121) );
  MUX21X1 U7208 ( .IN1(\mem0[243][7] ), .IN2(n844), .S(n7123), .Q(n18507) );
  MUX21X1 U7209 ( .IN1(\mem0[243][6] ), .IN2(n822), .S(n7123), .Q(n18506) );
  MUX21X1 U7210 ( .IN1(\mem0[243][5] ), .IN2(n800), .S(n7123), .Q(n18505) );
  MUX21X1 U7211 ( .IN1(\mem0[243][4] ), .IN2(n778), .S(n7123), .Q(n18504) );
  MUX21X1 U7212 ( .IN1(\mem0[243][3] ), .IN2(n756), .S(n7123), .Q(n18503) );
  MUX21X1 U7213 ( .IN1(\mem0[243][2] ), .IN2(n734), .S(n7123), .Q(n18502) );
  MUX21X1 U7214 ( .IN1(\mem0[243][1] ), .IN2(n712), .S(n7123), .Q(n18501) );
  MUX21X1 U7215 ( .IN1(\mem0[243][0] ), .IN2(n690), .S(n7123), .Q(n18500) );
  AND2X1 U7216 ( .IN1(n7124), .IN2(n7100), .Q(n7123) );
  MUX21X1 U7217 ( .IN1(\mem0[242][7] ), .IN2(n844), .S(n7125), .Q(n18499) );
  MUX21X1 U7218 ( .IN1(\mem0[242][6] ), .IN2(n822), .S(n7125), .Q(n18498) );
  MUX21X1 U7219 ( .IN1(\mem0[242][5] ), .IN2(n800), .S(n7125), .Q(n18497) );
  MUX21X1 U7220 ( .IN1(\mem0[242][4] ), .IN2(n778), .S(n7125), .Q(n18496) );
  MUX21X1 U7221 ( .IN1(\mem0[242][3] ), .IN2(n756), .S(n7125), .Q(n18495) );
  MUX21X1 U7222 ( .IN1(\mem0[242][2] ), .IN2(n734), .S(n7125), .Q(n18494) );
  MUX21X1 U7223 ( .IN1(\mem0[242][1] ), .IN2(n712), .S(n7125), .Q(n18493) );
  MUX21X1 U7224 ( .IN1(\mem0[242][0] ), .IN2(n690), .S(n7125), .Q(n18492) );
  AND2X1 U7225 ( .IN1(n7126), .IN2(n7100), .Q(n7125) );
  MUX21X1 U7226 ( .IN1(\mem0[241][7] ), .IN2(n844), .S(n7127), .Q(n18491) );
  MUX21X1 U7227 ( .IN1(\mem0[241][6] ), .IN2(n822), .S(n7127), .Q(n18490) );
  MUX21X1 U7228 ( .IN1(\mem0[241][5] ), .IN2(n800), .S(n7127), .Q(n18489) );
  MUX21X1 U7229 ( .IN1(\mem0[241][4] ), .IN2(n778), .S(n7127), .Q(n18488) );
  MUX21X1 U7230 ( .IN1(\mem0[241][3] ), .IN2(n756), .S(n7127), .Q(n18487) );
  MUX21X1 U7231 ( .IN1(\mem0[241][2] ), .IN2(n734), .S(n7127), .Q(n18486) );
  MUX21X1 U7232 ( .IN1(\mem0[241][1] ), .IN2(n712), .S(n7127), .Q(n18485) );
  MUX21X1 U7233 ( .IN1(\mem0[241][0] ), .IN2(n690), .S(n7127), .Q(n18484) );
  AND2X1 U7234 ( .IN1(n7128), .IN2(n7100), .Q(n7127) );
  MUX21X1 U7235 ( .IN1(\mem0[240][7] ), .IN2(n844), .S(n7129), .Q(n18483) );
  MUX21X1 U7236 ( .IN1(\mem0[240][6] ), .IN2(n822), .S(n7129), .Q(n18482) );
  MUX21X1 U7237 ( .IN1(\mem0[240][5] ), .IN2(n800), .S(n7129), .Q(n18481) );
  MUX21X1 U7238 ( .IN1(\mem0[240][4] ), .IN2(n778), .S(n7129), .Q(n18480) );
  MUX21X1 U7239 ( .IN1(\mem0[240][3] ), .IN2(n756), .S(n7129), .Q(n18479) );
  MUX21X1 U7240 ( .IN1(\mem0[240][2] ), .IN2(n734), .S(n7129), .Q(n18478) );
  MUX21X1 U7241 ( .IN1(\mem0[240][1] ), .IN2(n712), .S(n7129), .Q(n18477) );
  MUX21X1 U7242 ( .IN1(\mem0[240][0] ), .IN2(n690), .S(n7129), .Q(n18476) );
  AND2X1 U7243 ( .IN1(n7130), .IN2(n7100), .Q(n7129) );
  AND2X1 U7244 ( .IN1(n7131), .IN2(n7132), .Q(n7100) );
  MUX21X1 U7245 ( .IN1(\mem0[239][7] ), .IN2(n844), .S(n7133), .Q(n18475) );
  MUX21X1 U7246 ( .IN1(\mem0[239][6] ), .IN2(n822), .S(n7133), .Q(n18474) );
  MUX21X1 U7247 ( .IN1(\mem0[239][5] ), .IN2(n800), .S(n7133), .Q(n18473) );
  MUX21X1 U7248 ( .IN1(\mem0[239][4] ), .IN2(n778), .S(n7133), .Q(n18472) );
  MUX21X1 U7249 ( .IN1(\mem0[239][3] ), .IN2(n756), .S(n7133), .Q(n18471) );
  MUX21X1 U7250 ( .IN1(\mem0[239][2] ), .IN2(n734), .S(n7133), .Q(n18470) );
  MUX21X1 U7251 ( .IN1(\mem0[239][1] ), .IN2(n712), .S(n7133), .Q(n18469) );
  MUX21X1 U7252 ( .IN1(\mem0[239][0] ), .IN2(n690), .S(n7133), .Q(n18468) );
  AND2X1 U7253 ( .IN1(n7134), .IN2(n7099), .Q(n7133) );
  MUX21X1 U7254 ( .IN1(\mem0[238][7] ), .IN2(n844), .S(n7135), .Q(n18467) );
  MUX21X1 U7255 ( .IN1(\mem0[238][6] ), .IN2(n822), .S(n7135), .Q(n18466) );
  MUX21X1 U7256 ( .IN1(\mem0[238][5] ), .IN2(n800), .S(n7135), .Q(n18465) );
  MUX21X1 U7257 ( .IN1(\mem0[238][4] ), .IN2(n778), .S(n7135), .Q(n18464) );
  MUX21X1 U7258 ( .IN1(\mem0[238][3] ), .IN2(n756), .S(n7135), .Q(n18463) );
  MUX21X1 U7259 ( .IN1(\mem0[238][2] ), .IN2(n734), .S(n7135), .Q(n18462) );
  MUX21X1 U7260 ( .IN1(\mem0[238][1] ), .IN2(n712), .S(n7135), .Q(n18461) );
  MUX21X1 U7261 ( .IN1(\mem0[238][0] ), .IN2(n690), .S(n7135), .Q(n18460) );
  AND2X1 U7262 ( .IN1(n7134), .IN2(n7102), .Q(n7135) );
  MUX21X1 U7263 ( .IN1(\mem0[237][7] ), .IN2(n844), .S(n7136), .Q(n18459) );
  MUX21X1 U7264 ( .IN1(\mem0[237][6] ), .IN2(n822), .S(n7136), .Q(n18458) );
  MUX21X1 U7265 ( .IN1(\mem0[237][5] ), .IN2(n800), .S(n7136), .Q(n18457) );
  MUX21X1 U7266 ( .IN1(\mem0[237][4] ), .IN2(n778), .S(n7136), .Q(n18456) );
  MUX21X1 U7267 ( .IN1(\mem0[237][3] ), .IN2(n756), .S(n7136), .Q(n18455) );
  MUX21X1 U7268 ( .IN1(\mem0[237][2] ), .IN2(n734), .S(n7136), .Q(n18454) );
  MUX21X1 U7269 ( .IN1(\mem0[237][1] ), .IN2(n712), .S(n7136), .Q(n18453) );
  MUX21X1 U7270 ( .IN1(\mem0[237][0] ), .IN2(n690), .S(n7136), .Q(n18452) );
  AND2X1 U7271 ( .IN1(n7134), .IN2(n7104), .Q(n7136) );
  MUX21X1 U7272 ( .IN1(\mem0[236][7] ), .IN2(n844), .S(n7137), .Q(n18451) );
  MUX21X1 U7273 ( .IN1(\mem0[236][6] ), .IN2(n822), .S(n7137), .Q(n18450) );
  MUX21X1 U7274 ( .IN1(\mem0[236][5] ), .IN2(n800), .S(n7137), .Q(n18449) );
  MUX21X1 U7275 ( .IN1(\mem0[236][4] ), .IN2(n778), .S(n7137), .Q(n18448) );
  MUX21X1 U7276 ( .IN1(\mem0[236][3] ), .IN2(n756), .S(n7137), .Q(n18447) );
  MUX21X1 U7277 ( .IN1(\mem0[236][2] ), .IN2(n734), .S(n7137), .Q(n18446) );
  MUX21X1 U7278 ( .IN1(\mem0[236][1] ), .IN2(n712), .S(n7137), .Q(n18445) );
  MUX21X1 U7279 ( .IN1(\mem0[236][0] ), .IN2(n690), .S(n7137), .Q(n18444) );
  AND2X1 U7280 ( .IN1(n7134), .IN2(n7106), .Q(n7137) );
  MUX21X1 U7281 ( .IN1(\mem0[235][7] ), .IN2(n844), .S(n7138), .Q(n18443) );
  MUX21X1 U7282 ( .IN1(\mem0[235][6] ), .IN2(n822), .S(n7138), .Q(n18442) );
  MUX21X1 U7283 ( .IN1(\mem0[235][5] ), .IN2(n800), .S(n7138), .Q(n18441) );
  MUX21X1 U7284 ( .IN1(\mem0[235][4] ), .IN2(n778), .S(n7138), .Q(n18440) );
  MUX21X1 U7285 ( .IN1(\mem0[235][3] ), .IN2(n756), .S(n7138), .Q(n18439) );
  MUX21X1 U7286 ( .IN1(\mem0[235][2] ), .IN2(n734), .S(n7138), .Q(n18438) );
  MUX21X1 U7287 ( .IN1(\mem0[235][1] ), .IN2(n712), .S(n7138), .Q(n18437) );
  MUX21X1 U7288 ( .IN1(\mem0[235][0] ), .IN2(n690), .S(n7138), .Q(n18436) );
  AND2X1 U7289 ( .IN1(n7134), .IN2(n7108), .Q(n7138) );
  MUX21X1 U7290 ( .IN1(\mem0[234][7] ), .IN2(n844), .S(n7139), .Q(n18435) );
  MUX21X1 U7291 ( .IN1(\mem0[234][6] ), .IN2(n822), .S(n7139), .Q(n18434) );
  MUX21X1 U7292 ( .IN1(\mem0[234][5] ), .IN2(n800), .S(n7139), .Q(n18433) );
  MUX21X1 U7293 ( .IN1(\mem0[234][4] ), .IN2(n778), .S(n7139), .Q(n18432) );
  MUX21X1 U7294 ( .IN1(\mem0[234][3] ), .IN2(n756), .S(n7139), .Q(n18431) );
  MUX21X1 U7295 ( .IN1(\mem0[234][2] ), .IN2(n734), .S(n7139), .Q(n18430) );
  MUX21X1 U7296 ( .IN1(\mem0[234][1] ), .IN2(n712), .S(n7139), .Q(n18429) );
  MUX21X1 U7297 ( .IN1(\mem0[234][0] ), .IN2(n690), .S(n7139), .Q(n18428) );
  AND2X1 U7298 ( .IN1(n7134), .IN2(n7110), .Q(n7139) );
  MUX21X1 U7299 ( .IN1(\mem0[233][7] ), .IN2(n844), .S(n7140), .Q(n18427) );
  MUX21X1 U7300 ( .IN1(\mem0[233][6] ), .IN2(n822), .S(n7140), .Q(n18426) );
  MUX21X1 U7301 ( .IN1(\mem0[233][5] ), .IN2(n800), .S(n7140), .Q(n18425) );
  MUX21X1 U7302 ( .IN1(\mem0[233][4] ), .IN2(n778), .S(n7140), .Q(n18424) );
  MUX21X1 U7303 ( .IN1(\mem0[233][3] ), .IN2(n756), .S(n7140), .Q(n18423) );
  MUX21X1 U7304 ( .IN1(\mem0[233][2] ), .IN2(n734), .S(n7140), .Q(n18422) );
  MUX21X1 U7305 ( .IN1(\mem0[233][1] ), .IN2(n712), .S(n7140), .Q(n18421) );
  MUX21X1 U7306 ( .IN1(\mem0[233][0] ), .IN2(n690), .S(n7140), .Q(n18420) );
  AND2X1 U7307 ( .IN1(n7134), .IN2(n7112), .Q(n7140) );
  MUX21X1 U7308 ( .IN1(\mem0[232][7] ), .IN2(n844), .S(n7141), .Q(n18419) );
  MUX21X1 U7309 ( .IN1(\mem0[232][6] ), .IN2(n822), .S(n7141), .Q(n18418) );
  MUX21X1 U7310 ( .IN1(\mem0[232][5] ), .IN2(n800), .S(n7141), .Q(n18417) );
  MUX21X1 U7311 ( .IN1(\mem0[232][4] ), .IN2(n778), .S(n7141), .Q(n18416) );
  MUX21X1 U7312 ( .IN1(\mem0[232][3] ), .IN2(n756), .S(n7141), .Q(n18415) );
  MUX21X1 U7313 ( .IN1(\mem0[232][2] ), .IN2(n734), .S(n7141), .Q(n18414) );
  MUX21X1 U7314 ( .IN1(\mem0[232][1] ), .IN2(n712), .S(n7141), .Q(n18413) );
  MUX21X1 U7315 ( .IN1(\mem0[232][0] ), .IN2(n690), .S(n7141), .Q(n18412) );
  AND2X1 U7316 ( .IN1(n7134), .IN2(n7114), .Q(n7141) );
  MUX21X1 U7317 ( .IN1(\mem0[231][7] ), .IN2(n845), .S(n7142), .Q(n18411) );
  MUX21X1 U7318 ( .IN1(\mem0[231][6] ), .IN2(n823), .S(n7142), .Q(n18410) );
  MUX21X1 U7319 ( .IN1(\mem0[231][5] ), .IN2(n801), .S(n7142), .Q(n18409) );
  MUX21X1 U7320 ( .IN1(\mem0[231][4] ), .IN2(n779), .S(n7142), .Q(n18408) );
  MUX21X1 U7321 ( .IN1(\mem0[231][3] ), .IN2(n757), .S(n7142), .Q(n18407) );
  MUX21X1 U7322 ( .IN1(\mem0[231][2] ), .IN2(n735), .S(n7142), .Q(n18406) );
  MUX21X1 U7323 ( .IN1(\mem0[231][1] ), .IN2(n713), .S(n7142), .Q(n18405) );
  MUX21X1 U7324 ( .IN1(\mem0[231][0] ), .IN2(n691), .S(n7142), .Q(n18404) );
  AND2X1 U7325 ( .IN1(n7134), .IN2(n7116), .Q(n7142) );
  MUX21X1 U7326 ( .IN1(\mem0[230][7] ), .IN2(n845), .S(n7143), .Q(n18403) );
  MUX21X1 U7327 ( .IN1(\mem0[230][6] ), .IN2(n823), .S(n7143), .Q(n18402) );
  MUX21X1 U7328 ( .IN1(\mem0[230][5] ), .IN2(n801), .S(n7143), .Q(n18401) );
  MUX21X1 U7329 ( .IN1(\mem0[230][4] ), .IN2(n779), .S(n7143), .Q(n18400) );
  MUX21X1 U7330 ( .IN1(\mem0[230][3] ), .IN2(n757), .S(n7143), .Q(n18399) );
  MUX21X1 U7331 ( .IN1(\mem0[230][2] ), .IN2(n735), .S(n7143), .Q(n18398) );
  MUX21X1 U7332 ( .IN1(\mem0[230][1] ), .IN2(n713), .S(n7143), .Q(n18397) );
  MUX21X1 U7333 ( .IN1(\mem0[230][0] ), .IN2(n691), .S(n7143), .Q(n18396) );
  AND2X1 U7334 ( .IN1(n7134), .IN2(n7118), .Q(n7143) );
  MUX21X1 U7335 ( .IN1(\mem0[229][7] ), .IN2(n845), .S(n7144), .Q(n18395) );
  MUX21X1 U7336 ( .IN1(\mem0[229][6] ), .IN2(n823), .S(n7144), .Q(n18394) );
  MUX21X1 U7337 ( .IN1(\mem0[229][5] ), .IN2(n801), .S(n7144), .Q(n18393) );
  MUX21X1 U7338 ( .IN1(\mem0[229][4] ), .IN2(n779), .S(n7144), .Q(n18392) );
  MUX21X1 U7339 ( .IN1(\mem0[229][3] ), .IN2(n757), .S(n7144), .Q(n18391) );
  MUX21X1 U7340 ( .IN1(\mem0[229][2] ), .IN2(n735), .S(n7144), .Q(n18390) );
  MUX21X1 U7341 ( .IN1(\mem0[229][1] ), .IN2(n713), .S(n7144), .Q(n18389) );
  MUX21X1 U7342 ( .IN1(\mem0[229][0] ), .IN2(n691), .S(n7144), .Q(n18388) );
  AND2X1 U7343 ( .IN1(n7134), .IN2(n7120), .Q(n7144) );
  MUX21X1 U7344 ( .IN1(\mem0[228][7] ), .IN2(n845), .S(n7145), .Q(n18387) );
  MUX21X1 U7345 ( .IN1(\mem0[228][6] ), .IN2(n823), .S(n7145), .Q(n18386) );
  MUX21X1 U7346 ( .IN1(\mem0[228][5] ), .IN2(n801), .S(n7145), .Q(n18385) );
  MUX21X1 U7347 ( .IN1(\mem0[228][4] ), .IN2(n779), .S(n7145), .Q(n18384) );
  MUX21X1 U7348 ( .IN1(\mem0[228][3] ), .IN2(n757), .S(n7145), .Q(n18383) );
  MUX21X1 U7349 ( .IN1(\mem0[228][2] ), .IN2(n735), .S(n7145), .Q(n18382) );
  MUX21X1 U7350 ( .IN1(\mem0[228][1] ), .IN2(n713), .S(n7145), .Q(n18381) );
  MUX21X1 U7351 ( .IN1(\mem0[228][0] ), .IN2(n691), .S(n7145), .Q(n18380) );
  AND2X1 U7352 ( .IN1(n7134), .IN2(n7122), .Q(n7145) );
  MUX21X1 U7353 ( .IN1(\mem0[227][7] ), .IN2(n845), .S(n7146), .Q(n18379) );
  MUX21X1 U7354 ( .IN1(\mem0[227][6] ), .IN2(n823), .S(n7146), .Q(n18378) );
  MUX21X1 U7355 ( .IN1(\mem0[227][5] ), .IN2(n801), .S(n7146), .Q(n18377) );
  MUX21X1 U7356 ( .IN1(\mem0[227][4] ), .IN2(n779), .S(n7146), .Q(n18376) );
  MUX21X1 U7357 ( .IN1(\mem0[227][3] ), .IN2(n757), .S(n7146), .Q(n18375) );
  MUX21X1 U7358 ( .IN1(\mem0[227][2] ), .IN2(n735), .S(n7146), .Q(n18374) );
  MUX21X1 U7359 ( .IN1(\mem0[227][1] ), .IN2(n713), .S(n7146), .Q(n18373) );
  MUX21X1 U7360 ( .IN1(\mem0[227][0] ), .IN2(n691), .S(n7146), .Q(n18372) );
  AND2X1 U7361 ( .IN1(n7134), .IN2(n7124), .Q(n7146) );
  MUX21X1 U7362 ( .IN1(\mem0[226][7] ), .IN2(n845), .S(n7147), .Q(n18371) );
  MUX21X1 U7363 ( .IN1(\mem0[226][6] ), .IN2(n823), .S(n7147), .Q(n18370) );
  MUX21X1 U7364 ( .IN1(\mem0[226][5] ), .IN2(n801), .S(n7147), .Q(n18369) );
  MUX21X1 U7365 ( .IN1(\mem0[226][4] ), .IN2(n779), .S(n7147), .Q(n18368) );
  MUX21X1 U7366 ( .IN1(\mem0[226][3] ), .IN2(n757), .S(n7147), .Q(n18367) );
  MUX21X1 U7367 ( .IN1(\mem0[226][2] ), .IN2(n735), .S(n7147), .Q(n18366) );
  MUX21X1 U7368 ( .IN1(\mem0[226][1] ), .IN2(n713), .S(n7147), .Q(n18365) );
  MUX21X1 U7369 ( .IN1(\mem0[226][0] ), .IN2(n691), .S(n7147), .Q(n18364) );
  AND2X1 U7370 ( .IN1(n7134), .IN2(n7126), .Q(n7147) );
  MUX21X1 U7371 ( .IN1(\mem0[225][7] ), .IN2(n845), .S(n7148), .Q(n18363) );
  MUX21X1 U7372 ( .IN1(\mem0[225][6] ), .IN2(n823), .S(n7148), .Q(n18362) );
  MUX21X1 U7373 ( .IN1(\mem0[225][5] ), .IN2(n801), .S(n7148), .Q(n18361) );
  MUX21X1 U7374 ( .IN1(\mem0[225][4] ), .IN2(n779), .S(n7148), .Q(n18360) );
  MUX21X1 U7375 ( .IN1(\mem0[225][3] ), .IN2(n757), .S(n7148), .Q(n18359) );
  MUX21X1 U7376 ( .IN1(\mem0[225][2] ), .IN2(n735), .S(n7148), .Q(n18358) );
  MUX21X1 U7377 ( .IN1(\mem0[225][1] ), .IN2(n713), .S(n7148), .Q(n18357) );
  MUX21X1 U7378 ( .IN1(\mem0[225][0] ), .IN2(n691), .S(n7148), .Q(n18356) );
  AND2X1 U7379 ( .IN1(n7134), .IN2(n7128), .Q(n7148) );
  MUX21X1 U7380 ( .IN1(\mem0[224][7] ), .IN2(n845), .S(n7149), .Q(n18355) );
  MUX21X1 U7381 ( .IN1(\mem0[224][6] ), .IN2(n823), .S(n7149), .Q(n18354) );
  MUX21X1 U7382 ( .IN1(\mem0[224][5] ), .IN2(n801), .S(n7149), .Q(n18353) );
  MUX21X1 U7383 ( .IN1(\mem0[224][4] ), .IN2(n779), .S(n7149), .Q(n18352) );
  MUX21X1 U7384 ( .IN1(\mem0[224][3] ), .IN2(n757), .S(n7149), .Q(n18351) );
  MUX21X1 U7385 ( .IN1(\mem0[224][2] ), .IN2(n735), .S(n7149), .Q(n18350) );
  MUX21X1 U7386 ( .IN1(\mem0[224][1] ), .IN2(n713), .S(n7149), .Q(n18349) );
  MUX21X1 U7387 ( .IN1(\mem0[224][0] ), .IN2(n691), .S(n7149), .Q(n18348) );
  AND2X1 U7388 ( .IN1(n7134), .IN2(n7130), .Q(n7149) );
  AND2X1 U7389 ( .IN1(n7150), .IN2(n7132), .Q(n7134) );
  MUX21X1 U7390 ( .IN1(\mem0[223][7] ), .IN2(n845), .S(n7151), .Q(n18347) );
  MUX21X1 U7391 ( .IN1(\mem0[223][6] ), .IN2(n823), .S(n7151), .Q(n18346) );
  MUX21X1 U7392 ( .IN1(\mem0[223][5] ), .IN2(n801), .S(n7151), .Q(n18345) );
  MUX21X1 U7393 ( .IN1(\mem0[223][4] ), .IN2(n779), .S(n7151), .Q(n18344) );
  MUX21X1 U7394 ( .IN1(\mem0[223][3] ), .IN2(n757), .S(n7151), .Q(n18343) );
  MUX21X1 U7395 ( .IN1(\mem0[223][2] ), .IN2(n735), .S(n7151), .Q(n18342) );
  MUX21X1 U7396 ( .IN1(\mem0[223][1] ), .IN2(n713), .S(n7151), .Q(n18341) );
  MUX21X1 U7397 ( .IN1(\mem0[223][0] ), .IN2(n691), .S(n7151), .Q(n18340) );
  AND2X1 U7398 ( .IN1(n7152), .IN2(n7099), .Q(n7151) );
  MUX21X1 U7399 ( .IN1(\mem0[222][7] ), .IN2(n845), .S(n7153), .Q(n18339) );
  MUX21X1 U7400 ( .IN1(\mem0[222][6] ), .IN2(n823), .S(n7153), .Q(n18338) );
  MUX21X1 U7401 ( .IN1(\mem0[222][5] ), .IN2(n801), .S(n7153), .Q(n18337) );
  MUX21X1 U7402 ( .IN1(\mem0[222][4] ), .IN2(n779), .S(n7153), .Q(n18336) );
  MUX21X1 U7403 ( .IN1(\mem0[222][3] ), .IN2(n757), .S(n7153), .Q(n18335) );
  MUX21X1 U7404 ( .IN1(\mem0[222][2] ), .IN2(n735), .S(n7153), .Q(n18334) );
  MUX21X1 U7405 ( .IN1(\mem0[222][1] ), .IN2(n713), .S(n7153), .Q(n18333) );
  MUX21X1 U7406 ( .IN1(\mem0[222][0] ), .IN2(n691), .S(n7153), .Q(n18332) );
  AND2X1 U7407 ( .IN1(n7152), .IN2(n7102), .Q(n7153) );
  MUX21X1 U7408 ( .IN1(\mem0[221][7] ), .IN2(n845), .S(n7154), .Q(n18331) );
  MUX21X1 U7409 ( .IN1(\mem0[221][6] ), .IN2(n823), .S(n7154), .Q(n18330) );
  MUX21X1 U7410 ( .IN1(\mem0[221][5] ), .IN2(n801), .S(n7154), .Q(n18329) );
  MUX21X1 U7411 ( .IN1(\mem0[221][4] ), .IN2(n779), .S(n7154), .Q(n18328) );
  MUX21X1 U7412 ( .IN1(\mem0[221][3] ), .IN2(n757), .S(n7154), .Q(n18327) );
  MUX21X1 U7413 ( .IN1(\mem0[221][2] ), .IN2(n735), .S(n7154), .Q(n18326) );
  MUX21X1 U7414 ( .IN1(\mem0[221][1] ), .IN2(n713), .S(n7154), .Q(n18325) );
  MUX21X1 U7415 ( .IN1(\mem0[221][0] ), .IN2(n691), .S(n7154), .Q(n18324) );
  AND2X1 U7416 ( .IN1(n7152), .IN2(n7104), .Q(n7154) );
  MUX21X1 U7417 ( .IN1(\mem0[220][7] ), .IN2(n845), .S(n7155), .Q(n18323) );
  MUX21X1 U7418 ( .IN1(\mem0[220][6] ), .IN2(n823), .S(n7155), .Q(n18322) );
  MUX21X1 U7419 ( .IN1(\mem0[220][5] ), .IN2(n801), .S(n7155), .Q(n18321) );
  MUX21X1 U7420 ( .IN1(\mem0[220][4] ), .IN2(n779), .S(n7155), .Q(n18320) );
  MUX21X1 U7421 ( .IN1(\mem0[220][3] ), .IN2(n757), .S(n7155), .Q(n18319) );
  MUX21X1 U7422 ( .IN1(\mem0[220][2] ), .IN2(n735), .S(n7155), .Q(n18318) );
  MUX21X1 U7423 ( .IN1(\mem0[220][1] ), .IN2(n713), .S(n7155), .Q(n18317) );
  MUX21X1 U7424 ( .IN1(\mem0[220][0] ), .IN2(n691), .S(n7155), .Q(n18316) );
  AND2X1 U7425 ( .IN1(n7152), .IN2(n7106), .Q(n7155) );
  MUX21X1 U7426 ( .IN1(\mem0[219][7] ), .IN2(n846), .S(n7156), .Q(n18315) );
  MUX21X1 U7427 ( .IN1(\mem0[219][6] ), .IN2(n824), .S(n7156), .Q(n18314) );
  MUX21X1 U7428 ( .IN1(\mem0[219][5] ), .IN2(n802), .S(n7156), .Q(n18313) );
  MUX21X1 U7429 ( .IN1(\mem0[219][4] ), .IN2(n780), .S(n7156), .Q(n18312) );
  MUX21X1 U7430 ( .IN1(\mem0[219][3] ), .IN2(n758), .S(n7156), .Q(n18311) );
  MUX21X1 U7431 ( .IN1(\mem0[219][2] ), .IN2(n736), .S(n7156), .Q(n18310) );
  MUX21X1 U7432 ( .IN1(\mem0[219][1] ), .IN2(n714), .S(n7156), .Q(n18309) );
  MUX21X1 U7433 ( .IN1(\mem0[219][0] ), .IN2(n692), .S(n7156), .Q(n18308) );
  AND2X1 U7434 ( .IN1(n7152), .IN2(n7108), .Q(n7156) );
  MUX21X1 U7435 ( .IN1(\mem0[218][7] ), .IN2(n846), .S(n7157), .Q(n18307) );
  MUX21X1 U7436 ( .IN1(\mem0[218][6] ), .IN2(n824), .S(n7157), .Q(n18306) );
  MUX21X1 U7437 ( .IN1(\mem0[218][5] ), .IN2(n802), .S(n7157), .Q(n18305) );
  MUX21X1 U7438 ( .IN1(\mem0[218][4] ), .IN2(n780), .S(n7157), .Q(n18304) );
  MUX21X1 U7439 ( .IN1(\mem0[218][3] ), .IN2(n758), .S(n7157), .Q(n18303) );
  MUX21X1 U7440 ( .IN1(\mem0[218][2] ), .IN2(n736), .S(n7157), .Q(n18302) );
  MUX21X1 U7441 ( .IN1(\mem0[218][1] ), .IN2(n714), .S(n7157), .Q(n18301) );
  MUX21X1 U7442 ( .IN1(\mem0[218][0] ), .IN2(n692), .S(n7157), .Q(n18300) );
  AND2X1 U7443 ( .IN1(n7152), .IN2(n7110), .Q(n7157) );
  MUX21X1 U7444 ( .IN1(\mem0[217][7] ), .IN2(n846), .S(n7158), .Q(n18299) );
  MUX21X1 U7445 ( .IN1(\mem0[217][6] ), .IN2(n824), .S(n7158), .Q(n18298) );
  MUX21X1 U7446 ( .IN1(\mem0[217][5] ), .IN2(n802), .S(n7158), .Q(n18297) );
  MUX21X1 U7447 ( .IN1(\mem0[217][4] ), .IN2(n780), .S(n7158), .Q(n18296) );
  MUX21X1 U7448 ( .IN1(\mem0[217][3] ), .IN2(n758), .S(n7158), .Q(n18295) );
  MUX21X1 U7449 ( .IN1(\mem0[217][2] ), .IN2(n736), .S(n7158), .Q(n18294) );
  MUX21X1 U7450 ( .IN1(\mem0[217][1] ), .IN2(n714), .S(n7158), .Q(n18293) );
  MUX21X1 U7451 ( .IN1(\mem0[217][0] ), .IN2(n692), .S(n7158), .Q(n18292) );
  AND2X1 U7452 ( .IN1(n7152), .IN2(n7112), .Q(n7158) );
  MUX21X1 U7453 ( .IN1(\mem0[216][7] ), .IN2(n846), .S(n7159), .Q(n18291) );
  MUX21X1 U7454 ( .IN1(\mem0[216][6] ), .IN2(n824), .S(n7159), .Q(n18290) );
  MUX21X1 U7455 ( .IN1(\mem0[216][5] ), .IN2(n802), .S(n7159), .Q(n18289) );
  MUX21X1 U7456 ( .IN1(\mem0[216][4] ), .IN2(n780), .S(n7159), .Q(n18288) );
  MUX21X1 U7457 ( .IN1(\mem0[216][3] ), .IN2(n758), .S(n7159), .Q(n18287) );
  MUX21X1 U7458 ( .IN1(\mem0[216][2] ), .IN2(n736), .S(n7159), .Q(n18286) );
  MUX21X1 U7459 ( .IN1(\mem0[216][1] ), .IN2(n714), .S(n7159), .Q(n18285) );
  MUX21X1 U7460 ( .IN1(\mem0[216][0] ), .IN2(n692), .S(n7159), .Q(n18284) );
  AND2X1 U7461 ( .IN1(n7152), .IN2(n7114), .Q(n7159) );
  MUX21X1 U7462 ( .IN1(\mem0[215][7] ), .IN2(n846), .S(n7160), .Q(n18283) );
  MUX21X1 U7463 ( .IN1(\mem0[215][6] ), .IN2(n824), .S(n7160), .Q(n18282) );
  MUX21X1 U7464 ( .IN1(\mem0[215][5] ), .IN2(n802), .S(n7160), .Q(n18281) );
  MUX21X1 U7465 ( .IN1(\mem0[215][4] ), .IN2(n780), .S(n7160), .Q(n18280) );
  MUX21X1 U7466 ( .IN1(\mem0[215][3] ), .IN2(n758), .S(n7160), .Q(n18279) );
  MUX21X1 U7467 ( .IN1(\mem0[215][2] ), .IN2(n736), .S(n7160), .Q(n18278) );
  MUX21X1 U7468 ( .IN1(\mem0[215][1] ), .IN2(n714), .S(n7160), .Q(n18277) );
  MUX21X1 U7469 ( .IN1(\mem0[215][0] ), .IN2(n692), .S(n7160), .Q(n18276) );
  AND2X1 U7470 ( .IN1(n7152), .IN2(n7116), .Q(n7160) );
  MUX21X1 U7471 ( .IN1(\mem0[214][7] ), .IN2(n846), .S(n7161), .Q(n18275) );
  MUX21X1 U7472 ( .IN1(\mem0[214][6] ), .IN2(n824), .S(n7161), .Q(n18274) );
  MUX21X1 U7473 ( .IN1(\mem0[214][5] ), .IN2(n802), .S(n7161), .Q(n18273) );
  MUX21X1 U7474 ( .IN1(\mem0[214][4] ), .IN2(n780), .S(n7161), .Q(n18272) );
  MUX21X1 U7475 ( .IN1(\mem0[214][3] ), .IN2(n758), .S(n7161), .Q(n18271) );
  MUX21X1 U7476 ( .IN1(\mem0[214][2] ), .IN2(n736), .S(n7161), .Q(n18270) );
  MUX21X1 U7477 ( .IN1(\mem0[214][1] ), .IN2(n714), .S(n7161), .Q(n18269) );
  MUX21X1 U7478 ( .IN1(\mem0[214][0] ), .IN2(n692), .S(n7161), .Q(n18268) );
  AND2X1 U7479 ( .IN1(n7152), .IN2(n7118), .Q(n7161) );
  MUX21X1 U7480 ( .IN1(\mem0[213][7] ), .IN2(n846), .S(n7162), .Q(n18267) );
  MUX21X1 U7481 ( .IN1(\mem0[213][6] ), .IN2(n824), .S(n7162), .Q(n18266) );
  MUX21X1 U7482 ( .IN1(\mem0[213][5] ), .IN2(n802), .S(n7162), .Q(n18265) );
  MUX21X1 U7483 ( .IN1(\mem0[213][4] ), .IN2(n780), .S(n7162), .Q(n18264) );
  MUX21X1 U7484 ( .IN1(\mem0[213][3] ), .IN2(n758), .S(n7162), .Q(n18263) );
  MUX21X1 U7485 ( .IN1(\mem0[213][2] ), .IN2(n736), .S(n7162), .Q(n18262) );
  MUX21X1 U7486 ( .IN1(\mem0[213][1] ), .IN2(n714), .S(n7162), .Q(n18261) );
  MUX21X1 U7487 ( .IN1(\mem0[213][0] ), .IN2(n692), .S(n7162), .Q(n18260) );
  AND2X1 U7488 ( .IN1(n7152), .IN2(n7120), .Q(n7162) );
  MUX21X1 U7489 ( .IN1(\mem0[212][7] ), .IN2(n846), .S(n7163), .Q(n18259) );
  MUX21X1 U7490 ( .IN1(\mem0[212][6] ), .IN2(n824), .S(n7163), .Q(n18258) );
  MUX21X1 U7491 ( .IN1(\mem0[212][5] ), .IN2(n802), .S(n7163), .Q(n18257) );
  MUX21X1 U7492 ( .IN1(\mem0[212][4] ), .IN2(n780), .S(n7163), .Q(n18256) );
  MUX21X1 U7493 ( .IN1(\mem0[212][3] ), .IN2(n758), .S(n7163), .Q(n18255) );
  MUX21X1 U7494 ( .IN1(\mem0[212][2] ), .IN2(n736), .S(n7163), .Q(n18254) );
  MUX21X1 U7495 ( .IN1(\mem0[212][1] ), .IN2(n714), .S(n7163), .Q(n18253) );
  MUX21X1 U7496 ( .IN1(\mem0[212][0] ), .IN2(n692), .S(n7163), .Q(n18252) );
  AND2X1 U7497 ( .IN1(n7152), .IN2(n7122), .Q(n7163) );
  MUX21X1 U7498 ( .IN1(\mem0[211][7] ), .IN2(n846), .S(n7164), .Q(n18251) );
  MUX21X1 U7499 ( .IN1(\mem0[211][6] ), .IN2(n824), .S(n7164), .Q(n18250) );
  MUX21X1 U7500 ( .IN1(\mem0[211][5] ), .IN2(n802), .S(n7164), .Q(n18249) );
  MUX21X1 U7501 ( .IN1(\mem0[211][4] ), .IN2(n780), .S(n7164), .Q(n18248) );
  MUX21X1 U7502 ( .IN1(\mem0[211][3] ), .IN2(n758), .S(n7164), .Q(n18247) );
  MUX21X1 U7503 ( .IN1(\mem0[211][2] ), .IN2(n736), .S(n7164), .Q(n18246) );
  MUX21X1 U7504 ( .IN1(\mem0[211][1] ), .IN2(n714), .S(n7164), .Q(n18245) );
  MUX21X1 U7505 ( .IN1(\mem0[211][0] ), .IN2(n692), .S(n7164), .Q(n18244) );
  AND2X1 U7506 ( .IN1(n7152), .IN2(n7124), .Q(n7164) );
  MUX21X1 U7507 ( .IN1(\mem0[210][7] ), .IN2(n846), .S(n7165), .Q(n18243) );
  MUX21X1 U7508 ( .IN1(\mem0[210][6] ), .IN2(n824), .S(n7165), .Q(n18242) );
  MUX21X1 U7509 ( .IN1(\mem0[210][5] ), .IN2(n802), .S(n7165), .Q(n18241) );
  MUX21X1 U7510 ( .IN1(\mem0[210][4] ), .IN2(n780), .S(n7165), .Q(n18240) );
  MUX21X1 U7511 ( .IN1(\mem0[210][3] ), .IN2(n758), .S(n7165), .Q(n18239) );
  MUX21X1 U7512 ( .IN1(\mem0[210][2] ), .IN2(n736), .S(n7165), .Q(n18238) );
  MUX21X1 U7513 ( .IN1(\mem0[210][1] ), .IN2(n714), .S(n7165), .Q(n18237) );
  MUX21X1 U7514 ( .IN1(\mem0[210][0] ), .IN2(n692), .S(n7165), .Q(n18236) );
  AND2X1 U7515 ( .IN1(n7152), .IN2(n7126), .Q(n7165) );
  MUX21X1 U7516 ( .IN1(\mem0[209][7] ), .IN2(n846), .S(n7166), .Q(n18235) );
  MUX21X1 U7517 ( .IN1(\mem0[209][6] ), .IN2(n824), .S(n7166), .Q(n18234) );
  MUX21X1 U7518 ( .IN1(\mem0[209][5] ), .IN2(n802), .S(n7166), .Q(n18233) );
  MUX21X1 U7519 ( .IN1(\mem0[209][4] ), .IN2(n780), .S(n7166), .Q(n18232) );
  MUX21X1 U7520 ( .IN1(\mem0[209][3] ), .IN2(n758), .S(n7166), .Q(n18231) );
  MUX21X1 U7521 ( .IN1(\mem0[209][2] ), .IN2(n736), .S(n7166), .Q(n18230) );
  MUX21X1 U7522 ( .IN1(\mem0[209][1] ), .IN2(n714), .S(n7166), .Q(n18229) );
  MUX21X1 U7523 ( .IN1(\mem0[209][0] ), .IN2(n692), .S(n7166), .Q(n18228) );
  AND2X1 U7524 ( .IN1(n7152), .IN2(n7128), .Q(n7166) );
  MUX21X1 U7525 ( .IN1(\mem0[208][7] ), .IN2(n846), .S(n7167), .Q(n18227) );
  MUX21X1 U7526 ( .IN1(\mem0[208][6] ), .IN2(n824), .S(n7167), .Q(n18226) );
  MUX21X1 U7527 ( .IN1(\mem0[208][5] ), .IN2(n802), .S(n7167), .Q(n18225) );
  MUX21X1 U7528 ( .IN1(\mem0[208][4] ), .IN2(n780), .S(n7167), .Q(n18224) );
  MUX21X1 U7529 ( .IN1(\mem0[208][3] ), .IN2(n758), .S(n7167), .Q(n18223) );
  MUX21X1 U7530 ( .IN1(\mem0[208][2] ), .IN2(n736), .S(n7167), .Q(n18222) );
  MUX21X1 U7531 ( .IN1(\mem0[208][1] ), .IN2(n714), .S(n7167), .Q(n18221) );
  MUX21X1 U7532 ( .IN1(\mem0[208][0] ), .IN2(n692), .S(n7167), .Q(n18220) );
  AND2X1 U7533 ( .IN1(n7152), .IN2(n7130), .Q(n7167) );
  AND2X1 U7534 ( .IN1(n7168), .IN2(n7132), .Q(n7152) );
  MUX21X1 U7535 ( .IN1(\mem0[207][7] ), .IN2(n847), .S(n7169), .Q(n18219) );
  MUX21X1 U7536 ( .IN1(\mem0[207][6] ), .IN2(n825), .S(n7169), .Q(n18218) );
  MUX21X1 U7537 ( .IN1(\mem0[207][5] ), .IN2(n803), .S(n7169), .Q(n18217) );
  MUX21X1 U7538 ( .IN1(\mem0[207][4] ), .IN2(n781), .S(n7169), .Q(n18216) );
  MUX21X1 U7539 ( .IN1(\mem0[207][3] ), .IN2(n759), .S(n7169), .Q(n18215) );
  MUX21X1 U7540 ( .IN1(\mem0[207][2] ), .IN2(n737), .S(n7169), .Q(n18214) );
  MUX21X1 U7541 ( .IN1(\mem0[207][1] ), .IN2(n715), .S(n7169), .Q(n18213) );
  MUX21X1 U7542 ( .IN1(\mem0[207][0] ), .IN2(n693), .S(n7169), .Q(n18212) );
  AND2X1 U7543 ( .IN1(n7170), .IN2(n7099), .Q(n7169) );
  MUX21X1 U7544 ( .IN1(\mem0[206][7] ), .IN2(n847), .S(n7171), .Q(n18211) );
  MUX21X1 U7545 ( .IN1(\mem0[206][6] ), .IN2(n825), .S(n7171), .Q(n18210) );
  MUX21X1 U7546 ( .IN1(\mem0[206][5] ), .IN2(n803), .S(n7171), .Q(n18209) );
  MUX21X1 U7547 ( .IN1(\mem0[206][4] ), .IN2(n781), .S(n7171), .Q(n18208) );
  MUX21X1 U7548 ( .IN1(\mem0[206][3] ), .IN2(n759), .S(n7171), .Q(n18207) );
  MUX21X1 U7549 ( .IN1(\mem0[206][2] ), .IN2(n737), .S(n7171), .Q(n18206) );
  MUX21X1 U7550 ( .IN1(\mem0[206][1] ), .IN2(n715), .S(n7171), .Q(n18205) );
  MUX21X1 U7551 ( .IN1(\mem0[206][0] ), .IN2(n693), .S(n7171), .Q(n18204) );
  AND2X1 U7552 ( .IN1(n7170), .IN2(n7102), .Q(n7171) );
  MUX21X1 U7553 ( .IN1(\mem0[205][7] ), .IN2(n847), .S(n7172), .Q(n18203) );
  MUX21X1 U7554 ( .IN1(\mem0[205][6] ), .IN2(n825), .S(n7172), .Q(n18202) );
  MUX21X1 U7555 ( .IN1(\mem0[205][5] ), .IN2(n803), .S(n7172), .Q(n18201) );
  MUX21X1 U7556 ( .IN1(\mem0[205][4] ), .IN2(n781), .S(n7172), .Q(n18200) );
  MUX21X1 U7557 ( .IN1(\mem0[205][3] ), .IN2(n759), .S(n7172), .Q(n18199) );
  MUX21X1 U7558 ( .IN1(\mem0[205][2] ), .IN2(n737), .S(n7172), .Q(n18198) );
  MUX21X1 U7559 ( .IN1(\mem0[205][1] ), .IN2(n715), .S(n7172), .Q(n18197) );
  MUX21X1 U7560 ( .IN1(\mem0[205][0] ), .IN2(n693), .S(n7172), .Q(n18196) );
  AND2X1 U7561 ( .IN1(n7170), .IN2(n7104), .Q(n7172) );
  MUX21X1 U7562 ( .IN1(\mem0[204][7] ), .IN2(n847), .S(n7173), .Q(n18195) );
  MUX21X1 U7563 ( .IN1(\mem0[204][6] ), .IN2(n825), .S(n7173), .Q(n18194) );
  MUX21X1 U7564 ( .IN1(\mem0[204][5] ), .IN2(n803), .S(n7173), .Q(n18193) );
  MUX21X1 U7565 ( .IN1(\mem0[204][4] ), .IN2(n781), .S(n7173), .Q(n18192) );
  MUX21X1 U7566 ( .IN1(\mem0[204][3] ), .IN2(n759), .S(n7173), .Q(n18191) );
  MUX21X1 U7567 ( .IN1(\mem0[204][2] ), .IN2(n737), .S(n7173), .Q(n18190) );
  MUX21X1 U7568 ( .IN1(\mem0[204][1] ), .IN2(n715), .S(n7173), .Q(n18189) );
  MUX21X1 U7569 ( .IN1(\mem0[204][0] ), .IN2(n693), .S(n7173), .Q(n18188) );
  AND2X1 U7570 ( .IN1(n7170), .IN2(n7106), .Q(n7173) );
  MUX21X1 U7571 ( .IN1(\mem0[203][7] ), .IN2(n847), .S(n7174), .Q(n18187) );
  MUX21X1 U7572 ( .IN1(\mem0[203][6] ), .IN2(n825), .S(n7174), .Q(n18186) );
  MUX21X1 U7573 ( .IN1(\mem0[203][5] ), .IN2(n803), .S(n7174), .Q(n18185) );
  MUX21X1 U7574 ( .IN1(\mem0[203][4] ), .IN2(n781), .S(n7174), .Q(n18184) );
  MUX21X1 U7575 ( .IN1(\mem0[203][3] ), .IN2(n759), .S(n7174), .Q(n18183) );
  MUX21X1 U7576 ( .IN1(\mem0[203][2] ), .IN2(n737), .S(n7174), .Q(n18182) );
  MUX21X1 U7577 ( .IN1(\mem0[203][1] ), .IN2(n715), .S(n7174), .Q(n18181) );
  MUX21X1 U7578 ( .IN1(\mem0[203][0] ), .IN2(n693), .S(n7174), .Q(n18180) );
  AND2X1 U7579 ( .IN1(n7170), .IN2(n7108), .Q(n7174) );
  MUX21X1 U7580 ( .IN1(\mem0[202][7] ), .IN2(n847), .S(n7175), .Q(n18179) );
  MUX21X1 U7581 ( .IN1(\mem0[202][6] ), .IN2(n825), .S(n7175), .Q(n18178) );
  MUX21X1 U7582 ( .IN1(\mem0[202][5] ), .IN2(n803), .S(n7175), .Q(n18177) );
  MUX21X1 U7583 ( .IN1(\mem0[202][4] ), .IN2(n781), .S(n7175), .Q(n18176) );
  MUX21X1 U7584 ( .IN1(\mem0[202][3] ), .IN2(n759), .S(n7175), .Q(n18175) );
  MUX21X1 U7585 ( .IN1(\mem0[202][2] ), .IN2(n737), .S(n7175), .Q(n18174) );
  MUX21X1 U7586 ( .IN1(\mem0[202][1] ), .IN2(n715), .S(n7175), .Q(n18173) );
  MUX21X1 U7587 ( .IN1(\mem0[202][0] ), .IN2(n693), .S(n7175), .Q(n18172) );
  AND2X1 U7588 ( .IN1(n7170), .IN2(n7110), .Q(n7175) );
  MUX21X1 U7589 ( .IN1(\mem0[201][7] ), .IN2(n847), .S(n7176), .Q(n18171) );
  MUX21X1 U7590 ( .IN1(\mem0[201][6] ), .IN2(n825), .S(n7176), .Q(n18170) );
  MUX21X1 U7591 ( .IN1(\mem0[201][5] ), .IN2(n803), .S(n7176), .Q(n18169) );
  MUX21X1 U7592 ( .IN1(\mem0[201][4] ), .IN2(n781), .S(n7176), .Q(n18168) );
  MUX21X1 U7593 ( .IN1(\mem0[201][3] ), .IN2(n759), .S(n7176), .Q(n18167) );
  MUX21X1 U7594 ( .IN1(\mem0[201][2] ), .IN2(n737), .S(n7176), .Q(n18166) );
  MUX21X1 U7595 ( .IN1(\mem0[201][1] ), .IN2(n715), .S(n7176), .Q(n18165) );
  MUX21X1 U7596 ( .IN1(\mem0[201][0] ), .IN2(n693), .S(n7176), .Q(n18164) );
  AND2X1 U7597 ( .IN1(n7170), .IN2(n7112), .Q(n7176) );
  MUX21X1 U7598 ( .IN1(\mem0[200][7] ), .IN2(n847), .S(n7177), .Q(n18163) );
  MUX21X1 U7599 ( .IN1(\mem0[200][6] ), .IN2(n825), .S(n7177), .Q(n18162) );
  MUX21X1 U7600 ( .IN1(\mem0[200][5] ), .IN2(n803), .S(n7177), .Q(n18161) );
  MUX21X1 U7601 ( .IN1(\mem0[200][4] ), .IN2(n781), .S(n7177), .Q(n18160) );
  MUX21X1 U7602 ( .IN1(\mem0[200][3] ), .IN2(n759), .S(n7177), .Q(n18159) );
  MUX21X1 U7603 ( .IN1(\mem0[200][2] ), .IN2(n737), .S(n7177), .Q(n18158) );
  MUX21X1 U7604 ( .IN1(\mem0[200][1] ), .IN2(n715), .S(n7177), .Q(n18157) );
  MUX21X1 U7605 ( .IN1(\mem0[200][0] ), .IN2(n693), .S(n7177), .Q(n18156) );
  AND2X1 U7606 ( .IN1(n7170), .IN2(n7114), .Q(n7177) );
  MUX21X1 U7607 ( .IN1(\mem0[199][7] ), .IN2(n847), .S(n7178), .Q(n18155) );
  MUX21X1 U7608 ( .IN1(\mem0[199][6] ), .IN2(n825), .S(n7178), .Q(n18154) );
  MUX21X1 U7609 ( .IN1(\mem0[199][5] ), .IN2(n803), .S(n7178), .Q(n18153) );
  MUX21X1 U7610 ( .IN1(\mem0[199][4] ), .IN2(n781), .S(n7178), .Q(n18152) );
  MUX21X1 U7611 ( .IN1(\mem0[199][3] ), .IN2(n759), .S(n7178), .Q(n18151) );
  MUX21X1 U7612 ( .IN1(\mem0[199][2] ), .IN2(n737), .S(n7178), .Q(n18150) );
  MUX21X1 U7613 ( .IN1(\mem0[199][1] ), .IN2(n715), .S(n7178), .Q(n18149) );
  MUX21X1 U7614 ( .IN1(\mem0[199][0] ), .IN2(n693), .S(n7178), .Q(n18148) );
  AND2X1 U7615 ( .IN1(n7170), .IN2(n7116), .Q(n7178) );
  MUX21X1 U7616 ( .IN1(\mem0[198][7] ), .IN2(n847), .S(n7179), .Q(n18147) );
  MUX21X1 U7617 ( .IN1(\mem0[198][6] ), .IN2(n825), .S(n7179), .Q(n18146) );
  MUX21X1 U7618 ( .IN1(\mem0[198][5] ), .IN2(n803), .S(n7179), .Q(n18145) );
  MUX21X1 U7619 ( .IN1(\mem0[198][4] ), .IN2(n781), .S(n7179), .Q(n18144) );
  MUX21X1 U7620 ( .IN1(\mem0[198][3] ), .IN2(n759), .S(n7179), .Q(n18143) );
  MUX21X1 U7621 ( .IN1(\mem0[198][2] ), .IN2(n737), .S(n7179), .Q(n18142) );
  MUX21X1 U7622 ( .IN1(\mem0[198][1] ), .IN2(n715), .S(n7179), .Q(n18141) );
  MUX21X1 U7623 ( .IN1(\mem0[198][0] ), .IN2(n693), .S(n7179), .Q(n18140) );
  AND2X1 U7624 ( .IN1(n7170), .IN2(n7118), .Q(n7179) );
  MUX21X1 U7625 ( .IN1(\mem0[197][7] ), .IN2(n847), .S(n7180), .Q(n18139) );
  MUX21X1 U7626 ( .IN1(\mem0[197][6] ), .IN2(n825), .S(n7180), .Q(n18138) );
  MUX21X1 U7627 ( .IN1(\mem0[197][5] ), .IN2(n803), .S(n7180), .Q(n18137) );
  MUX21X1 U7628 ( .IN1(\mem0[197][4] ), .IN2(n781), .S(n7180), .Q(n18136) );
  MUX21X1 U7629 ( .IN1(\mem0[197][3] ), .IN2(n759), .S(n7180), .Q(n18135) );
  MUX21X1 U7630 ( .IN1(\mem0[197][2] ), .IN2(n737), .S(n7180), .Q(n18134) );
  MUX21X1 U7631 ( .IN1(\mem0[197][1] ), .IN2(n715), .S(n7180), .Q(n18133) );
  MUX21X1 U7632 ( .IN1(\mem0[197][0] ), .IN2(n693), .S(n7180), .Q(n18132) );
  AND2X1 U7633 ( .IN1(n7170), .IN2(n7120), .Q(n7180) );
  MUX21X1 U7634 ( .IN1(\mem0[196][7] ), .IN2(n847), .S(n7181), .Q(n18131) );
  MUX21X1 U7635 ( .IN1(\mem0[196][6] ), .IN2(n825), .S(n7181), .Q(n18130) );
  MUX21X1 U7636 ( .IN1(\mem0[196][5] ), .IN2(n803), .S(n7181), .Q(n18129) );
  MUX21X1 U7637 ( .IN1(\mem0[196][4] ), .IN2(n781), .S(n7181), .Q(n18128) );
  MUX21X1 U7638 ( .IN1(\mem0[196][3] ), .IN2(n759), .S(n7181), .Q(n18127) );
  MUX21X1 U7639 ( .IN1(\mem0[196][2] ), .IN2(n737), .S(n7181), .Q(n18126) );
  MUX21X1 U7640 ( .IN1(\mem0[196][1] ), .IN2(n715), .S(n7181), .Q(n18125) );
  MUX21X1 U7641 ( .IN1(\mem0[196][0] ), .IN2(n693), .S(n7181), .Q(n18124) );
  AND2X1 U7642 ( .IN1(n7170), .IN2(n7122), .Q(n7181) );
  MUX21X1 U7643 ( .IN1(\mem0[195][7] ), .IN2(n848), .S(n7182), .Q(n18123) );
  MUX21X1 U7644 ( .IN1(\mem0[195][6] ), .IN2(n826), .S(n7182), .Q(n18122) );
  MUX21X1 U7645 ( .IN1(\mem0[195][5] ), .IN2(n804), .S(n7182), .Q(n18121) );
  MUX21X1 U7646 ( .IN1(\mem0[195][4] ), .IN2(n782), .S(n7182), .Q(n18120) );
  MUX21X1 U7647 ( .IN1(\mem0[195][3] ), .IN2(n760), .S(n7182), .Q(n18119) );
  MUX21X1 U7648 ( .IN1(\mem0[195][2] ), .IN2(n738), .S(n7182), .Q(n18118) );
  MUX21X1 U7649 ( .IN1(\mem0[195][1] ), .IN2(n716), .S(n7182), .Q(n18117) );
  MUX21X1 U7650 ( .IN1(\mem0[195][0] ), .IN2(n694), .S(n7182), .Q(n18116) );
  AND2X1 U7651 ( .IN1(n7170), .IN2(n7124), .Q(n7182) );
  MUX21X1 U7652 ( .IN1(\mem0[194][7] ), .IN2(n848), .S(n7183), .Q(n18115) );
  MUX21X1 U7653 ( .IN1(\mem0[194][6] ), .IN2(n826), .S(n7183), .Q(n18114) );
  MUX21X1 U7654 ( .IN1(\mem0[194][5] ), .IN2(n804), .S(n7183), .Q(n18113) );
  MUX21X1 U7655 ( .IN1(\mem0[194][4] ), .IN2(n782), .S(n7183), .Q(n18112) );
  MUX21X1 U7656 ( .IN1(\mem0[194][3] ), .IN2(n760), .S(n7183), .Q(n18111) );
  MUX21X1 U7657 ( .IN1(\mem0[194][2] ), .IN2(n738), .S(n7183), .Q(n18110) );
  MUX21X1 U7658 ( .IN1(\mem0[194][1] ), .IN2(n716), .S(n7183), .Q(n18109) );
  MUX21X1 U7659 ( .IN1(\mem0[194][0] ), .IN2(n694), .S(n7183), .Q(n18108) );
  AND2X1 U7660 ( .IN1(n7170), .IN2(n7126), .Q(n7183) );
  MUX21X1 U7661 ( .IN1(\mem0[193][7] ), .IN2(n848), .S(n7184), .Q(n18107) );
  MUX21X1 U7662 ( .IN1(\mem0[193][6] ), .IN2(n826), .S(n7184), .Q(n18106) );
  MUX21X1 U7663 ( .IN1(\mem0[193][5] ), .IN2(n804), .S(n7184), .Q(n18105) );
  MUX21X1 U7664 ( .IN1(\mem0[193][4] ), .IN2(n782), .S(n7184), .Q(n18104) );
  MUX21X1 U7665 ( .IN1(\mem0[193][3] ), .IN2(n760), .S(n7184), .Q(n18103) );
  MUX21X1 U7666 ( .IN1(\mem0[193][2] ), .IN2(n738), .S(n7184), .Q(n18102) );
  MUX21X1 U7667 ( .IN1(\mem0[193][1] ), .IN2(n716), .S(n7184), .Q(n18101) );
  MUX21X1 U7668 ( .IN1(\mem0[193][0] ), .IN2(n694), .S(n7184), .Q(n18100) );
  AND2X1 U7669 ( .IN1(n7170), .IN2(n7128), .Q(n7184) );
  MUX21X1 U7670 ( .IN1(\mem0[192][7] ), .IN2(n848), .S(n7185), .Q(n18099) );
  MUX21X1 U7671 ( .IN1(\mem0[192][6] ), .IN2(n826), .S(n7185), .Q(n18098) );
  MUX21X1 U7672 ( .IN1(\mem0[192][5] ), .IN2(n804), .S(n7185), .Q(n18097) );
  MUX21X1 U7673 ( .IN1(\mem0[192][4] ), .IN2(n782), .S(n7185), .Q(n18096) );
  MUX21X1 U7674 ( .IN1(\mem0[192][3] ), .IN2(n760), .S(n7185), .Q(n18095) );
  MUX21X1 U7675 ( .IN1(\mem0[192][2] ), .IN2(n738), .S(n7185), .Q(n18094) );
  MUX21X1 U7676 ( .IN1(\mem0[192][1] ), .IN2(n716), .S(n7185), .Q(n18093) );
  MUX21X1 U7677 ( .IN1(\mem0[192][0] ), .IN2(n694), .S(n7185), .Q(n18092) );
  AND2X1 U7678 ( .IN1(n7170), .IN2(n7130), .Q(n7185) );
  AND2X1 U7679 ( .IN1(n7186), .IN2(n7132), .Q(n7170) );
  MUX21X1 U7680 ( .IN1(\mem0[191][7] ), .IN2(n848), .S(n7187), .Q(n18091) );
  MUX21X1 U7681 ( .IN1(\mem0[191][6] ), .IN2(n826), .S(n7187), .Q(n18090) );
  MUX21X1 U7682 ( .IN1(\mem0[191][5] ), .IN2(n804), .S(n7187), .Q(n18089) );
  MUX21X1 U7683 ( .IN1(\mem0[191][4] ), .IN2(n782), .S(n7187), .Q(n18088) );
  MUX21X1 U7684 ( .IN1(\mem0[191][3] ), .IN2(n760), .S(n7187), .Q(n18087) );
  MUX21X1 U7685 ( .IN1(\mem0[191][2] ), .IN2(n738), .S(n7187), .Q(n18086) );
  MUX21X1 U7686 ( .IN1(\mem0[191][1] ), .IN2(n716), .S(n7187), .Q(n18085) );
  MUX21X1 U7687 ( .IN1(\mem0[191][0] ), .IN2(n694), .S(n7187), .Q(n18084) );
  AND2X1 U7688 ( .IN1(n7188), .IN2(n7099), .Q(n7187) );
  MUX21X1 U7689 ( .IN1(\mem0[190][7] ), .IN2(n848), .S(n7189), .Q(n18083) );
  MUX21X1 U7690 ( .IN1(\mem0[190][6] ), .IN2(n826), .S(n7189), .Q(n18082) );
  MUX21X1 U7691 ( .IN1(\mem0[190][5] ), .IN2(n804), .S(n7189), .Q(n18081) );
  MUX21X1 U7692 ( .IN1(\mem0[190][4] ), .IN2(n782), .S(n7189), .Q(n18080) );
  MUX21X1 U7693 ( .IN1(\mem0[190][3] ), .IN2(n760), .S(n7189), .Q(n18079) );
  MUX21X1 U7694 ( .IN1(\mem0[190][2] ), .IN2(n738), .S(n7189), .Q(n18078) );
  MUX21X1 U7695 ( .IN1(\mem0[190][1] ), .IN2(n716), .S(n7189), .Q(n18077) );
  MUX21X1 U7696 ( .IN1(\mem0[190][0] ), .IN2(n694), .S(n7189), .Q(n18076) );
  AND2X1 U7697 ( .IN1(n7188), .IN2(n7102), .Q(n7189) );
  MUX21X1 U7698 ( .IN1(\mem0[189][7] ), .IN2(n848), .S(n7190), .Q(n18075) );
  MUX21X1 U7699 ( .IN1(\mem0[189][6] ), .IN2(n826), .S(n7190), .Q(n18074) );
  MUX21X1 U7700 ( .IN1(\mem0[189][5] ), .IN2(n804), .S(n7190), .Q(n18073) );
  MUX21X1 U7701 ( .IN1(\mem0[189][4] ), .IN2(n782), .S(n7190), .Q(n18072) );
  MUX21X1 U7702 ( .IN1(\mem0[189][3] ), .IN2(n760), .S(n7190), .Q(n18071) );
  MUX21X1 U7703 ( .IN1(\mem0[189][2] ), .IN2(n738), .S(n7190), .Q(n18070) );
  MUX21X1 U7704 ( .IN1(\mem0[189][1] ), .IN2(n716), .S(n7190), .Q(n18069) );
  MUX21X1 U7705 ( .IN1(\mem0[189][0] ), .IN2(n694), .S(n7190), .Q(n18068) );
  AND2X1 U7706 ( .IN1(n7188), .IN2(n7104), .Q(n7190) );
  MUX21X1 U7707 ( .IN1(\mem0[188][7] ), .IN2(n848), .S(n7191), .Q(n18067) );
  MUX21X1 U7708 ( .IN1(\mem0[188][6] ), .IN2(n826), .S(n7191), .Q(n18066) );
  MUX21X1 U7709 ( .IN1(\mem0[188][5] ), .IN2(n804), .S(n7191), .Q(n18065) );
  MUX21X1 U7710 ( .IN1(\mem0[188][4] ), .IN2(n782), .S(n7191), .Q(n18064) );
  MUX21X1 U7711 ( .IN1(\mem0[188][3] ), .IN2(n760), .S(n7191), .Q(n18063) );
  MUX21X1 U7712 ( .IN1(\mem0[188][2] ), .IN2(n738), .S(n7191), .Q(n18062) );
  MUX21X1 U7713 ( .IN1(\mem0[188][1] ), .IN2(n716), .S(n7191), .Q(n18061) );
  MUX21X1 U7714 ( .IN1(\mem0[188][0] ), .IN2(n694), .S(n7191), .Q(n18060) );
  AND2X1 U7715 ( .IN1(n7188), .IN2(n7106), .Q(n7191) );
  MUX21X1 U7716 ( .IN1(\mem0[187][7] ), .IN2(n848), .S(n7192), .Q(n18059) );
  MUX21X1 U7717 ( .IN1(\mem0[187][6] ), .IN2(n826), .S(n7192), .Q(n18058) );
  MUX21X1 U7718 ( .IN1(\mem0[187][5] ), .IN2(n804), .S(n7192), .Q(n18057) );
  MUX21X1 U7719 ( .IN1(\mem0[187][4] ), .IN2(n782), .S(n7192), .Q(n18056) );
  MUX21X1 U7720 ( .IN1(\mem0[187][3] ), .IN2(n760), .S(n7192), .Q(n18055) );
  MUX21X1 U7721 ( .IN1(\mem0[187][2] ), .IN2(n738), .S(n7192), .Q(n18054) );
  MUX21X1 U7722 ( .IN1(\mem0[187][1] ), .IN2(n716), .S(n7192), .Q(n18053) );
  MUX21X1 U7723 ( .IN1(\mem0[187][0] ), .IN2(n694), .S(n7192), .Q(n18052) );
  AND2X1 U7724 ( .IN1(n7188), .IN2(n7108), .Q(n7192) );
  MUX21X1 U7725 ( .IN1(\mem0[186][7] ), .IN2(n848), .S(n7193), .Q(n18051) );
  MUX21X1 U7726 ( .IN1(\mem0[186][6] ), .IN2(n826), .S(n7193), .Q(n18050) );
  MUX21X1 U7727 ( .IN1(\mem0[186][5] ), .IN2(n804), .S(n7193), .Q(n18049) );
  MUX21X1 U7728 ( .IN1(\mem0[186][4] ), .IN2(n782), .S(n7193), .Q(n18048) );
  MUX21X1 U7729 ( .IN1(\mem0[186][3] ), .IN2(n760), .S(n7193), .Q(n18047) );
  MUX21X1 U7730 ( .IN1(\mem0[186][2] ), .IN2(n738), .S(n7193), .Q(n18046) );
  MUX21X1 U7731 ( .IN1(\mem0[186][1] ), .IN2(n716), .S(n7193), .Q(n18045) );
  MUX21X1 U7732 ( .IN1(\mem0[186][0] ), .IN2(n694), .S(n7193), .Q(n18044) );
  AND2X1 U7733 ( .IN1(n7188), .IN2(n7110), .Q(n7193) );
  MUX21X1 U7734 ( .IN1(\mem0[185][7] ), .IN2(n848), .S(n7194), .Q(n18043) );
  MUX21X1 U7735 ( .IN1(\mem0[185][6] ), .IN2(n826), .S(n7194), .Q(n18042) );
  MUX21X1 U7736 ( .IN1(\mem0[185][5] ), .IN2(n804), .S(n7194), .Q(n18041) );
  MUX21X1 U7737 ( .IN1(\mem0[185][4] ), .IN2(n782), .S(n7194), .Q(n18040) );
  MUX21X1 U7738 ( .IN1(\mem0[185][3] ), .IN2(n760), .S(n7194), .Q(n18039) );
  MUX21X1 U7739 ( .IN1(\mem0[185][2] ), .IN2(n738), .S(n7194), .Q(n18038) );
  MUX21X1 U7740 ( .IN1(\mem0[185][1] ), .IN2(n716), .S(n7194), .Q(n18037) );
  MUX21X1 U7741 ( .IN1(\mem0[185][0] ), .IN2(n694), .S(n7194), .Q(n18036) );
  AND2X1 U7742 ( .IN1(n7188), .IN2(n7112), .Q(n7194) );
  MUX21X1 U7743 ( .IN1(\mem0[184][7] ), .IN2(n848), .S(n7195), .Q(n18035) );
  MUX21X1 U7744 ( .IN1(\mem0[184][6] ), .IN2(n826), .S(n7195), .Q(n18034) );
  MUX21X1 U7745 ( .IN1(\mem0[184][5] ), .IN2(n804), .S(n7195), .Q(n18033) );
  MUX21X1 U7746 ( .IN1(\mem0[184][4] ), .IN2(n782), .S(n7195), .Q(n18032) );
  MUX21X1 U7747 ( .IN1(\mem0[184][3] ), .IN2(n760), .S(n7195), .Q(n18031) );
  MUX21X1 U7748 ( .IN1(\mem0[184][2] ), .IN2(n738), .S(n7195), .Q(n18030) );
  MUX21X1 U7749 ( .IN1(\mem0[184][1] ), .IN2(n716), .S(n7195), .Q(n18029) );
  MUX21X1 U7750 ( .IN1(\mem0[184][0] ), .IN2(n694), .S(n7195), .Q(n18028) );
  AND2X1 U7751 ( .IN1(n7188), .IN2(n7114), .Q(n7195) );
  MUX21X1 U7752 ( .IN1(\mem0[183][7] ), .IN2(n849), .S(n7196), .Q(n18027) );
  MUX21X1 U7753 ( .IN1(\mem0[183][6] ), .IN2(n827), .S(n7196), .Q(n18026) );
  MUX21X1 U7754 ( .IN1(\mem0[183][5] ), .IN2(n805), .S(n7196), .Q(n18025) );
  MUX21X1 U7755 ( .IN1(\mem0[183][4] ), .IN2(n783), .S(n7196), .Q(n18024) );
  MUX21X1 U7756 ( .IN1(\mem0[183][3] ), .IN2(n761), .S(n7196), .Q(n18023) );
  MUX21X1 U7757 ( .IN1(\mem0[183][2] ), .IN2(n739), .S(n7196), .Q(n18022) );
  MUX21X1 U7758 ( .IN1(\mem0[183][1] ), .IN2(n717), .S(n7196), .Q(n18021) );
  MUX21X1 U7759 ( .IN1(\mem0[183][0] ), .IN2(n695), .S(n7196), .Q(n18020) );
  AND2X1 U7760 ( .IN1(n7188), .IN2(n7116), .Q(n7196) );
  MUX21X1 U7761 ( .IN1(\mem0[182][7] ), .IN2(n849), .S(n7197), .Q(n18019) );
  MUX21X1 U7762 ( .IN1(\mem0[182][6] ), .IN2(n827), .S(n7197), .Q(n18018) );
  MUX21X1 U7763 ( .IN1(\mem0[182][5] ), .IN2(n805), .S(n7197), .Q(n18017) );
  MUX21X1 U7764 ( .IN1(\mem0[182][4] ), .IN2(n783), .S(n7197), .Q(n18016) );
  MUX21X1 U7765 ( .IN1(\mem0[182][3] ), .IN2(n761), .S(n7197), .Q(n18015) );
  MUX21X1 U7766 ( .IN1(\mem0[182][2] ), .IN2(n739), .S(n7197), .Q(n18014) );
  MUX21X1 U7767 ( .IN1(\mem0[182][1] ), .IN2(n717), .S(n7197), .Q(n18013) );
  MUX21X1 U7768 ( .IN1(\mem0[182][0] ), .IN2(n695), .S(n7197), .Q(n18012) );
  AND2X1 U7769 ( .IN1(n7188), .IN2(n7118), .Q(n7197) );
  MUX21X1 U7770 ( .IN1(\mem0[181][7] ), .IN2(n849), .S(n7198), .Q(n18011) );
  MUX21X1 U7771 ( .IN1(\mem0[181][6] ), .IN2(n827), .S(n7198), .Q(n18010) );
  MUX21X1 U7772 ( .IN1(\mem0[181][5] ), .IN2(n805), .S(n7198), .Q(n18009) );
  MUX21X1 U7773 ( .IN1(\mem0[181][4] ), .IN2(n783), .S(n7198), .Q(n18008) );
  MUX21X1 U7774 ( .IN1(\mem0[181][3] ), .IN2(n761), .S(n7198), .Q(n18007) );
  MUX21X1 U7775 ( .IN1(\mem0[181][2] ), .IN2(n739), .S(n7198), .Q(n18006) );
  MUX21X1 U7776 ( .IN1(\mem0[181][1] ), .IN2(n717), .S(n7198), .Q(n18005) );
  MUX21X1 U7777 ( .IN1(\mem0[181][0] ), .IN2(n695), .S(n7198), .Q(n18004) );
  AND2X1 U7778 ( .IN1(n7188), .IN2(n7120), .Q(n7198) );
  MUX21X1 U7779 ( .IN1(\mem0[180][7] ), .IN2(n849), .S(n7199), .Q(n18003) );
  MUX21X1 U7780 ( .IN1(\mem0[180][6] ), .IN2(n827), .S(n7199), .Q(n18002) );
  MUX21X1 U7781 ( .IN1(\mem0[180][5] ), .IN2(n805), .S(n7199), .Q(n18001) );
  MUX21X1 U7782 ( .IN1(\mem0[180][4] ), .IN2(n783), .S(n7199), .Q(n18000) );
  MUX21X1 U7783 ( .IN1(\mem0[180][3] ), .IN2(n761), .S(n7199), .Q(n17999) );
  MUX21X1 U7784 ( .IN1(\mem0[180][2] ), .IN2(n739), .S(n7199), .Q(n17998) );
  MUX21X1 U7785 ( .IN1(\mem0[180][1] ), .IN2(n717), .S(n7199), .Q(n17997) );
  MUX21X1 U7786 ( .IN1(\mem0[180][0] ), .IN2(n695), .S(n7199), .Q(n17996) );
  AND2X1 U7787 ( .IN1(n7188), .IN2(n7122), .Q(n7199) );
  MUX21X1 U7788 ( .IN1(\mem0[179][7] ), .IN2(n849), .S(n7200), .Q(n17995) );
  MUX21X1 U7789 ( .IN1(\mem0[179][6] ), .IN2(n827), .S(n7200), .Q(n17994) );
  MUX21X1 U7790 ( .IN1(\mem0[179][5] ), .IN2(n805), .S(n7200), .Q(n17993) );
  MUX21X1 U7791 ( .IN1(\mem0[179][4] ), .IN2(n783), .S(n7200), .Q(n17992) );
  MUX21X1 U7792 ( .IN1(\mem0[179][3] ), .IN2(n761), .S(n7200), .Q(n17991) );
  MUX21X1 U7793 ( .IN1(\mem0[179][2] ), .IN2(n739), .S(n7200), .Q(n17990) );
  MUX21X1 U7794 ( .IN1(\mem0[179][1] ), .IN2(n717), .S(n7200), .Q(n17989) );
  MUX21X1 U7795 ( .IN1(\mem0[179][0] ), .IN2(n695), .S(n7200), .Q(n17988) );
  AND2X1 U7796 ( .IN1(n7188), .IN2(n7124), .Q(n7200) );
  MUX21X1 U7797 ( .IN1(\mem0[178][7] ), .IN2(n849), .S(n7201), .Q(n17987) );
  MUX21X1 U7798 ( .IN1(\mem0[178][6] ), .IN2(n827), .S(n7201), .Q(n17986) );
  MUX21X1 U7799 ( .IN1(\mem0[178][5] ), .IN2(n805), .S(n7201), .Q(n17985) );
  MUX21X1 U7800 ( .IN1(\mem0[178][4] ), .IN2(n783), .S(n7201), .Q(n17984) );
  MUX21X1 U7801 ( .IN1(\mem0[178][3] ), .IN2(n761), .S(n7201), .Q(n17983) );
  MUX21X1 U7802 ( .IN1(\mem0[178][2] ), .IN2(n739), .S(n7201), .Q(n17982) );
  MUX21X1 U7803 ( .IN1(\mem0[178][1] ), .IN2(n717), .S(n7201), .Q(n17981) );
  MUX21X1 U7804 ( .IN1(\mem0[178][0] ), .IN2(n695), .S(n7201), .Q(n17980) );
  AND2X1 U7805 ( .IN1(n7188), .IN2(n7126), .Q(n7201) );
  MUX21X1 U7806 ( .IN1(\mem0[177][7] ), .IN2(n849), .S(n7202), .Q(n17979) );
  MUX21X1 U7807 ( .IN1(\mem0[177][6] ), .IN2(n827), .S(n7202), .Q(n17978) );
  MUX21X1 U7808 ( .IN1(\mem0[177][5] ), .IN2(n805), .S(n7202), .Q(n17977) );
  MUX21X1 U7809 ( .IN1(\mem0[177][4] ), .IN2(n783), .S(n7202), .Q(n17976) );
  MUX21X1 U7810 ( .IN1(\mem0[177][3] ), .IN2(n761), .S(n7202), .Q(n17975) );
  MUX21X1 U7811 ( .IN1(\mem0[177][2] ), .IN2(n739), .S(n7202), .Q(n17974) );
  MUX21X1 U7812 ( .IN1(\mem0[177][1] ), .IN2(n717), .S(n7202), .Q(n17973) );
  MUX21X1 U7813 ( .IN1(\mem0[177][0] ), .IN2(n695), .S(n7202), .Q(n17972) );
  AND2X1 U7814 ( .IN1(n7188), .IN2(n7128), .Q(n7202) );
  MUX21X1 U7815 ( .IN1(\mem0[176][7] ), .IN2(n849), .S(n7203), .Q(n17971) );
  MUX21X1 U7816 ( .IN1(\mem0[176][6] ), .IN2(n827), .S(n7203), .Q(n17970) );
  MUX21X1 U7817 ( .IN1(\mem0[176][5] ), .IN2(n805), .S(n7203), .Q(n17969) );
  MUX21X1 U7818 ( .IN1(\mem0[176][4] ), .IN2(n783), .S(n7203), .Q(n17968) );
  MUX21X1 U7819 ( .IN1(\mem0[176][3] ), .IN2(n761), .S(n7203), .Q(n17967) );
  MUX21X1 U7820 ( .IN1(\mem0[176][2] ), .IN2(n739), .S(n7203), .Q(n17966) );
  MUX21X1 U7821 ( .IN1(\mem0[176][1] ), .IN2(n717), .S(n7203), .Q(n17965) );
  MUX21X1 U7822 ( .IN1(\mem0[176][0] ), .IN2(n695), .S(n7203), .Q(n17964) );
  AND2X1 U7823 ( .IN1(n7188), .IN2(n7130), .Q(n7203) );
  AND2X1 U7824 ( .IN1(n7204), .IN2(n7132), .Q(n7188) );
  MUX21X1 U7825 ( .IN1(\mem0[175][7] ), .IN2(n849), .S(n7205), .Q(n17963) );
  MUX21X1 U7826 ( .IN1(\mem0[175][6] ), .IN2(n827), .S(n7205), .Q(n17962) );
  MUX21X1 U7827 ( .IN1(\mem0[175][5] ), .IN2(n805), .S(n7205), .Q(n17961) );
  MUX21X1 U7828 ( .IN1(\mem0[175][4] ), .IN2(n783), .S(n7205), .Q(n17960) );
  MUX21X1 U7829 ( .IN1(\mem0[175][3] ), .IN2(n761), .S(n7205), .Q(n17959) );
  MUX21X1 U7830 ( .IN1(\mem0[175][2] ), .IN2(n739), .S(n7205), .Q(n17958) );
  MUX21X1 U7831 ( .IN1(\mem0[175][1] ), .IN2(n717), .S(n7205), .Q(n17957) );
  MUX21X1 U7832 ( .IN1(\mem0[175][0] ), .IN2(n695), .S(n7205), .Q(n17956) );
  AND2X1 U7833 ( .IN1(n7206), .IN2(n7099), .Q(n7205) );
  MUX21X1 U7834 ( .IN1(\mem0[174][7] ), .IN2(n849), .S(n7207), .Q(n17955) );
  MUX21X1 U7835 ( .IN1(\mem0[174][6] ), .IN2(n827), .S(n7207), .Q(n17954) );
  MUX21X1 U7836 ( .IN1(\mem0[174][5] ), .IN2(n805), .S(n7207), .Q(n17953) );
  MUX21X1 U7837 ( .IN1(\mem0[174][4] ), .IN2(n783), .S(n7207), .Q(n17952) );
  MUX21X1 U7838 ( .IN1(\mem0[174][3] ), .IN2(n761), .S(n7207), .Q(n17951) );
  MUX21X1 U7839 ( .IN1(\mem0[174][2] ), .IN2(n739), .S(n7207), .Q(n17950) );
  MUX21X1 U7840 ( .IN1(\mem0[174][1] ), .IN2(n717), .S(n7207), .Q(n17949) );
  MUX21X1 U7841 ( .IN1(\mem0[174][0] ), .IN2(n695), .S(n7207), .Q(n17948) );
  AND2X1 U7842 ( .IN1(n7206), .IN2(n7102), .Q(n7207) );
  MUX21X1 U7843 ( .IN1(\mem0[173][7] ), .IN2(n849), .S(n7208), .Q(n17947) );
  MUX21X1 U7844 ( .IN1(\mem0[173][6] ), .IN2(n827), .S(n7208), .Q(n17946) );
  MUX21X1 U7845 ( .IN1(\mem0[173][5] ), .IN2(n805), .S(n7208), .Q(n17945) );
  MUX21X1 U7846 ( .IN1(\mem0[173][4] ), .IN2(n783), .S(n7208), .Q(n17944) );
  MUX21X1 U7847 ( .IN1(\mem0[173][3] ), .IN2(n761), .S(n7208), .Q(n17943) );
  MUX21X1 U7848 ( .IN1(\mem0[173][2] ), .IN2(n739), .S(n7208), .Q(n17942) );
  MUX21X1 U7849 ( .IN1(\mem0[173][1] ), .IN2(n717), .S(n7208), .Q(n17941) );
  MUX21X1 U7850 ( .IN1(\mem0[173][0] ), .IN2(n695), .S(n7208), .Q(n17940) );
  AND2X1 U7851 ( .IN1(n7206), .IN2(n7104), .Q(n7208) );
  MUX21X1 U7852 ( .IN1(\mem0[172][7] ), .IN2(n849), .S(n7209), .Q(n17939) );
  MUX21X1 U7853 ( .IN1(\mem0[172][6] ), .IN2(n827), .S(n7209), .Q(n17938) );
  MUX21X1 U7854 ( .IN1(\mem0[172][5] ), .IN2(n805), .S(n7209), .Q(n17937) );
  MUX21X1 U7855 ( .IN1(\mem0[172][4] ), .IN2(n783), .S(n7209), .Q(n17936) );
  MUX21X1 U7856 ( .IN1(\mem0[172][3] ), .IN2(n761), .S(n7209), .Q(n17935) );
  MUX21X1 U7857 ( .IN1(\mem0[172][2] ), .IN2(n739), .S(n7209), .Q(n17934) );
  MUX21X1 U7858 ( .IN1(\mem0[172][1] ), .IN2(n717), .S(n7209), .Q(n17933) );
  MUX21X1 U7859 ( .IN1(\mem0[172][0] ), .IN2(n695), .S(n7209), .Q(n17932) );
  AND2X1 U7860 ( .IN1(n7206), .IN2(n7106), .Q(n7209) );
  MUX21X1 U7861 ( .IN1(\mem0[171][7] ), .IN2(n850), .S(n7210), .Q(n17931) );
  MUX21X1 U7862 ( .IN1(\mem0[171][6] ), .IN2(n828), .S(n7210), .Q(n17930) );
  MUX21X1 U7863 ( .IN1(\mem0[171][5] ), .IN2(n806), .S(n7210), .Q(n17929) );
  MUX21X1 U7864 ( .IN1(\mem0[171][4] ), .IN2(n784), .S(n7210), .Q(n17928) );
  MUX21X1 U7865 ( .IN1(\mem0[171][3] ), .IN2(n762), .S(n7210), .Q(n17927) );
  MUX21X1 U7866 ( .IN1(\mem0[171][2] ), .IN2(n740), .S(n7210), .Q(n17926) );
  MUX21X1 U7867 ( .IN1(\mem0[171][1] ), .IN2(n718), .S(n7210), .Q(n17925) );
  MUX21X1 U7868 ( .IN1(\mem0[171][0] ), .IN2(n696), .S(n7210), .Q(n17924) );
  AND2X1 U7869 ( .IN1(n7206), .IN2(n7108), .Q(n7210) );
  MUX21X1 U7870 ( .IN1(\mem0[170][7] ), .IN2(n850), .S(n7211), .Q(n17923) );
  MUX21X1 U7871 ( .IN1(\mem0[170][6] ), .IN2(n828), .S(n7211), .Q(n17922) );
  MUX21X1 U7872 ( .IN1(\mem0[170][5] ), .IN2(n806), .S(n7211), .Q(n17921) );
  MUX21X1 U7873 ( .IN1(\mem0[170][4] ), .IN2(n784), .S(n7211), .Q(n17920) );
  MUX21X1 U7874 ( .IN1(\mem0[170][3] ), .IN2(n762), .S(n7211), .Q(n17919) );
  MUX21X1 U7875 ( .IN1(\mem0[170][2] ), .IN2(n740), .S(n7211), .Q(n17918) );
  MUX21X1 U7876 ( .IN1(\mem0[170][1] ), .IN2(n718), .S(n7211), .Q(n17917) );
  MUX21X1 U7877 ( .IN1(\mem0[170][0] ), .IN2(n696), .S(n7211), .Q(n17916) );
  AND2X1 U7878 ( .IN1(n7206), .IN2(n7110), .Q(n7211) );
  MUX21X1 U7879 ( .IN1(\mem0[169][7] ), .IN2(n850), .S(n7212), .Q(n17915) );
  MUX21X1 U7880 ( .IN1(\mem0[169][6] ), .IN2(n828), .S(n7212), .Q(n17914) );
  MUX21X1 U7881 ( .IN1(\mem0[169][5] ), .IN2(n806), .S(n7212), .Q(n17913) );
  MUX21X1 U7882 ( .IN1(\mem0[169][4] ), .IN2(n784), .S(n7212), .Q(n17912) );
  MUX21X1 U7883 ( .IN1(\mem0[169][3] ), .IN2(n762), .S(n7212), .Q(n17911) );
  MUX21X1 U7884 ( .IN1(\mem0[169][2] ), .IN2(n740), .S(n7212), .Q(n17910) );
  MUX21X1 U7885 ( .IN1(\mem0[169][1] ), .IN2(n718), .S(n7212), .Q(n17909) );
  MUX21X1 U7886 ( .IN1(\mem0[169][0] ), .IN2(n696), .S(n7212), .Q(n17908) );
  AND2X1 U7887 ( .IN1(n7206), .IN2(n7112), .Q(n7212) );
  MUX21X1 U7888 ( .IN1(\mem0[168][7] ), .IN2(n850), .S(n7213), .Q(n17907) );
  MUX21X1 U7889 ( .IN1(\mem0[168][6] ), .IN2(n828), .S(n7213), .Q(n17906) );
  MUX21X1 U7890 ( .IN1(\mem0[168][5] ), .IN2(n806), .S(n7213), .Q(n17905) );
  MUX21X1 U7891 ( .IN1(\mem0[168][4] ), .IN2(n784), .S(n7213), .Q(n17904) );
  MUX21X1 U7892 ( .IN1(\mem0[168][3] ), .IN2(n762), .S(n7213), .Q(n17903) );
  MUX21X1 U7893 ( .IN1(\mem0[168][2] ), .IN2(n740), .S(n7213), .Q(n17902) );
  MUX21X1 U7894 ( .IN1(\mem0[168][1] ), .IN2(n718), .S(n7213), .Q(n17901) );
  MUX21X1 U7895 ( .IN1(\mem0[168][0] ), .IN2(n696), .S(n7213), .Q(n17900) );
  AND2X1 U7896 ( .IN1(n7206), .IN2(n7114), .Q(n7213) );
  MUX21X1 U7897 ( .IN1(\mem0[167][7] ), .IN2(n850), .S(n7214), .Q(n17899) );
  MUX21X1 U7898 ( .IN1(\mem0[167][6] ), .IN2(n828), .S(n7214), .Q(n17898) );
  MUX21X1 U7899 ( .IN1(\mem0[167][5] ), .IN2(n806), .S(n7214), .Q(n17897) );
  MUX21X1 U7900 ( .IN1(\mem0[167][4] ), .IN2(n784), .S(n7214), .Q(n17896) );
  MUX21X1 U7901 ( .IN1(\mem0[167][3] ), .IN2(n762), .S(n7214), .Q(n17895) );
  MUX21X1 U7902 ( .IN1(\mem0[167][2] ), .IN2(n740), .S(n7214), .Q(n17894) );
  MUX21X1 U7903 ( .IN1(\mem0[167][1] ), .IN2(n718), .S(n7214), .Q(n17893) );
  MUX21X1 U7904 ( .IN1(\mem0[167][0] ), .IN2(n696), .S(n7214), .Q(n17892) );
  AND2X1 U7905 ( .IN1(n7206), .IN2(n7116), .Q(n7214) );
  MUX21X1 U7906 ( .IN1(\mem0[166][7] ), .IN2(n850), .S(n7215), .Q(n17891) );
  MUX21X1 U7907 ( .IN1(\mem0[166][6] ), .IN2(n828), .S(n7215), .Q(n17890) );
  MUX21X1 U7908 ( .IN1(\mem0[166][5] ), .IN2(n806), .S(n7215), .Q(n17889) );
  MUX21X1 U7909 ( .IN1(\mem0[166][4] ), .IN2(n784), .S(n7215), .Q(n17888) );
  MUX21X1 U7910 ( .IN1(\mem0[166][3] ), .IN2(n762), .S(n7215), .Q(n17887) );
  MUX21X1 U7911 ( .IN1(\mem0[166][2] ), .IN2(n740), .S(n7215), .Q(n17886) );
  MUX21X1 U7912 ( .IN1(\mem0[166][1] ), .IN2(n718), .S(n7215), .Q(n17885) );
  MUX21X1 U7913 ( .IN1(\mem0[166][0] ), .IN2(n696), .S(n7215), .Q(n17884) );
  AND2X1 U7914 ( .IN1(n7206), .IN2(n7118), .Q(n7215) );
  MUX21X1 U7915 ( .IN1(\mem0[165][7] ), .IN2(n850), .S(n7216), .Q(n17883) );
  MUX21X1 U7916 ( .IN1(\mem0[165][6] ), .IN2(n828), .S(n7216), .Q(n17882) );
  MUX21X1 U7917 ( .IN1(\mem0[165][5] ), .IN2(n806), .S(n7216), .Q(n17881) );
  MUX21X1 U7918 ( .IN1(\mem0[165][4] ), .IN2(n784), .S(n7216), .Q(n17880) );
  MUX21X1 U7919 ( .IN1(\mem0[165][3] ), .IN2(n762), .S(n7216), .Q(n17879) );
  MUX21X1 U7920 ( .IN1(\mem0[165][2] ), .IN2(n740), .S(n7216), .Q(n17878) );
  MUX21X1 U7921 ( .IN1(\mem0[165][1] ), .IN2(n718), .S(n7216), .Q(n17877) );
  MUX21X1 U7922 ( .IN1(\mem0[165][0] ), .IN2(n696), .S(n7216), .Q(n17876) );
  AND2X1 U7923 ( .IN1(n7206), .IN2(n7120), .Q(n7216) );
  MUX21X1 U7924 ( .IN1(\mem0[164][7] ), .IN2(n850), .S(n7217), .Q(n17875) );
  MUX21X1 U7925 ( .IN1(\mem0[164][6] ), .IN2(n828), .S(n7217), .Q(n17874) );
  MUX21X1 U7926 ( .IN1(\mem0[164][5] ), .IN2(n806), .S(n7217), .Q(n17873) );
  MUX21X1 U7927 ( .IN1(\mem0[164][4] ), .IN2(n784), .S(n7217), .Q(n17872) );
  MUX21X1 U7928 ( .IN1(\mem0[164][3] ), .IN2(n762), .S(n7217), .Q(n17871) );
  MUX21X1 U7929 ( .IN1(\mem0[164][2] ), .IN2(n740), .S(n7217), .Q(n17870) );
  MUX21X1 U7930 ( .IN1(\mem0[164][1] ), .IN2(n718), .S(n7217), .Q(n17869) );
  MUX21X1 U7931 ( .IN1(\mem0[164][0] ), .IN2(n696), .S(n7217), .Q(n17868) );
  AND2X1 U7932 ( .IN1(n7206), .IN2(n7122), .Q(n7217) );
  MUX21X1 U7933 ( .IN1(\mem0[163][7] ), .IN2(n850), .S(n7218), .Q(n17867) );
  MUX21X1 U7934 ( .IN1(\mem0[163][6] ), .IN2(n828), .S(n7218), .Q(n17866) );
  MUX21X1 U7935 ( .IN1(\mem0[163][5] ), .IN2(n806), .S(n7218), .Q(n17865) );
  MUX21X1 U7936 ( .IN1(\mem0[163][4] ), .IN2(n784), .S(n7218), .Q(n17864) );
  MUX21X1 U7937 ( .IN1(\mem0[163][3] ), .IN2(n762), .S(n7218), .Q(n17863) );
  MUX21X1 U7938 ( .IN1(\mem0[163][2] ), .IN2(n740), .S(n7218), .Q(n17862) );
  MUX21X1 U7939 ( .IN1(\mem0[163][1] ), .IN2(n718), .S(n7218), .Q(n17861) );
  MUX21X1 U7940 ( .IN1(\mem0[163][0] ), .IN2(n696), .S(n7218), .Q(n17860) );
  AND2X1 U7941 ( .IN1(n7206), .IN2(n7124), .Q(n7218) );
  MUX21X1 U7942 ( .IN1(\mem0[162][7] ), .IN2(n850), .S(n7219), .Q(n17859) );
  MUX21X1 U7943 ( .IN1(\mem0[162][6] ), .IN2(n828), .S(n7219), .Q(n17858) );
  MUX21X1 U7944 ( .IN1(\mem0[162][5] ), .IN2(n806), .S(n7219), .Q(n17857) );
  MUX21X1 U7945 ( .IN1(\mem0[162][4] ), .IN2(n784), .S(n7219), .Q(n17856) );
  MUX21X1 U7946 ( .IN1(\mem0[162][3] ), .IN2(n762), .S(n7219), .Q(n17855) );
  MUX21X1 U7947 ( .IN1(\mem0[162][2] ), .IN2(n740), .S(n7219), .Q(n17854) );
  MUX21X1 U7948 ( .IN1(\mem0[162][1] ), .IN2(n718), .S(n7219), .Q(n17853) );
  MUX21X1 U7949 ( .IN1(\mem0[162][0] ), .IN2(n696), .S(n7219), .Q(n17852) );
  AND2X1 U7950 ( .IN1(n7206), .IN2(n7126), .Q(n7219) );
  MUX21X1 U7951 ( .IN1(\mem0[161][7] ), .IN2(n850), .S(n7220), .Q(n17851) );
  MUX21X1 U7952 ( .IN1(\mem0[161][6] ), .IN2(n828), .S(n7220), .Q(n17850) );
  MUX21X1 U7953 ( .IN1(\mem0[161][5] ), .IN2(n806), .S(n7220), .Q(n17849) );
  MUX21X1 U7954 ( .IN1(\mem0[161][4] ), .IN2(n784), .S(n7220), .Q(n17848) );
  MUX21X1 U7955 ( .IN1(\mem0[161][3] ), .IN2(n762), .S(n7220), .Q(n17847) );
  MUX21X1 U7956 ( .IN1(\mem0[161][2] ), .IN2(n740), .S(n7220), .Q(n17846) );
  MUX21X1 U7957 ( .IN1(\mem0[161][1] ), .IN2(n718), .S(n7220), .Q(n17845) );
  MUX21X1 U7958 ( .IN1(\mem0[161][0] ), .IN2(n696), .S(n7220), .Q(n17844) );
  AND2X1 U7959 ( .IN1(n7206), .IN2(n7128), .Q(n7220) );
  MUX21X1 U7960 ( .IN1(\mem0[160][7] ), .IN2(n850), .S(n7221), .Q(n17843) );
  MUX21X1 U7961 ( .IN1(\mem0[160][6] ), .IN2(n828), .S(n7221), .Q(n17842) );
  MUX21X1 U7962 ( .IN1(\mem0[160][5] ), .IN2(n806), .S(n7221), .Q(n17841) );
  MUX21X1 U7963 ( .IN1(\mem0[160][4] ), .IN2(n784), .S(n7221), .Q(n17840) );
  MUX21X1 U7964 ( .IN1(\mem0[160][3] ), .IN2(n762), .S(n7221), .Q(n17839) );
  MUX21X1 U7965 ( .IN1(\mem0[160][2] ), .IN2(n740), .S(n7221), .Q(n17838) );
  MUX21X1 U7966 ( .IN1(\mem0[160][1] ), .IN2(n718), .S(n7221), .Q(n17837) );
  MUX21X1 U7967 ( .IN1(\mem0[160][0] ), .IN2(n696), .S(n7221), .Q(n17836) );
  AND2X1 U7968 ( .IN1(n7206), .IN2(n7130), .Q(n7221) );
  AND2X1 U7969 ( .IN1(n7222), .IN2(n7132), .Q(n7206) );
  MUX21X1 U7970 ( .IN1(\mem0[159][7] ), .IN2(n851), .S(n7223), .Q(n17835) );
  MUX21X1 U7971 ( .IN1(\mem0[159][6] ), .IN2(n829), .S(n7223), .Q(n17834) );
  MUX21X1 U7972 ( .IN1(\mem0[159][5] ), .IN2(n807), .S(n7223), .Q(n17833) );
  MUX21X1 U7973 ( .IN1(\mem0[159][4] ), .IN2(n785), .S(n7223), .Q(n17832) );
  MUX21X1 U7974 ( .IN1(\mem0[159][3] ), .IN2(n763), .S(n7223), .Q(n17831) );
  MUX21X1 U7975 ( .IN1(\mem0[159][2] ), .IN2(n741), .S(n7223), .Q(n17830) );
  MUX21X1 U7976 ( .IN1(\mem0[159][1] ), .IN2(n719), .S(n7223), .Q(n17829) );
  MUX21X1 U7977 ( .IN1(\mem0[159][0] ), .IN2(n697), .S(n7223), .Q(n17828) );
  AND2X1 U7978 ( .IN1(n7224), .IN2(n7099), .Q(n7223) );
  MUX21X1 U7979 ( .IN1(\mem0[158][7] ), .IN2(n851), .S(n7225), .Q(n17827) );
  MUX21X1 U7980 ( .IN1(\mem0[158][6] ), .IN2(n829), .S(n7225), .Q(n17826) );
  MUX21X1 U7981 ( .IN1(\mem0[158][5] ), .IN2(n807), .S(n7225), .Q(n17825) );
  MUX21X1 U7982 ( .IN1(\mem0[158][4] ), .IN2(n785), .S(n7225), .Q(n17824) );
  MUX21X1 U7983 ( .IN1(\mem0[158][3] ), .IN2(n763), .S(n7225), .Q(n17823) );
  MUX21X1 U7984 ( .IN1(\mem0[158][2] ), .IN2(n741), .S(n7225), .Q(n17822) );
  MUX21X1 U7985 ( .IN1(\mem0[158][1] ), .IN2(n719), .S(n7225), .Q(n17821) );
  MUX21X1 U7986 ( .IN1(\mem0[158][0] ), .IN2(n697), .S(n7225), .Q(n17820) );
  AND2X1 U7987 ( .IN1(n7224), .IN2(n7102), .Q(n7225) );
  MUX21X1 U7988 ( .IN1(\mem0[157][7] ), .IN2(n851), .S(n7226), .Q(n17819) );
  MUX21X1 U7989 ( .IN1(\mem0[157][6] ), .IN2(n829), .S(n7226), .Q(n17818) );
  MUX21X1 U7990 ( .IN1(\mem0[157][5] ), .IN2(n807), .S(n7226), .Q(n17817) );
  MUX21X1 U7991 ( .IN1(\mem0[157][4] ), .IN2(n785), .S(n7226), .Q(n17816) );
  MUX21X1 U7992 ( .IN1(\mem0[157][3] ), .IN2(n763), .S(n7226), .Q(n17815) );
  MUX21X1 U7993 ( .IN1(\mem0[157][2] ), .IN2(n741), .S(n7226), .Q(n17814) );
  MUX21X1 U7994 ( .IN1(\mem0[157][1] ), .IN2(n719), .S(n7226), .Q(n17813) );
  MUX21X1 U7995 ( .IN1(\mem0[157][0] ), .IN2(n697), .S(n7226), .Q(n17812) );
  AND2X1 U7996 ( .IN1(n7224), .IN2(n7104), .Q(n7226) );
  MUX21X1 U7997 ( .IN1(\mem0[156][7] ), .IN2(n851), .S(n7227), .Q(n17811) );
  MUX21X1 U7998 ( .IN1(\mem0[156][6] ), .IN2(n829), .S(n7227), .Q(n17810) );
  MUX21X1 U7999 ( .IN1(\mem0[156][5] ), .IN2(n807), .S(n7227), .Q(n17809) );
  MUX21X1 U8000 ( .IN1(\mem0[156][4] ), .IN2(n785), .S(n7227), .Q(n17808) );
  MUX21X1 U8001 ( .IN1(\mem0[156][3] ), .IN2(n763), .S(n7227), .Q(n17807) );
  MUX21X1 U8002 ( .IN1(\mem0[156][2] ), .IN2(n741), .S(n7227), .Q(n17806) );
  MUX21X1 U8003 ( .IN1(\mem0[156][1] ), .IN2(n719), .S(n7227), .Q(n17805) );
  MUX21X1 U8004 ( .IN1(\mem0[156][0] ), .IN2(n697), .S(n7227), .Q(n17804) );
  AND2X1 U8005 ( .IN1(n7224), .IN2(n7106), .Q(n7227) );
  MUX21X1 U8006 ( .IN1(\mem0[155][7] ), .IN2(n851), .S(n7228), .Q(n17803) );
  MUX21X1 U8007 ( .IN1(\mem0[155][6] ), .IN2(n829), .S(n7228), .Q(n17802) );
  MUX21X1 U8008 ( .IN1(\mem0[155][5] ), .IN2(n807), .S(n7228), .Q(n17801) );
  MUX21X1 U8009 ( .IN1(\mem0[155][4] ), .IN2(n785), .S(n7228), .Q(n17800) );
  MUX21X1 U8010 ( .IN1(\mem0[155][3] ), .IN2(n763), .S(n7228), .Q(n17799) );
  MUX21X1 U8011 ( .IN1(\mem0[155][2] ), .IN2(n741), .S(n7228), .Q(n17798) );
  MUX21X1 U8012 ( .IN1(\mem0[155][1] ), .IN2(n719), .S(n7228), .Q(n17797) );
  MUX21X1 U8013 ( .IN1(\mem0[155][0] ), .IN2(n697), .S(n7228), .Q(n17796) );
  AND2X1 U8014 ( .IN1(n7224), .IN2(n7108), .Q(n7228) );
  MUX21X1 U8015 ( .IN1(\mem0[154][7] ), .IN2(n851), .S(n7229), .Q(n17795) );
  MUX21X1 U8016 ( .IN1(\mem0[154][6] ), .IN2(n829), .S(n7229), .Q(n17794) );
  MUX21X1 U8017 ( .IN1(\mem0[154][5] ), .IN2(n807), .S(n7229), .Q(n17793) );
  MUX21X1 U8018 ( .IN1(\mem0[154][4] ), .IN2(n785), .S(n7229), .Q(n17792) );
  MUX21X1 U8019 ( .IN1(\mem0[154][3] ), .IN2(n763), .S(n7229), .Q(n17791) );
  MUX21X1 U8020 ( .IN1(\mem0[154][2] ), .IN2(n741), .S(n7229), .Q(n17790) );
  MUX21X1 U8021 ( .IN1(\mem0[154][1] ), .IN2(n719), .S(n7229), .Q(n17789) );
  MUX21X1 U8022 ( .IN1(\mem0[154][0] ), .IN2(n697), .S(n7229), .Q(n17788) );
  AND2X1 U8023 ( .IN1(n7224), .IN2(n7110), .Q(n7229) );
  MUX21X1 U8024 ( .IN1(\mem0[153][7] ), .IN2(n851), .S(n7230), .Q(n17787) );
  MUX21X1 U8025 ( .IN1(\mem0[153][6] ), .IN2(n829), .S(n7230), .Q(n17786) );
  MUX21X1 U8026 ( .IN1(\mem0[153][5] ), .IN2(n807), .S(n7230), .Q(n17785) );
  MUX21X1 U8027 ( .IN1(\mem0[153][4] ), .IN2(n785), .S(n7230), .Q(n17784) );
  MUX21X1 U8028 ( .IN1(\mem0[153][3] ), .IN2(n763), .S(n7230), .Q(n17783) );
  MUX21X1 U8029 ( .IN1(\mem0[153][2] ), .IN2(n741), .S(n7230), .Q(n17782) );
  MUX21X1 U8030 ( .IN1(\mem0[153][1] ), .IN2(n719), .S(n7230), .Q(n17781) );
  MUX21X1 U8031 ( .IN1(\mem0[153][0] ), .IN2(n697), .S(n7230), .Q(n17780) );
  AND2X1 U8032 ( .IN1(n7224), .IN2(n7112), .Q(n7230) );
  MUX21X1 U8033 ( .IN1(\mem0[152][7] ), .IN2(n851), .S(n7231), .Q(n17779) );
  MUX21X1 U8034 ( .IN1(\mem0[152][6] ), .IN2(n829), .S(n7231), .Q(n17778) );
  MUX21X1 U8035 ( .IN1(\mem0[152][5] ), .IN2(n807), .S(n7231), .Q(n17777) );
  MUX21X1 U8036 ( .IN1(\mem0[152][4] ), .IN2(n785), .S(n7231), .Q(n17776) );
  MUX21X1 U8037 ( .IN1(\mem0[152][3] ), .IN2(n763), .S(n7231), .Q(n17775) );
  MUX21X1 U8038 ( .IN1(\mem0[152][2] ), .IN2(n741), .S(n7231), .Q(n17774) );
  MUX21X1 U8039 ( .IN1(\mem0[152][1] ), .IN2(n719), .S(n7231), .Q(n17773) );
  MUX21X1 U8040 ( .IN1(\mem0[152][0] ), .IN2(n697), .S(n7231), .Q(n17772) );
  AND2X1 U8041 ( .IN1(n7224), .IN2(n7114), .Q(n7231) );
  MUX21X1 U8042 ( .IN1(\mem0[151][7] ), .IN2(n851), .S(n7232), .Q(n17771) );
  MUX21X1 U8043 ( .IN1(\mem0[151][6] ), .IN2(n829), .S(n7232), .Q(n17770) );
  MUX21X1 U8044 ( .IN1(\mem0[151][5] ), .IN2(n807), .S(n7232), .Q(n17769) );
  MUX21X1 U8045 ( .IN1(\mem0[151][4] ), .IN2(n785), .S(n7232), .Q(n17768) );
  MUX21X1 U8046 ( .IN1(\mem0[151][3] ), .IN2(n763), .S(n7232), .Q(n17767) );
  MUX21X1 U8047 ( .IN1(\mem0[151][2] ), .IN2(n741), .S(n7232), .Q(n17766) );
  MUX21X1 U8048 ( .IN1(\mem0[151][1] ), .IN2(n719), .S(n7232), .Q(n17765) );
  MUX21X1 U8049 ( .IN1(\mem0[151][0] ), .IN2(n697), .S(n7232), .Q(n17764) );
  AND2X1 U8050 ( .IN1(n7224), .IN2(n7116), .Q(n7232) );
  MUX21X1 U8051 ( .IN1(\mem0[150][7] ), .IN2(n851), .S(n7233), .Q(n17763) );
  MUX21X1 U8052 ( .IN1(\mem0[150][6] ), .IN2(n829), .S(n7233), .Q(n17762) );
  MUX21X1 U8053 ( .IN1(\mem0[150][5] ), .IN2(n807), .S(n7233), .Q(n17761) );
  MUX21X1 U8054 ( .IN1(\mem0[150][4] ), .IN2(n785), .S(n7233), .Q(n17760) );
  MUX21X1 U8055 ( .IN1(\mem0[150][3] ), .IN2(n763), .S(n7233), .Q(n17759) );
  MUX21X1 U8056 ( .IN1(\mem0[150][2] ), .IN2(n741), .S(n7233), .Q(n17758) );
  MUX21X1 U8057 ( .IN1(\mem0[150][1] ), .IN2(n719), .S(n7233), .Q(n17757) );
  MUX21X1 U8058 ( .IN1(\mem0[150][0] ), .IN2(n697), .S(n7233), .Q(n17756) );
  AND2X1 U8059 ( .IN1(n7224), .IN2(n7118), .Q(n7233) );
  MUX21X1 U8060 ( .IN1(\mem0[149][7] ), .IN2(n851), .S(n7234), .Q(n17755) );
  MUX21X1 U8061 ( .IN1(\mem0[149][6] ), .IN2(n829), .S(n7234), .Q(n17754) );
  MUX21X1 U8062 ( .IN1(\mem0[149][5] ), .IN2(n807), .S(n7234), .Q(n17753) );
  MUX21X1 U8063 ( .IN1(\mem0[149][4] ), .IN2(n785), .S(n7234), .Q(n17752) );
  MUX21X1 U8064 ( .IN1(\mem0[149][3] ), .IN2(n763), .S(n7234), .Q(n17751) );
  MUX21X1 U8065 ( .IN1(\mem0[149][2] ), .IN2(n741), .S(n7234), .Q(n17750) );
  MUX21X1 U8066 ( .IN1(\mem0[149][1] ), .IN2(n719), .S(n7234), .Q(n17749) );
  MUX21X1 U8067 ( .IN1(\mem0[149][0] ), .IN2(n697), .S(n7234), .Q(n17748) );
  AND2X1 U8068 ( .IN1(n7224), .IN2(n7120), .Q(n7234) );
  MUX21X1 U8069 ( .IN1(\mem0[148][7] ), .IN2(n851), .S(n7235), .Q(n17747) );
  MUX21X1 U8070 ( .IN1(\mem0[148][6] ), .IN2(n829), .S(n7235), .Q(n17746) );
  MUX21X1 U8071 ( .IN1(\mem0[148][5] ), .IN2(n807), .S(n7235), .Q(n17745) );
  MUX21X1 U8072 ( .IN1(\mem0[148][4] ), .IN2(n785), .S(n7235), .Q(n17744) );
  MUX21X1 U8073 ( .IN1(\mem0[148][3] ), .IN2(n763), .S(n7235), .Q(n17743) );
  MUX21X1 U8074 ( .IN1(\mem0[148][2] ), .IN2(n741), .S(n7235), .Q(n17742) );
  MUX21X1 U8075 ( .IN1(\mem0[148][1] ), .IN2(n719), .S(n7235), .Q(n17741) );
  MUX21X1 U8076 ( .IN1(\mem0[148][0] ), .IN2(n697), .S(n7235), .Q(n17740) );
  AND2X1 U8077 ( .IN1(n7224), .IN2(n7122), .Q(n7235) );
  MUX21X1 U8078 ( .IN1(\mem0[147][7] ), .IN2(n852), .S(n7236), .Q(n17739) );
  MUX21X1 U8079 ( .IN1(\mem0[147][6] ), .IN2(n830), .S(n7236), .Q(n17738) );
  MUX21X1 U8080 ( .IN1(\mem0[147][5] ), .IN2(n808), .S(n7236), .Q(n17737) );
  MUX21X1 U8081 ( .IN1(\mem0[147][4] ), .IN2(n786), .S(n7236), .Q(n17736) );
  MUX21X1 U8082 ( .IN1(\mem0[147][3] ), .IN2(n764), .S(n7236), .Q(n17735) );
  MUX21X1 U8083 ( .IN1(\mem0[147][2] ), .IN2(n742), .S(n7236), .Q(n17734) );
  MUX21X1 U8084 ( .IN1(\mem0[147][1] ), .IN2(n720), .S(n7236), .Q(n17733) );
  MUX21X1 U8085 ( .IN1(\mem0[147][0] ), .IN2(n698), .S(n7236), .Q(n17732) );
  AND2X1 U8086 ( .IN1(n7224), .IN2(n7124), .Q(n7236) );
  MUX21X1 U8087 ( .IN1(\mem0[146][7] ), .IN2(n852), .S(n7237), .Q(n17731) );
  MUX21X1 U8088 ( .IN1(\mem0[146][6] ), .IN2(n830), .S(n7237), .Q(n17730) );
  MUX21X1 U8089 ( .IN1(\mem0[146][5] ), .IN2(n808), .S(n7237), .Q(n17729) );
  MUX21X1 U8090 ( .IN1(\mem0[146][4] ), .IN2(n786), .S(n7237), .Q(n17728) );
  MUX21X1 U8091 ( .IN1(\mem0[146][3] ), .IN2(n764), .S(n7237), .Q(n17727) );
  MUX21X1 U8092 ( .IN1(\mem0[146][2] ), .IN2(n742), .S(n7237), .Q(n17726) );
  MUX21X1 U8093 ( .IN1(\mem0[146][1] ), .IN2(n720), .S(n7237), .Q(n17725) );
  MUX21X1 U8094 ( .IN1(\mem0[146][0] ), .IN2(n698), .S(n7237), .Q(n17724) );
  AND2X1 U8095 ( .IN1(n7224), .IN2(n7126), .Q(n7237) );
  MUX21X1 U8096 ( .IN1(\mem0[145][7] ), .IN2(n852), .S(n7238), .Q(n17723) );
  MUX21X1 U8097 ( .IN1(\mem0[145][6] ), .IN2(n830), .S(n7238), .Q(n17722) );
  MUX21X1 U8098 ( .IN1(\mem0[145][5] ), .IN2(n808), .S(n7238), .Q(n17721) );
  MUX21X1 U8099 ( .IN1(\mem0[145][4] ), .IN2(n786), .S(n7238), .Q(n17720) );
  MUX21X1 U8100 ( .IN1(\mem0[145][3] ), .IN2(n764), .S(n7238), .Q(n17719) );
  MUX21X1 U8101 ( .IN1(\mem0[145][2] ), .IN2(n742), .S(n7238), .Q(n17718) );
  MUX21X1 U8102 ( .IN1(\mem0[145][1] ), .IN2(n720), .S(n7238), .Q(n17717) );
  MUX21X1 U8103 ( .IN1(\mem0[145][0] ), .IN2(n698), .S(n7238), .Q(n17716) );
  AND2X1 U8104 ( .IN1(n7224), .IN2(n7128), .Q(n7238) );
  MUX21X1 U8105 ( .IN1(\mem0[144][7] ), .IN2(n852), .S(n7239), .Q(n17715) );
  MUX21X1 U8106 ( .IN1(\mem0[144][6] ), .IN2(n830), .S(n7239), .Q(n17714) );
  MUX21X1 U8107 ( .IN1(\mem0[144][5] ), .IN2(n808), .S(n7239), .Q(n17713) );
  MUX21X1 U8108 ( .IN1(\mem0[144][4] ), .IN2(n786), .S(n7239), .Q(n17712) );
  MUX21X1 U8109 ( .IN1(\mem0[144][3] ), .IN2(n764), .S(n7239), .Q(n17711) );
  MUX21X1 U8110 ( .IN1(\mem0[144][2] ), .IN2(n742), .S(n7239), .Q(n17710) );
  MUX21X1 U8111 ( .IN1(\mem0[144][1] ), .IN2(n720), .S(n7239), .Q(n17709) );
  MUX21X1 U8112 ( .IN1(\mem0[144][0] ), .IN2(n698), .S(n7239), .Q(n17708) );
  AND2X1 U8113 ( .IN1(n7224), .IN2(n7130), .Q(n7239) );
  AND2X1 U8114 ( .IN1(n7240), .IN2(n7132), .Q(n7224) );
  MUX21X1 U8115 ( .IN1(\mem0[143][7] ), .IN2(n852), .S(n7241), .Q(n17707) );
  MUX21X1 U8116 ( .IN1(\mem0[143][6] ), .IN2(n830), .S(n7241), .Q(n17706) );
  MUX21X1 U8117 ( .IN1(\mem0[143][5] ), .IN2(n808), .S(n7241), .Q(n17705) );
  MUX21X1 U8118 ( .IN1(\mem0[143][4] ), .IN2(n786), .S(n7241), .Q(n17704) );
  MUX21X1 U8119 ( .IN1(\mem0[143][3] ), .IN2(n764), .S(n7241), .Q(n17703) );
  MUX21X1 U8120 ( .IN1(\mem0[143][2] ), .IN2(n742), .S(n7241), .Q(n17702) );
  MUX21X1 U8121 ( .IN1(\mem0[143][1] ), .IN2(n720), .S(n7241), .Q(n17701) );
  MUX21X1 U8122 ( .IN1(\mem0[143][0] ), .IN2(n698), .S(n7241), .Q(n17700) );
  AND2X1 U8123 ( .IN1(n7242), .IN2(n7099), .Q(n7241) );
  MUX21X1 U8124 ( .IN1(\mem0[142][7] ), .IN2(n852), .S(n7243), .Q(n17699) );
  MUX21X1 U8125 ( .IN1(\mem0[142][6] ), .IN2(n830), .S(n7243), .Q(n17698) );
  MUX21X1 U8126 ( .IN1(\mem0[142][5] ), .IN2(n808), .S(n7243), .Q(n17697) );
  MUX21X1 U8127 ( .IN1(\mem0[142][4] ), .IN2(n786), .S(n7243), .Q(n17696) );
  MUX21X1 U8128 ( .IN1(\mem0[142][3] ), .IN2(n764), .S(n7243), .Q(n17695) );
  MUX21X1 U8129 ( .IN1(\mem0[142][2] ), .IN2(n742), .S(n7243), .Q(n17694) );
  MUX21X1 U8130 ( .IN1(\mem0[142][1] ), .IN2(n720), .S(n7243), .Q(n17693) );
  MUX21X1 U8131 ( .IN1(\mem0[142][0] ), .IN2(n698), .S(n7243), .Q(n17692) );
  AND2X1 U8132 ( .IN1(n7242), .IN2(n7102), .Q(n7243) );
  MUX21X1 U8133 ( .IN1(\mem0[141][7] ), .IN2(n852), .S(n7244), .Q(n17691) );
  MUX21X1 U8134 ( .IN1(\mem0[141][6] ), .IN2(n830), .S(n7244), .Q(n17690) );
  MUX21X1 U8135 ( .IN1(\mem0[141][5] ), .IN2(n808), .S(n7244), .Q(n17689) );
  MUX21X1 U8136 ( .IN1(\mem0[141][4] ), .IN2(n786), .S(n7244), .Q(n17688) );
  MUX21X1 U8137 ( .IN1(\mem0[141][3] ), .IN2(n764), .S(n7244), .Q(n17687) );
  MUX21X1 U8138 ( .IN1(\mem0[141][2] ), .IN2(n742), .S(n7244), .Q(n17686) );
  MUX21X1 U8139 ( .IN1(\mem0[141][1] ), .IN2(n720), .S(n7244), .Q(n17685) );
  MUX21X1 U8140 ( .IN1(\mem0[141][0] ), .IN2(n698), .S(n7244), .Q(n17684) );
  AND2X1 U8141 ( .IN1(n7242), .IN2(n7104), .Q(n7244) );
  MUX21X1 U8142 ( .IN1(\mem0[140][7] ), .IN2(n852), .S(n7245), .Q(n17683) );
  MUX21X1 U8143 ( .IN1(\mem0[140][6] ), .IN2(n830), .S(n7245), .Q(n17682) );
  MUX21X1 U8144 ( .IN1(\mem0[140][5] ), .IN2(n808), .S(n7245), .Q(n17681) );
  MUX21X1 U8145 ( .IN1(\mem0[140][4] ), .IN2(n786), .S(n7245), .Q(n17680) );
  MUX21X1 U8146 ( .IN1(\mem0[140][3] ), .IN2(n764), .S(n7245), .Q(n17679) );
  MUX21X1 U8147 ( .IN1(\mem0[140][2] ), .IN2(n742), .S(n7245), .Q(n17678) );
  MUX21X1 U8148 ( .IN1(\mem0[140][1] ), .IN2(n720), .S(n7245), .Q(n17677) );
  MUX21X1 U8149 ( .IN1(\mem0[140][0] ), .IN2(n698), .S(n7245), .Q(n17676) );
  AND2X1 U8150 ( .IN1(n7242), .IN2(n7106), .Q(n7245) );
  MUX21X1 U8151 ( .IN1(\mem0[139][7] ), .IN2(n852), .S(n7246), .Q(n17675) );
  MUX21X1 U8152 ( .IN1(\mem0[139][6] ), .IN2(n830), .S(n7246), .Q(n17674) );
  MUX21X1 U8153 ( .IN1(\mem0[139][5] ), .IN2(n808), .S(n7246), .Q(n17673) );
  MUX21X1 U8154 ( .IN1(\mem0[139][4] ), .IN2(n786), .S(n7246), .Q(n17672) );
  MUX21X1 U8155 ( .IN1(\mem0[139][3] ), .IN2(n764), .S(n7246), .Q(n17671) );
  MUX21X1 U8156 ( .IN1(\mem0[139][2] ), .IN2(n742), .S(n7246), .Q(n17670) );
  MUX21X1 U8157 ( .IN1(\mem0[139][1] ), .IN2(n720), .S(n7246), .Q(n17669) );
  MUX21X1 U8158 ( .IN1(\mem0[139][0] ), .IN2(n698), .S(n7246), .Q(n17668) );
  AND2X1 U8159 ( .IN1(n7242), .IN2(n7108), .Q(n7246) );
  MUX21X1 U8160 ( .IN1(\mem0[138][7] ), .IN2(n852), .S(n7247), .Q(n17667) );
  MUX21X1 U8161 ( .IN1(\mem0[138][6] ), .IN2(n830), .S(n7247), .Q(n17666) );
  MUX21X1 U8162 ( .IN1(\mem0[138][5] ), .IN2(n808), .S(n7247), .Q(n17665) );
  MUX21X1 U8163 ( .IN1(\mem0[138][4] ), .IN2(n786), .S(n7247), .Q(n17664) );
  MUX21X1 U8164 ( .IN1(\mem0[138][3] ), .IN2(n764), .S(n7247), .Q(n17663) );
  MUX21X1 U8165 ( .IN1(\mem0[138][2] ), .IN2(n742), .S(n7247), .Q(n17662) );
  MUX21X1 U8166 ( .IN1(\mem0[138][1] ), .IN2(n720), .S(n7247), .Q(n17661) );
  MUX21X1 U8167 ( .IN1(\mem0[138][0] ), .IN2(n698), .S(n7247), .Q(n17660) );
  AND2X1 U8168 ( .IN1(n7242), .IN2(n7110), .Q(n7247) );
  MUX21X1 U8169 ( .IN1(\mem0[137][7] ), .IN2(n852), .S(n7248), .Q(n17659) );
  MUX21X1 U8170 ( .IN1(\mem0[137][6] ), .IN2(n830), .S(n7248), .Q(n17658) );
  MUX21X1 U8171 ( .IN1(\mem0[137][5] ), .IN2(n808), .S(n7248), .Q(n17657) );
  MUX21X1 U8172 ( .IN1(\mem0[137][4] ), .IN2(n786), .S(n7248), .Q(n17656) );
  MUX21X1 U8173 ( .IN1(\mem0[137][3] ), .IN2(n764), .S(n7248), .Q(n17655) );
  MUX21X1 U8174 ( .IN1(\mem0[137][2] ), .IN2(n742), .S(n7248), .Q(n17654) );
  MUX21X1 U8175 ( .IN1(\mem0[137][1] ), .IN2(n720), .S(n7248), .Q(n17653) );
  MUX21X1 U8176 ( .IN1(\mem0[137][0] ), .IN2(n698), .S(n7248), .Q(n17652) );
  AND2X1 U8177 ( .IN1(n7242), .IN2(n7112), .Q(n7248) );
  MUX21X1 U8178 ( .IN1(\mem0[136][7] ), .IN2(n852), .S(n7249), .Q(n17651) );
  MUX21X1 U8179 ( .IN1(\mem0[136][6] ), .IN2(n830), .S(n7249), .Q(n17650) );
  MUX21X1 U8180 ( .IN1(\mem0[136][5] ), .IN2(n808), .S(n7249), .Q(n17649) );
  MUX21X1 U8181 ( .IN1(\mem0[136][4] ), .IN2(n786), .S(n7249), .Q(n17648) );
  MUX21X1 U8182 ( .IN1(\mem0[136][3] ), .IN2(n764), .S(n7249), .Q(n17647) );
  MUX21X1 U8183 ( .IN1(\mem0[136][2] ), .IN2(n742), .S(n7249), .Q(n17646) );
  MUX21X1 U8184 ( .IN1(\mem0[136][1] ), .IN2(n720), .S(n7249), .Q(n17645) );
  MUX21X1 U8185 ( .IN1(\mem0[136][0] ), .IN2(n698), .S(n7249), .Q(n17644) );
  AND2X1 U8186 ( .IN1(n7242), .IN2(n7114), .Q(n7249) );
  MUX21X1 U8187 ( .IN1(\mem0[135][7] ), .IN2(n853), .S(n7250), .Q(n17643) );
  MUX21X1 U8188 ( .IN1(\mem0[135][6] ), .IN2(n831), .S(n7250), .Q(n17642) );
  MUX21X1 U8189 ( .IN1(\mem0[135][5] ), .IN2(n809), .S(n7250), .Q(n17641) );
  MUX21X1 U8190 ( .IN1(\mem0[135][4] ), .IN2(n787), .S(n7250), .Q(n17640) );
  MUX21X1 U8191 ( .IN1(\mem0[135][3] ), .IN2(n765), .S(n7250), .Q(n17639) );
  MUX21X1 U8192 ( .IN1(\mem0[135][2] ), .IN2(n743), .S(n7250), .Q(n17638) );
  MUX21X1 U8193 ( .IN1(\mem0[135][1] ), .IN2(n721), .S(n7250), .Q(n17637) );
  MUX21X1 U8194 ( .IN1(\mem0[135][0] ), .IN2(n699), .S(n7250), .Q(n17636) );
  AND2X1 U8195 ( .IN1(n7242), .IN2(n7116), .Q(n7250) );
  MUX21X1 U8196 ( .IN1(\mem0[134][7] ), .IN2(n853), .S(n7251), .Q(n17635) );
  MUX21X1 U8197 ( .IN1(\mem0[134][6] ), .IN2(n831), .S(n7251), .Q(n17634) );
  MUX21X1 U8198 ( .IN1(\mem0[134][5] ), .IN2(n809), .S(n7251), .Q(n17633) );
  MUX21X1 U8199 ( .IN1(\mem0[134][4] ), .IN2(n787), .S(n7251), .Q(n17632) );
  MUX21X1 U8200 ( .IN1(\mem0[134][3] ), .IN2(n765), .S(n7251), .Q(n17631) );
  MUX21X1 U8201 ( .IN1(\mem0[134][2] ), .IN2(n743), .S(n7251), .Q(n17630) );
  MUX21X1 U8202 ( .IN1(\mem0[134][1] ), .IN2(n721), .S(n7251), .Q(n17629) );
  MUX21X1 U8203 ( .IN1(\mem0[134][0] ), .IN2(n699), .S(n7251), .Q(n17628) );
  AND2X1 U8204 ( .IN1(n7242), .IN2(n7118), .Q(n7251) );
  MUX21X1 U8205 ( .IN1(\mem0[133][7] ), .IN2(n853), .S(n7252), .Q(n17627) );
  MUX21X1 U8206 ( .IN1(\mem0[133][6] ), .IN2(n831), .S(n7252), .Q(n17626) );
  MUX21X1 U8207 ( .IN1(\mem0[133][5] ), .IN2(n809), .S(n7252), .Q(n17625) );
  MUX21X1 U8208 ( .IN1(\mem0[133][4] ), .IN2(n787), .S(n7252), .Q(n17624) );
  MUX21X1 U8209 ( .IN1(\mem0[133][3] ), .IN2(n765), .S(n7252), .Q(n17623) );
  MUX21X1 U8210 ( .IN1(\mem0[133][2] ), .IN2(n743), .S(n7252), .Q(n17622) );
  MUX21X1 U8211 ( .IN1(\mem0[133][1] ), .IN2(n721), .S(n7252), .Q(n17621) );
  MUX21X1 U8212 ( .IN1(\mem0[133][0] ), .IN2(n699), .S(n7252), .Q(n17620) );
  AND2X1 U8213 ( .IN1(n7242), .IN2(n7120), .Q(n7252) );
  MUX21X1 U8214 ( .IN1(\mem0[132][7] ), .IN2(n853), .S(n7253), .Q(n17619) );
  MUX21X1 U8215 ( .IN1(\mem0[132][6] ), .IN2(n831), .S(n7253), .Q(n17618) );
  MUX21X1 U8216 ( .IN1(\mem0[132][5] ), .IN2(n809), .S(n7253), .Q(n17617) );
  MUX21X1 U8217 ( .IN1(\mem0[132][4] ), .IN2(n787), .S(n7253), .Q(n17616) );
  MUX21X1 U8218 ( .IN1(\mem0[132][3] ), .IN2(n765), .S(n7253), .Q(n17615) );
  MUX21X1 U8219 ( .IN1(\mem0[132][2] ), .IN2(n743), .S(n7253), .Q(n17614) );
  MUX21X1 U8220 ( .IN1(\mem0[132][1] ), .IN2(n721), .S(n7253), .Q(n17613) );
  MUX21X1 U8221 ( .IN1(\mem0[132][0] ), .IN2(n699), .S(n7253), .Q(n17612) );
  AND2X1 U8222 ( .IN1(n7242), .IN2(n7122), .Q(n7253) );
  MUX21X1 U8223 ( .IN1(\mem0[131][7] ), .IN2(n853), .S(n7254), .Q(n17611) );
  MUX21X1 U8224 ( .IN1(\mem0[131][6] ), .IN2(n831), .S(n7254), .Q(n17610) );
  MUX21X1 U8225 ( .IN1(\mem0[131][5] ), .IN2(n809), .S(n7254), .Q(n17609) );
  MUX21X1 U8226 ( .IN1(\mem0[131][4] ), .IN2(n787), .S(n7254), .Q(n17608) );
  MUX21X1 U8227 ( .IN1(\mem0[131][3] ), .IN2(n765), .S(n7254), .Q(n17607) );
  MUX21X1 U8228 ( .IN1(\mem0[131][2] ), .IN2(n743), .S(n7254), .Q(n17606) );
  MUX21X1 U8229 ( .IN1(\mem0[131][1] ), .IN2(n721), .S(n7254), .Q(n17605) );
  MUX21X1 U8230 ( .IN1(\mem0[131][0] ), .IN2(n699), .S(n7254), .Q(n17604) );
  AND2X1 U8231 ( .IN1(n7242), .IN2(n7124), .Q(n7254) );
  MUX21X1 U8232 ( .IN1(\mem0[130][7] ), .IN2(n853), .S(n7255), .Q(n17603) );
  MUX21X1 U8233 ( .IN1(\mem0[130][6] ), .IN2(n831), .S(n7255), .Q(n17602) );
  MUX21X1 U8234 ( .IN1(\mem0[130][5] ), .IN2(n809), .S(n7255), .Q(n17601) );
  MUX21X1 U8235 ( .IN1(\mem0[130][4] ), .IN2(n787), .S(n7255), .Q(n17600) );
  MUX21X1 U8236 ( .IN1(\mem0[130][3] ), .IN2(n765), .S(n7255), .Q(n17599) );
  MUX21X1 U8237 ( .IN1(\mem0[130][2] ), .IN2(n743), .S(n7255), .Q(n17598) );
  MUX21X1 U8238 ( .IN1(\mem0[130][1] ), .IN2(n721), .S(n7255), .Q(n17597) );
  MUX21X1 U8239 ( .IN1(\mem0[130][0] ), .IN2(n699), .S(n7255), .Q(n17596) );
  AND2X1 U8240 ( .IN1(n7242), .IN2(n7126), .Q(n7255) );
  MUX21X1 U8241 ( .IN1(\mem0[129][7] ), .IN2(n853), .S(n7256), .Q(n17595) );
  MUX21X1 U8242 ( .IN1(\mem0[129][6] ), .IN2(n831), .S(n7256), .Q(n17594) );
  MUX21X1 U8243 ( .IN1(\mem0[129][5] ), .IN2(n809), .S(n7256), .Q(n17593) );
  MUX21X1 U8244 ( .IN1(\mem0[129][4] ), .IN2(n787), .S(n7256), .Q(n17592) );
  MUX21X1 U8245 ( .IN1(\mem0[129][3] ), .IN2(n765), .S(n7256), .Q(n17591) );
  MUX21X1 U8246 ( .IN1(\mem0[129][2] ), .IN2(n743), .S(n7256), .Q(n17590) );
  MUX21X1 U8247 ( .IN1(\mem0[129][1] ), .IN2(n721), .S(n7256), .Q(n17589) );
  MUX21X1 U8248 ( .IN1(\mem0[129][0] ), .IN2(n699), .S(n7256), .Q(n17588) );
  AND2X1 U8249 ( .IN1(n7242), .IN2(n7128), .Q(n7256) );
  MUX21X1 U8250 ( .IN1(\mem0[128][7] ), .IN2(n853), .S(n7257), .Q(n17587) );
  MUX21X1 U8251 ( .IN1(\mem0[128][6] ), .IN2(n831), .S(n7257), .Q(n17586) );
  MUX21X1 U8252 ( .IN1(\mem0[128][5] ), .IN2(n809), .S(n7257), .Q(n17585) );
  MUX21X1 U8253 ( .IN1(\mem0[128][4] ), .IN2(n787), .S(n7257), .Q(n17584) );
  MUX21X1 U8254 ( .IN1(\mem0[128][3] ), .IN2(n765), .S(n7257), .Q(n17583) );
  MUX21X1 U8255 ( .IN1(\mem0[128][2] ), .IN2(n743), .S(n7257), .Q(n17582) );
  MUX21X1 U8256 ( .IN1(\mem0[128][1] ), .IN2(n721), .S(n7257), .Q(n17581) );
  MUX21X1 U8257 ( .IN1(\mem0[128][0] ), .IN2(n699), .S(n7257), .Q(n17580) );
  AND2X1 U8258 ( .IN1(n7242), .IN2(n7130), .Q(n7257) );
  AND2X1 U8259 ( .IN1(n7258), .IN2(n7132), .Q(n7242) );
  MUX21X1 U8260 ( .IN1(\mem0[127][7] ), .IN2(n853), .S(n7259), .Q(n17579) );
  MUX21X1 U8261 ( .IN1(\mem0[127][6] ), .IN2(n831), .S(n7259), .Q(n17578) );
  MUX21X1 U8262 ( .IN1(\mem0[127][5] ), .IN2(n809), .S(n7259), .Q(n17577) );
  MUX21X1 U8263 ( .IN1(\mem0[127][4] ), .IN2(n787), .S(n7259), .Q(n17576) );
  MUX21X1 U8264 ( .IN1(\mem0[127][3] ), .IN2(n765), .S(n7259), .Q(n17575) );
  MUX21X1 U8265 ( .IN1(\mem0[127][2] ), .IN2(n743), .S(n7259), .Q(n17574) );
  MUX21X1 U8266 ( .IN1(\mem0[127][1] ), .IN2(n721), .S(n7259), .Q(n17573) );
  MUX21X1 U8267 ( .IN1(\mem0[127][0] ), .IN2(n699), .S(n7259), .Q(n17572) );
  AND2X1 U8268 ( .IN1(n7260), .IN2(n7099), .Q(n7259) );
  MUX21X1 U8269 ( .IN1(\mem0[126][7] ), .IN2(n853), .S(n7261), .Q(n17571) );
  MUX21X1 U8270 ( .IN1(\mem0[126][6] ), .IN2(n831), .S(n7261), .Q(n17570) );
  MUX21X1 U8271 ( .IN1(\mem0[126][5] ), .IN2(n809), .S(n7261), .Q(n17569) );
  MUX21X1 U8272 ( .IN1(\mem0[126][4] ), .IN2(n787), .S(n7261), .Q(n17568) );
  MUX21X1 U8273 ( .IN1(\mem0[126][3] ), .IN2(n765), .S(n7261), .Q(n17567) );
  MUX21X1 U8274 ( .IN1(\mem0[126][2] ), .IN2(n743), .S(n7261), .Q(n17566) );
  MUX21X1 U8275 ( .IN1(\mem0[126][1] ), .IN2(n721), .S(n7261), .Q(n17565) );
  MUX21X1 U8276 ( .IN1(\mem0[126][0] ), .IN2(n699), .S(n7261), .Q(n17564) );
  AND2X1 U8277 ( .IN1(n7260), .IN2(n7102), .Q(n7261) );
  MUX21X1 U8278 ( .IN1(\mem0[125][7] ), .IN2(n853), .S(n7262), .Q(n17563) );
  MUX21X1 U8279 ( .IN1(\mem0[125][6] ), .IN2(n831), .S(n7262), .Q(n17562) );
  MUX21X1 U8280 ( .IN1(\mem0[125][5] ), .IN2(n809), .S(n7262), .Q(n17561) );
  MUX21X1 U8281 ( .IN1(\mem0[125][4] ), .IN2(n787), .S(n7262), .Q(n17560) );
  MUX21X1 U8282 ( .IN1(\mem0[125][3] ), .IN2(n765), .S(n7262), .Q(n17559) );
  MUX21X1 U8283 ( .IN1(\mem0[125][2] ), .IN2(n743), .S(n7262), .Q(n17558) );
  MUX21X1 U8284 ( .IN1(\mem0[125][1] ), .IN2(n721), .S(n7262), .Q(n17557) );
  MUX21X1 U8285 ( .IN1(\mem0[125][0] ), .IN2(n699), .S(n7262), .Q(n17556) );
  AND2X1 U8286 ( .IN1(n7260), .IN2(n7104), .Q(n7262) );
  MUX21X1 U8287 ( .IN1(\mem0[124][7] ), .IN2(n853), .S(n7263), .Q(n17555) );
  MUX21X1 U8288 ( .IN1(\mem0[124][6] ), .IN2(n831), .S(n7263), .Q(n17554) );
  MUX21X1 U8289 ( .IN1(\mem0[124][5] ), .IN2(n809), .S(n7263), .Q(n17553) );
  MUX21X1 U8290 ( .IN1(\mem0[124][4] ), .IN2(n787), .S(n7263), .Q(n17552) );
  MUX21X1 U8291 ( .IN1(\mem0[124][3] ), .IN2(n765), .S(n7263), .Q(n17551) );
  MUX21X1 U8292 ( .IN1(\mem0[124][2] ), .IN2(n743), .S(n7263), .Q(n17550) );
  MUX21X1 U8293 ( .IN1(\mem0[124][1] ), .IN2(n721), .S(n7263), .Q(n17549) );
  MUX21X1 U8294 ( .IN1(\mem0[124][0] ), .IN2(n699), .S(n7263), .Q(n17548) );
  AND2X1 U8295 ( .IN1(n7260), .IN2(n7106), .Q(n7263) );
  MUX21X1 U8296 ( .IN1(\mem0[123][7] ), .IN2(n854), .S(n7264), .Q(n17547) );
  MUX21X1 U8297 ( .IN1(\mem0[123][6] ), .IN2(n832), .S(n7264), .Q(n17546) );
  MUX21X1 U8298 ( .IN1(\mem0[123][5] ), .IN2(n810), .S(n7264), .Q(n17545) );
  MUX21X1 U8299 ( .IN1(\mem0[123][4] ), .IN2(n788), .S(n7264), .Q(n17544) );
  MUX21X1 U8300 ( .IN1(\mem0[123][3] ), .IN2(n766), .S(n7264), .Q(n17543) );
  MUX21X1 U8301 ( .IN1(\mem0[123][2] ), .IN2(n744), .S(n7264), .Q(n17542) );
  MUX21X1 U8302 ( .IN1(\mem0[123][1] ), .IN2(n722), .S(n7264), .Q(n17541) );
  MUX21X1 U8303 ( .IN1(\mem0[123][0] ), .IN2(n700), .S(n7264), .Q(n17540) );
  AND2X1 U8304 ( .IN1(n7260), .IN2(n7108), .Q(n7264) );
  MUX21X1 U8305 ( .IN1(\mem0[122][7] ), .IN2(n854), .S(n7265), .Q(n17539) );
  MUX21X1 U8306 ( .IN1(\mem0[122][6] ), .IN2(n832), .S(n7265), .Q(n17538) );
  MUX21X1 U8307 ( .IN1(\mem0[122][5] ), .IN2(n810), .S(n7265), .Q(n17537) );
  MUX21X1 U8308 ( .IN1(\mem0[122][4] ), .IN2(n788), .S(n7265), .Q(n17536) );
  MUX21X1 U8309 ( .IN1(\mem0[122][3] ), .IN2(n766), .S(n7265), .Q(n17535) );
  MUX21X1 U8310 ( .IN1(\mem0[122][2] ), .IN2(n744), .S(n7265), .Q(n17534) );
  MUX21X1 U8311 ( .IN1(\mem0[122][1] ), .IN2(n722), .S(n7265), .Q(n17533) );
  MUX21X1 U8312 ( .IN1(\mem0[122][0] ), .IN2(n700), .S(n7265), .Q(n17532) );
  AND2X1 U8313 ( .IN1(n7260), .IN2(n7110), .Q(n7265) );
  MUX21X1 U8314 ( .IN1(\mem0[121][7] ), .IN2(n854), .S(n7266), .Q(n17531) );
  MUX21X1 U8315 ( .IN1(\mem0[121][6] ), .IN2(n832), .S(n7266), .Q(n17530) );
  MUX21X1 U8316 ( .IN1(\mem0[121][5] ), .IN2(n810), .S(n7266), .Q(n17529) );
  MUX21X1 U8317 ( .IN1(\mem0[121][4] ), .IN2(n788), .S(n7266), .Q(n17528) );
  MUX21X1 U8318 ( .IN1(\mem0[121][3] ), .IN2(n766), .S(n7266), .Q(n17527) );
  MUX21X1 U8319 ( .IN1(\mem0[121][2] ), .IN2(n744), .S(n7266), .Q(n17526) );
  MUX21X1 U8320 ( .IN1(\mem0[121][1] ), .IN2(n722), .S(n7266), .Q(n17525) );
  MUX21X1 U8321 ( .IN1(\mem0[121][0] ), .IN2(n700), .S(n7266), .Q(n17524) );
  AND2X1 U8322 ( .IN1(n7260), .IN2(n7112), .Q(n7266) );
  MUX21X1 U8323 ( .IN1(\mem0[120][7] ), .IN2(n854), .S(n7267), .Q(n17523) );
  MUX21X1 U8324 ( .IN1(\mem0[120][6] ), .IN2(n832), .S(n7267), .Q(n17522) );
  MUX21X1 U8325 ( .IN1(\mem0[120][5] ), .IN2(n810), .S(n7267), .Q(n17521) );
  MUX21X1 U8326 ( .IN1(\mem0[120][4] ), .IN2(n788), .S(n7267), .Q(n17520) );
  MUX21X1 U8327 ( .IN1(\mem0[120][3] ), .IN2(n766), .S(n7267), .Q(n17519) );
  MUX21X1 U8328 ( .IN1(\mem0[120][2] ), .IN2(n744), .S(n7267), .Q(n17518) );
  MUX21X1 U8329 ( .IN1(\mem0[120][1] ), .IN2(n722), .S(n7267), .Q(n17517) );
  MUX21X1 U8330 ( .IN1(\mem0[120][0] ), .IN2(n700), .S(n7267), .Q(n17516) );
  AND2X1 U8331 ( .IN1(n7260), .IN2(n7114), .Q(n7267) );
  MUX21X1 U8332 ( .IN1(\mem0[119][7] ), .IN2(n854), .S(n7268), .Q(n17515) );
  MUX21X1 U8333 ( .IN1(\mem0[119][6] ), .IN2(n832), .S(n7268), .Q(n17514) );
  MUX21X1 U8334 ( .IN1(\mem0[119][5] ), .IN2(n810), .S(n7268), .Q(n17513) );
  MUX21X1 U8335 ( .IN1(\mem0[119][4] ), .IN2(n788), .S(n7268), .Q(n17512) );
  MUX21X1 U8336 ( .IN1(\mem0[119][3] ), .IN2(n766), .S(n7268), .Q(n17511) );
  MUX21X1 U8337 ( .IN1(\mem0[119][2] ), .IN2(n744), .S(n7268), .Q(n17510) );
  MUX21X1 U8338 ( .IN1(\mem0[119][1] ), .IN2(n722), .S(n7268), .Q(n17509) );
  MUX21X1 U8339 ( .IN1(\mem0[119][0] ), .IN2(n700), .S(n7268), .Q(n17508) );
  AND2X1 U8340 ( .IN1(n7260), .IN2(n7116), .Q(n7268) );
  MUX21X1 U8341 ( .IN1(\mem0[118][7] ), .IN2(n854), .S(n7269), .Q(n17507) );
  MUX21X1 U8342 ( .IN1(\mem0[118][6] ), .IN2(n832), .S(n7269), .Q(n17506) );
  MUX21X1 U8343 ( .IN1(\mem0[118][5] ), .IN2(n810), .S(n7269), .Q(n17505) );
  MUX21X1 U8344 ( .IN1(\mem0[118][4] ), .IN2(n788), .S(n7269), .Q(n17504) );
  MUX21X1 U8345 ( .IN1(\mem0[118][3] ), .IN2(n766), .S(n7269), .Q(n17503) );
  MUX21X1 U8346 ( .IN1(\mem0[118][2] ), .IN2(n744), .S(n7269), .Q(n17502) );
  MUX21X1 U8347 ( .IN1(\mem0[118][1] ), .IN2(n722), .S(n7269), .Q(n17501) );
  MUX21X1 U8348 ( .IN1(\mem0[118][0] ), .IN2(n700), .S(n7269), .Q(n17500) );
  AND2X1 U8349 ( .IN1(n7260), .IN2(n7118), .Q(n7269) );
  MUX21X1 U8350 ( .IN1(\mem0[117][7] ), .IN2(n854), .S(n7270), .Q(n17499) );
  MUX21X1 U8351 ( .IN1(\mem0[117][6] ), .IN2(n832), .S(n7270), .Q(n17498) );
  MUX21X1 U8352 ( .IN1(\mem0[117][5] ), .IN2(n810), .S(n7270), .Q(n17497) );
  MUX21X1 U8353 ( .IN1(\mem0[117][4] ), .IN2(n788), .S(n7270), .Q(n17496) );
  MUX21X1 U8354 ( .IN1(\mem0[117][3] ), .IN2(n766), .S(n7270), .Q(n17495) );
  MUX21X1 U8355 ( .IN1(\mem0[117][2] ), .IN2(n744), .S(n7270), .Q(n17494) );
  MUX21X1 U8356 ( .IN1(\mem0[117][1] ), .IN2(n722), .S(n7270), .Q(n17493) );
  MUX21X1 U8357 ( .IN1(\mem0[117][0] ), .IN2(n700), .S(n7270), .Q(n17492) );
  AND2X1 U8358 ( .IN1(n7260), .IN2(n7120), .Q(n7270) );
  MUX21X1 U8359 ( .IN1(\mem0[116][7] ), .IN2(n854), .S(n7271), .Q(n17491) );
  MUX21X1 U8360 ( .IN1(\mem0[116][6] ), .IN2(n832), .S(n7271), .Q(n17490) );
  MUX21X1 U8361 ( .IN1(\mem0[116][5] ), .IN2(n810), .S(n7271), .Q(n17489) );
  MUX21X1 U8362 ( .IN1(\mem0[116][4] ), .IN2(n788), .S(n7271), .Q(n17488) );
  MUX21X1 U8363 ( .IN1(\mem0[116][3] ), .IN2(n766), .S(n7271), .Q(n17487) );
  MUX21X1 U8364 ( .IN1(\mem0[116][2] ), .IN2(n744), .S(n7271), .Q(n17486) );
  MUX21X1 U8365 ( .IN1(\mem0[116][1] ), .IN2(n722), .S(n7271), .Q(n17485) );
  MUX21X1 U8366 ( .IN1(\mem0[116][0] ), .IN2(n700), .S(n7271), .Q(n17484) );
  AND2X1 U8367 ( .IN1(n7260), .IN2(n7122), .Q(n7271) );
  MUX21X1 U8368 ( .IN1(\mem0[115][7] ), .IN2(n854), .S(n7272), .Q(n17483) );
  MUX21X1 U8369 ( .IN1(\mem0[115][6] ), .IN2(n832), .S(n7272), .Q(n17482) );
  MUX21X1 U8370 ( .IN1(\mem0[115][5] ), .IN2(n810), .S(n7272), .Q(n17481) );
  MUX21X1 U8371 ( .IN1(\mem0[115][4] ), .IN2(n788), .S(n7272), .Q(n17480) );
  MUX21X1 U8372 ( .IN1(\mem0[115][3] ), .IN2(n766), .S(n7272), .Q(n17479) );
  MUX21X1 U8373 ( .IN1(\mem0[115][2] ), .IN2(n744), .S(n7272), .Q(n17478) );
  MUX21X1 U8374 ( .IN1(\mem0[115][1] ), .IN2(n722), .S(n7272), .Q(n17477) );
  MUX21X1 U8375 ( .IN1(\mem0[115][0] ), .IN2(n700), .S(n7272), .Q(n17476) );
  AND2X1 U8376 ( .IN1(n7260), .IN2(n7124), .Q(n7272) );
  MUX21X1 U8377 ( .IN1(\mem0[114][7] ), .IN2(n854), .S(n7273), .Q(n17475) );
  MUX21X1 U8378 ( .IN1(\mem0[114][6] ), .IN2(n832), .S(n7273), .Q(n17474) );
  MUX21X1 U8379 ( .IN1(\mem0[114][5] ), .IN2(n810), .S(n7273), .Q(n17473) );
  MUX21X1 U8380 ( .IN1(\mem0[114][4] ), .IN2(n788), .S(n7273), .Q(n17472) );
  MUX21X1 U8381 ( .IN1(\mem0[114][3] ), .IN2(n766), .S(n7273), .Q(n17471) );
  MUX21X1 U8382 ( .IN1(\mem0[114][2] ), .IN2(n744), .S(n7273), .Q(n17470) );
  MUX21X1 U8383 ( .IN1(\mem0[114][1] ), .IN2(n722), .S(n7273), .Q(n17469) );
  MUX21X1 U8384 ( .IN1(\mem0[114][0] ), .IN2(n700), .S(n7273), .Q(n17468) );
  AND2X1 U8385 ( .IN1(n7260), .IN2(n7126), .Q(n7273) );
  MUX21X1 U8386 ( .IN1(\mem0[113][7] ), .IN2(n854), .S(n7274), .Q(n17467) );
  MUX21X1 U8387 ( .IN1(\mem0[113][6] ), .IN2(n832), .S(n7274), .Q(n17466) );
  MUX21X1 U8388 ( .IN1(\mem0[113][5] ), .IN2(n810), .S(n7274), .Q(n17465) );
  MUX21X1 U8389 ( .IN1(\mem0[113][4] ), .IN2(n788), .S(n7274), .Q(n17464) );
  MUX21X1 U8390 ( .IN1(\mem0[113][3] ), .IN2(n766), .S(n7274), .Q(n17463) );
  MUX21X1 U8391 ( .IN1(\mem0[113][2] ), .IN2(n744), .S(n7274), .Q(n17462) );
  MUX21X1 U8392 ( .IN1(\mem0[113][1] ), .IN2(n722), .S(n7274), .Q(n17461) );
  MUX21X1 U8393 ( .IN1(\mem0[113][0] ), .IN2(n700), .S(n7274), .Q(n17460) );
  AND2X1 U8394 ( .IN1(n7260), .IN2(n7128), .Q(n7274) );
  MUX21X1 U8395 ( .IN1(\mem0[112][7] ), .IN2(n854), .S(n7275), .Q(n17459) );
  MUX21X1 U8396 ( .IN1(\mem0[112][6] ), .IN2(n832), .S(n7275), .Q(n17458) );
  MUX21X1 U8397 ( .IN1(\mem0[112][5] ), .IN2(n810), .S(n7275), .Q(n17457) );
  MUX21X1 U8398 ( .IN1(\mem0[112][4] ), .IN2(n788), .S(n7275), .Q(n17456) );
  MUX21X1 U8399 ( .IN1(\mem0[112][3] ), .IN2(n766), .S(n7275), .Q(n17455) );
  MUX21X1 U8400 ( .IN1(\mem0[112][2] ), .IN2(n744), .S(n7275), .Q(n17454) );
  MUX21X1 U8401 ( .IN1(\mem0[112][1] ), .IN2(n722), .S(n7275), .Q(n17453) );
  MUX21X1 U8402 ( .IN1(\mem0[112][0] ), .IN2(n700), .S(n7275), .Q(n17452) );
  AND2X1 U8403 ( .IN1(n7260), .IN2(n7130), .Q(n7275) );
  AND2X1 U8404 ( .IN1(n7276), .IN2(n7132), .Q(n7260) );
  MUX21X1 U8405 ( .IN1(\mem0[111][7] ), .IN2(n855), .S(n7277), .Q(n17451) );
  MUX21X1 U8406 ( .IN1(\mem0[111][6] ), .IN2(n833), .S(n7277), .Q(n17450) );
  MUX21X1 U8407 ( .IN1(\mem0[111][5] ), .IN2(n811), .S(n7277), .Q(n17449) );
  MUX21X1 U8408 ( .IN1(\mem0[111][4] ), .IN2(n789), .S(n7277), .Q(n17448) );
  MUX21X1 U8409 ( .IN1(\mem0[111][3] ), .IN2(n767), .S(n7277), .Q(n17447) );
  MUX21X1 U8410 ( .IN1(\mem0[111][2] ), .IN2(n745), .S(n7277), .Q(n17446) );
  MUX21X1 U8411 ( .IN1(\mem0[111][1] ), .IN2(n723), .S(n7277), .Q(n17445) );
  MUX21X1 U8412 ( .IN1(\mem0[111][0] ), .IN2(n701), .S(n7277), .Q(n17444) );
  AND2X1 U8413 ( .IN1(n7278), .IN2(n7099), .Q(n7277) );
  MUX21X1 U8414 ( .IN1(\mem0[110][7] ), .IN2(n855), .S(n7279), .Q(n17443) );
  MUX21X1 U8415 ( .IN1(\mem0[110][6] ), .IN2(n833), .S(n7279), .Q(n17442) );
  MUX21X1 U8416 ( .IN1(\mem0[110][5] ), .IN2(n811), .S(n7279), .Q(n17441) );
  MUX21X1 U8417 ( .IN1(\mem0[110][4] ), .IN2(n789), .S(n7279), .Q(n17440) );
  MUX21X1 U8418 ( .IN1(\mem0[110][3] ), .IN2(n767), .S(n7279), .Q(n17439) );
  MUX21X1 U8419 ( .IN1(\mem0[110][2] ), .IN2(n745), .S(n7279), .Q(n17438) );
  MUX21X1 U8420 ( .IN1(\mem0[110][1] ), .IN2(n723), .S(n7279), .Q(n17437) );
  MUX21X1 U8421 ( .IN1(\mem0[110][0] ), .IN2(n701), .S(n7279), .Q(n17436) );
  AND2X1 U8422 ( .IN1(n7278), .IN2(n7102), .Q(n7279) );
  MUX21X1 U8423 ( .IN1(\mem0[109][7] ), .IN2(n855), .S(n7280), .Q(n17435) );
  MUX21X1 U8424 ( .IN1(\mem0[109][6] ), .IN2(n833), .S(n7280), .Q(n17434) );
  MUX21X1 U8425 ( .IN1(\mem0[109][5] ), .IN2(n811), .S(n7280), .Q(n17433) );
  MUX21X1 U8426 ( .IN1(\mem0[109][4] ), .IN2(n789), .S(n7280), .Q(n17432) );
  MUX21X1 U8427 ( .IN1(\mem0[109][3] ), .IN2(n767), .S(n7280), .Q(n17431) );
  MUX21X1 U8428 ( .IN1(\mem0[109][2] ), .IN2(n745), .S(n7280), .Q(n17430) );
  MUX21X1 U8429 ( .IN1(\mem0[109][1] ), .IN2(n723), .S(n7280), .Q(n17429) );
  MUX21X1 U8430 ( .IN1(\mem0[109][0] ), .IN2(n701), .S(n7280), .Q(n17428) );
  AND2X1 U8431 ( .IN1(n7278), .IN2(n7104), .Q(n7280) );
  MUX21X1 U8432 ( .IN1(\mem0[108][7] ), .IN2(n855), .S(n7281), .Q(n17427) );
  MUX21X1 U8433 ( .IN1(\mem0[108][6] ), .IN2(n833), .S(n7281), .Q(n17426) );
  MUX21X1 U8434 ( .IN1(\mem0[108][5] ), .IN2(n811), .S(n7281), .Q(n17425) );
  MUX21X1 U8435 ( .IN1(\mem0[108][4] ), .IN2(n789), .S(n7281), .Q(n17424) );
  MUX21X1 U8436 ( .IN1(\mem0[108][3] ), .IN2(n767), .S(n7281), .Q(n17423) );
  MUX21X1 U8437 ( .IN1(\mem0[108][2] ), .IN2(n745), .S(n7281), .Q(n17422) );
  MUX21X1 U8438 ( .IN1(\mem0[108][1] ), .IN2(n723), .S(n7281), .Q(n17421) );
  MUX21X1 U8439 ( .IN1(\mem0[108][0] ), .IN2(n701), .S(n7281), .Q(n17420) );
  AND2X1 U8440 ( .IN1(n7278), .IN2(n7106), .Q(n7281) );
  MUX21X1 U8441 ( .IN1(\mem0[107][7] ), .IN2(n855), .S(n7282), .Q(n17419) );
  MUX21X1 U8442 ( .IN1(\mem0[107][6] ), .IN2(n833), .S(n7282), .Q(n17418) );
  MUX21X1 U8443 ( .IN1(\mem0[107][5] ), .IN2(n811), .S(n7282), .Q(n17417) );
  MUX21X1 U8444 ( .IN1(\mem0[107][4] ), .IN2(n789), .S(n7282), .Q(n17416) );
  MUX21X1 U8445 ( .IN1(\mem0[107][3] ), .IN2(n767), .S(n7282), .Q(n17415) );
  MUX21X1 U8446 ( .IN1(\mem0[107][2] ), .IN2(n745), .S(n7282), .Q(n17414) );
  MUX21X1 U8447 ( .IN1(\mem0[107][1] ), .IN2(n723), .S(n7282), .Q(n17413) );
  MUX21X1 U8448 ( .IN1(\mem0[107][0] ), .IN2(n701), .S(n7282), .Q(n17412) );
  AND2X1 U8449 ( .IN1(n7278), .IN2(n7108), .Q(n7282) );
  MUX21X1 U8450 ( .IN1(\mem0[106][7] ), .IN2(n855), .S(n7283), .Q(n17411) );
  MUX21X1 U8451 ( .IN1(\mem0[106][6] ), .IN2(n833), .S(n7283), .Q(n17410) );
  MUX21X1 U8452 ( .IN1(\mem0[106][5] ), .IN2(n811), .S(n7283), .Q(n17409) );
  MUX21X1 U8453 ( .IN1(\mem0[106][4] ), .IN2(n789), .S(n7283), .Q(n17408) );
  MUX21X1 U8454 ( .IN1(\mem0[106][3] ), .IN2(n767), .S(n7283), .Q(n17407) );
  MUX21X1 U8455 ( .IN1(\mem0[106][2] ), .IN2(n745), .S(n7283), .Q(n17406) );
  MUX21X1 U8456 ( .IN1(\mem0[106][1] ), .IN2(n723), .S(n7283), .Q(n17405) );
  MUX21X1 U8457 ( .IN1(\mem0[106][0] ), .IN2(n701), .S(n7283), .Q(n17404) );
  AND2X1 U8458 ( .IN1(n7278), .IN2(n7110), .Q(n7283) );
  MUX21X1 U8459 ( .IN1(\mem0[105][7] ), .IN2(n855), .S(n7284), .Q(n17403) );
  MUX21X1 U8460 ( .IN1(\mem0[105][6] ), .IN2(n833), .S(n7284), .Q(n17402) );
  MUX21X1 U8461 ( .IN1(\mem0[105][5] ), .IN2(n811), .S(n7284), .Q(n17401) );
  MUX21X1 U8462 ( .IN1(\mem0[105][4] ), .IN2(n789), .S(n7284), .Q(n17400) );
  MUX21X1 U8463 ( .IN1(\mem0[105][3] ), .IN2(n767), .S(n7284), .Q(n17399) );
  MUX21X1 U8464 ( .IN1(\mem0[105][2] ), .IN2(n745), .S(n7284), .Q(n17398) );
  MUX21X1 U8465 ( .IN1(\mem0[105][1] ), .IN2(n723), .S(n7284), .Q(n17397) );
  MUX21X1 U8466 ( .IN1(\mem0[105][0] ), .IN2(n701), .S(n7284), .Q(n17396) );
  AND2X1 U8467 ( .IN1(n7278), .IN2(n7112), .Q(n7284) );
  MUX21X1 U8468 ( .IN1(\mem0[104][7] ), .IN2(n855), .S(n7285), .Q(n17395) );
  MUX21X1 U8469 ( .IN1(\mem0[104][6] ), .IN2(n833), .S(n7285), .Q(n17394) );
  MUX21X1 U8470 ( .IN1(\mem0[104][5] ), .IN2(n811), .S(n7285), .Q(n17393) );
  MUX21X1 U8471 ( .IN1(\mem0[104][4] ), .IN2(n789), .S(n7285), .Q(n17392) );
  MUX21X1 U8472 ( .IN1(\mem0[104][3] ), .IN2(n767), .S(n7285), .Q(n17391) );
  MUX21X1 U8473 ( .IN1(\mem0[104][2] ), .IN2(n745), .S(n7285), .Q(n17390) );
  MUX21X1 U8474 ( .IN1(\mem0[104][1] ), .IN2(n723), .S(n7285), .Q(n17389) );
  MUX21X1 U8475 ( .IN1(\mem0[104][0] ), .IN2(n701), .S(n7285), .Q(n17388) );
  AND2X1 U8476 ( .IN1(n7278), .IN2(n7114), .Q(n7285) );
  MUX21X1 U8477 ( .IN1(\mem0[103][7] ), .IN2(n855), .S(n7286), .Q(n17387) );
  MUX21X1 U8478 ( .IN1(\mem0[103][6] ), .IN2(n833), .S(n7286), .Q(n17386) );
  MUX21X1 U8479 ( .IN1(\mem0[103][5] ), .IN2(n811), .S(n7286), .Q(n17385) );
  MUX21X1 U8480 ( .IN1(\mem0[103][4] ), .IN2(n789), .S(n7286), .Q(n17384) );
  MUX21X1 U8481 ( .IN1(\mem0[103][3] ), .IN2(n767), .S(n7286), .Q(n17383) );
  MUX21X1 U8482 ( .IN1(\mem0[103][2] ), .IN2(n745), .S(n7286), .Q(n17382) );
  MUX21X1 U8483 ( .IN1(\mem0[103][1] ), .IN2(n723), .S(n7286), .Q(n17381) );
  MUX21X1 U8484 ( .IN1(\mem0[103][0] ), .IN2(n701), .S(n7286), .Q(n17380) );
  AND2X1 U8485 ( .IN1(n7278), .IN2(n7116), .Q(n7286) );
  MUX21X1 U8486 ( .IN1(\mem0[102][7] ), .IN2(n855), .S(n7287), .Q(n17379) );
  MUX21X1 U8487 ( .IN1(\mem0[102][6] ), .IN2(n833), .S(n7287), .Q(n17378) );
  MUX21X1 U8488 ( .IN1(\mem0[102][5] ), .IN2(n811), .S(n7287), .Q(n17377) );
  MUX21X1 U8489 ( .IN1(\mem0[102][4] ), .IN2(n789), .S(n7287), .Q(n17376) );
  MUX21X1 U8490 ( .IN1(\mem0[102][3] ), .IN2(n767), .S(n7287), .Q(n17375) );
  MUX21X1 U8491 ( .IN1(\mem0[102][2] ), .IN2(n745), .S(n7287), .Q(n17374) );
  MUX21X1 U8492 ( .IN1(\mem0[102][1] ), .IN2(n723), .S(n7287), .Q(n17373) );
  MUX21X1 U8493 ( .IN1(\mem0[102][0] ), .IN2(n701), .S(n7287), .Q(n17372) );
  AND2X1 U8494 ( .IN1(n7278), .IN2(n7118), .Q(n7287) );
  MUX21X1 U8495 ( .IN1(\mem0[101][7] ), .IN2(n855), .S(n7288), .Q(n17371) );
  MUX21X1 U8496 ( .IN1(\mem0[101][6] ), .IN2(n833), .S(n7288), .Q(n17370) );
  MUX21X1 U8497 ( .IN1(\mem0[101][5] ), .IN2(n811), .S(n7288), .Q(n17369) );
  MUX21X1 U8498 ( .IN1(\mem0[101][4] ), .IN2(n789), .S(n7288), .Q(n17368) );
  MUX21X1 U8499 ( .IN1(\mem0[101][3] ), .IN2(n767), .S(n7288), .Q(n17367) );
  MUX21X1 U8500 ( .IN1(\mem0[101][2] ), .IN2(n745), .S(n7288), .Q(n17366) );
  MUX21X1 U8501 ( .IN1(\mem0[101][1] ), .IN2(n723), .S(n7288), .Q(n17365) );
  MUX21X1 U8502 ( .IN1(\mem0[101][0] ), .IN2(n701), .S(n7288), .Q(n17364) );
  AND2X1 U8503 ( .IN1(n7278), .IN2(n7120), .Q(n7288) );
  MUX21X1 U8504 ( .IN1(\mem0[100][7] ), .IN2(n855), .S(n7289), .Q(n17363) );
  MUX21X1 U8505 ( .IN1(\mem0[100][6] ), .IN2(n833), .S(n7289), .Q(n17362) );
  MUX21X1 U8506 ( .IN1(\mem0[100][5] ), .IN2(n811), .S(n7289), .Q(n17361) );
  MUX21X1 U8507 ( .IN1(\mem0[100][4] ), .IN2(n789), .S(n7289), .Q(n17360) );
  MUX21X1 U8508 ( .IN1(\mem0[100][3] ), .IN2(n767), .S(n7289), .Q(n17359) );
  MUX21X1 U8509 ( .IN1(\mem0[100][2] ), .IN2(n745), .S(n7289), .Q(n17358) );
  MUX21X1 U8510 ( .IN1(\mem0[100][1] ), .IN2(n723), .S(n7289), .Q(n17357) );
  MUX21X1 U8511 ( .IN1(\mem0[100][0] ), .IN2(n701), .S(n7289), .Q(n17356) );
  AND2X1 U8512 ( .IN1(n7278), .IN2(n7122), .Q(n7289) );
  MUX21X1 U8513 ( .IN1(\mem0[99][7] ), .IN2(n856), .S(n7290), .Q(n17355) );
  MUX21X1 U8514 ( .IN1(\mem0[99][6] ), .IN2(n834), .S(n7290), .Q(n17354) );
  MUX21X1 U8515 ( .IN1(\mem0[99][5] ), .IN2(n812), .S(n7290), .Q(n17353) );
  MUX21X1 U8516 ( .IN1(\mem0[99][4] ), .IN2(n790), .S(n7290), .Q(n17352) );
  MUX21X1 U8517 ( .IN1(\mem0[99][3] ), .IN2(n768), .S(n7290), .Q(n17351) );
  MUX21X1 U8518 ( .IN1(\mem0[99][2] ), .IN2(n746), .S(n7290), .Q(n17350) );
  MUX21X1 U8519 ( .IN1(\mem0[99][1] ), .IN2(n724), .S(n7290), .Q(n17349) );
  MUX21X1 U8520 ( .IN1(\mem0[99][0] ), .IN2(n702), .S(n7290), .Q(n17348) );
  AND2X1 U8521 ( .IN1(n7278), .IN2(n7124), .Q(n7290) );
  MUX21X1 U8522 ( .IN1(\mem0[98][7] ), .IN2(n856), .S(n7291), .Q(n17347) );
  MUX21X1 U8523 ( .IN1(\mem0[98][6] ), .IN2(n834), .S(n7291), .Q(n17346) );
  MUX21X1 U8524 ( .IN1(\mem0[98][5] ), .IN2(n812), .S(n7291), .Q(n17345) );
  MUX21X1 U8525 ( .IN1(\mem0[98][4] ), .IN2(n790), .S(n7291), .Q(n17344) );
  MUX21X1 U8526 ( .IN1(\mem0[98][3] ), .IN2(n768), .S(n7291), .Q(n17343) );
  MUX21X1 U8527 ( .IN1(\mem0[98][2] ), .IN2(n746), .S(n7291), .Q(n17342) );
  MUX21X1 U8528 ( .IN1(\mem0[98][1] ), .IN2(n724), .S(n7291), .Q(n17341) );
  MUX21X1 U8529 ( .IN1(\mem0[98][0] ), .IN2(n702), .S(n7291), .Q(n17340) );
  AND2X1 U8530 ( .IN1(n7278), .IN2(n7126), .Q(n7291) );
  MUX21X1 U8531 ( .IN1(\mem0[97][7] ), .IN2(n856), .S(n7292), .Q(n17339) );
  MUX21X1 U8532 ( .IN1(\mem0[97][6] ), .IN2(n834), .S(n7292), .Q(n17338) );
  MUX21X1 U8533 ( .IN1(\mem0[97][5] ), .IN2(n812), .S(n7292), .Q(n17337) );
  MUX21X1 U8534 ( .IN1(\mem0[97][4] ), .IN2(n790), .S(n7292), .Q(n17336) );
  MUX21X1 U8535 ( .IN1(\mem0[97][3] ), .IN2(n768), .S(n7292), .Q(n17335) );
  MUX21X1 U8536 ( .IN1(\mem0[97][2] ), .IN2(n746), .S(n7292), .Q(n17334) );
  MUX21X1 U8537 ( .IN1(\mem0[97][1] ), .IN2(n724), .S(n7292), .Q(n17333) );
  MUX21X1 U8538 ( .IN1(\mem0[97][0] ), .IN2(n702), .S(n7292), .Q(n17332) );
  AND2X1 U8539 ( .IN1(n7278), .IN2(n7128), .Q(n7292) );
  MUX21X1 U8540 ( .IN1(\mem0[96][7] ), .IN2(n856), .S(n7293), .Q(n17331) );
  MUX21X1 U8541 ( .IN1(\mem0[96][6] ), .IN2(n834), .S(n7293), .Q(n17330) );
  MUX21X1 U8542 ( .IN1(\mem0[96][5] ), .IN2(n812), .S(n7293), .Q(n17329) );
  MUX21X1 U8543 ( .IN1(\mem0[96][4] ), .IN2(n790), .S(n7293), .Q(n17328) );
  MUX21X1 U8544 ( .IN1(\mem0[96][3] ), .IN2(n768), .S(n7293), .Q(n17327) );
  MUX21X1 U8545 ( .IN1(\mem0[96][2] ), .IN2(n746), .S(n7293), .Q(n17326) );
  MUX21X1 U8546 ( .IN1(\mem0[96][1] ), .IN2(n724), .S(n7293), .Q(n17325) );
  MUX21X1 U8547 ( .IN1(\mem0[96][0] ), .IN2(n702), .S(n7293), .Q(n17324) );
  AND2X1 U8548 ( .IN1(n7278), .IN2(n7130), .Q(n7293) );
  AND2X1 U8549 ( .IN1(n7294), .IN2(n7132), .Q(n7278) );
  MUX21X1 U8550 ( .IN1(\mem0[95][7] ), .IN2(n856), .S(n7295), .Q(n17323) );
  MUX21X1 U8551 ( .IN1(\mem0[95][6] ), .IN2(n834), .S(n7295), .Q(n17322) );
  MUX21X1 U8552 ( .IN1(\mem0[95][5] ), .IN2(n812), .S(n7295), .Q(n17321) );
  MUX21X1 U8553 ( .IN1(\mem0[95][4] ), .IN2(n790), .S(n7295), .Q(n17320) );
  MUX21X1 U8554 ( .IN1(\mem0[95][3] ), .IN2(n768), .S(n7295), .Q(n17319) );
  MUX21X1 U8555 ( .IN1(\mem0[95][2] ), .IN2(n746), .S(n7295), .Q(n17318) );
  MUX21X1 U8556 ( .IN1(\mem0[95][1] ), .IN2(n724), .S(n7295), .Q(n17317) );
  MUX21X1 U8557 ( .IN1(\mem0[95][0] ), .IN2(n702), .S(n7295), .Q(n17316) );
  AND2X1 U8558 ( .IN1(n7296), .IN2(n7099), .Q(n7295) );
  MUX21X1 U8559 ( .IN1(\mem0[94][7] ), .IN2(n856), .S(n7297), .Q(n17315) );
  MUX21X1 U8560 ( .IN1(\mem0[94][6] ), .IN2(n834), .S(n7297), .Q(n17314) );
  MUX21X1 U8561 ( .IN1(\mem0[94][5] ), .IN2(n812), .S(n7297), .Q(n17313) );
  MUX21X1 U8562 ( .IN1(\mem0[94][4] ), .IN2(n790), .S(n7297), .Q(n17312) );
  MUX21X1 U8563 ( .IN1(\mem0[94][3] ), .IN2(n768), .S(n7297), .Q(n17311) );
  MUX21X1 U8564 ( .IN1(\mem0[94][2] ), .IN2(n746), .S(n7297), .Q(n17310) );
  MUX21X1 U8565 ( .IN1(\mem0[94][1] ), .IN2(n724), .S(n7297), .Q(n17309) );
  MUX21X1 U8566 ( .IN1(\mem0[94][0] ), .IN2(n702), .S(n7297), .Q(n17308) );
  AND2X1 U8567 ( .IN1(n7296), .IN2(n7102), .Q(n7297) );
  MUX21X1 U8568 ( .IN1(\mem0[93][7] ), .IN2(n856), .S(n7298), .Q(n17307) );
  MUX21X1 U8569 ( .IN1(\mem0[93][6] ), .IN2(n834), .S(n7298), .Q(n17306) );
  MUX21X1 U8570 ( .IN1(\mem0[93][5] ), .IN2(n812), .S(n7298), .Q(n17305) );
  MUX21X1 U8571 ( .IN1(\mem0[93][4] ), .IN2(n790), .S(n7298), .Q(n17304) );
  MUX21X1 U8572 ( .IN1(\mem0[93][3] ), .IN2(n768), .S(n7298), .Q(n17303) );
  MUX21X1 U8573 ( .IN1(\mem0[93][2] ), .IN2(n746), .S(n7298), .Q(n17302) );
  MUX21X1 U8574 ( .IN1(\mem0[93][1] ), .IN2(n724), .S(n7298), .Q(n17301) );
  MUX21X1 U8575 ( .IN1(\mem0[93][0] ), .IN2(n702), .S(n7298), .Q(n17300) );
  AND2X1 U8576 ( .IN1(n7296), .IN2(n7104), .Q(n7298) );
  MUX21X1 U8577 ( .IN1(\mem0[92][7] ), .IN2(n856), .S(n7299), .Q(n17299) );
  MUX21X1 U8578 ( .IN1(\mem0[92][6] ), .IN2(n834), .S(n7299), .Q(n17298) );
  MUX21X1 U8579 ( .IN1(\mem0[92][5] ), .IN2(n812), .S(n7299), .Q(n17297) );
  MUX21X1 U8580 ( .IN1(\mem0[92][4] ), .IN2(n790), .S(n7299), .Q(n17296) );
  MUX21X1 U8581 ( .IN1(\mem0[92][3] ), .IN2(n768), .S(n7299), .Q(n17295) );
  MUX21X1 U8582 ( .IN1(\mem0[92][2] ), .IN2(n746), .S(n7299), .Q(n17294) );
  MUX21X1 U8583 ( .IN1(\mem0[92][1] ), .IN2(n724), .S(n7299), .Q(n17293) );
  MUX21X1 U8584 ( .IN1(\mem0[92][0] ), .IN2(n702), .S(n7299), .Q(n17292) );
  AND2X1 U8585 ( .IN1(n7296), .IN2(n7106), .Q(n7299) );
  MUX21X1 U8586 ( .IN1(\mem0[91][7] ), .IN2(n856), .S(n7300), .Q(n17291) );
  MUX21X1 U8587 ( .IN1(\mem0[91][6] ), .IN2(n834), .S(n7300), .Q(n17290) );
  MUX21X1 U8588 ( .IN1(\mem0[91][5] ), .IN2(n812), .S(n7300), .Q(n17289) );
  MUX21X1 U8589 ( .IN1(\mem0[91][4] ), .IN2(n790), .S(n7300), .Q(n17288) );
  MUX21X1 U8590 ( .IN1(\mem0[91][3] ), .IN2(n768), .S(n7300), .Q(n17287) );
  MUX21X1 U8591 ( .IN1(\mem0[91][2] ), .IN2(n746), .S(n7300), .Q(n17286) );
  MUX21X1 U8592 ( .IN1(\mem0[91][1] ), .IN2(n724), .S(n7300), .Q(n17285) );
  MUX21X1 U8593 ( .IN1(\mem0[91][0] ), .IN2(n702), .S(n7300), .Q(n17284) );
  AND2X1 U8594 ( .IN1(n7296), .IN2(n7108), .Q(n7300) );
  MUX21X1 U8595 ( .IN1(\mem0[90][7] ), .IN2(n856), .S(n7301), .Q(n17283) );
  MUX21X1 U8596 ( .IN1(\mem0[90][6] ), .IN2(n834), .S(n7301), .Q(n17282) );
  MUX21X1 U8597 ( .IN1(\mem0[90][5] ), .IN2(n812), .S(n7301), .Q(n17281) );
  MUX21X1 U8598 ( .IN1(\mem0[90][4] ), .IN2(n790), .S(n7301), .Q(n17280) );
  MUX21X1 U8599 ( .IN1(\mem0[90][3] ), .IN2(n768), .S(n7301), .Q(n17279) );
  MUX21X1 U8600 ( .IN1(\mem0[90][2] ), .IN2(n746), .S(n7301), .Q(n17278) );
  MUX21X1 U8601 ( .IN1(\mem0[90][1] ), .IN2(n724), .S(n7301), .Q(n17277) );
  MUX21X1 U8602 ( .IN1(\mem0[90][0] ), .IN2(n702), .S(n7301), .Q(n17276) );
  AND2X1 U8603 ( .IN1(n7296), .IN2(n7110), .Q(n7301) );
  MUX21X1 U8604 ( .IN1(\mem0[89][7] ), .IN2(n856), .S(n7302), .Q(n17275) );
  MUX21X1 U8605 ( .IN1(\mem0[89][6] ), .IN2(n834), .S(n7302), .Q(n17274) );
  MUX21X1 U8606 ( .IN1(\mem0[89][5] ), .IN2(n812), .S(n7302), .Q(n17273) );
  MUX21X1 U8607 ( .IN1(\mem0[89][4] ), .IN2(n790), .S(n7302), .Q(n17272) );
  MUX21X1 U8608 ( .IN1(\mem0[89][3] ), .IN2(n768), .S(n7302), .Q(n17271) );
  MUX21X1 U8609 ( .IN1(\mem0[89][2] ), .IN2(n746), .S(n7302), .Q(n17270) );
  MUX21X1 U8610 ( .IN1(\mem0[89][1] ), .IN2(n724), .S(n7302), .Q(n17269) );
  MUX21X1 U8611 ( .IN1(\mem0[89][0] ), .IN2(n702), .S(n7302), .Q(n17268) );
  AND2X1 U8612 ( .IN1(n7296), .IN2(n7112), .Q(n7302) );
  MUX21X1 U8613 ( .IN1(\mem0[88][7] ), .IN2(n856), .S(n7303), .Q(n17267) );
  MUX21X1 U8614 ( .IN1(\mem0[88][6] ), .IN2(n834), .S(n7303), .Q(n17266) );
  MUX21X1 U8615 ( .IN1(\mem0[88][5] ), .IN2(n812), .S(n7303), .Q(n17265) );
  MUX21X1 U8616 ( .IN1(\mem0[88][4] ), .IN2(n790), .S(n7303), .Q(n17264) );
  MUX21X1 U8617 ( .IN1(\mem0[88][3] ), .IN2(n768), .S(n7303), .Q(n17263) );
  MUX21X1 U8618 ( .IN1(\mem0[88][2] ), .IN2(n746), .S(n7303), .Q(n17262) );
  MUX21X1 U8619 ( .IN1(\mem0[88][1] ), .IN2(n724), .S(n7303), .Q(n17261) );
  MUX21X1 U8620 ( .IN1(\mem0[88][0] ), .IN2(n702), .S(n7303), .Q(n17260) );
  AND2X1 U8621 ( .IN1(n7296), .IN2(n7114), .Q(n7303) );
  MUX21X1 U8622 ( .IN1(\mem0[87][7] ), .IN2(n857), .S(n7304), .Q(n17259) );
  MUX21X1 U8623 ( .IN1(\mem0[87][6] ), .IN2(n835), .S(n7304), .Q(n17258) );
  MUX21X1 U8624 ( .IN1(\mem0[87][5] ), .IN2(n813), .S(n7304), .Q(n17257) );
  MUX21X1 U8625 ( .IN1(\mem0[87][4] ), .IN2(n791), .S(n7304), .Q(n17256) );
  MUX21X1 U8626 ( .IN1(\mem0[87][3] ), .IN2(n769), .S(n7304), .Q(n17255) );
  MUX21X1 U8627 ( .IN1(\mem0[87][2] ), .IN2(n747), .S(n7304), .Q(n17254) );
  MUX21X1 U8628 ( .IN1(\mem0[87][1] ), .IN2(n725), .S(n7304), .Q(n17253) );
  MUX21X1 U8629 ( .IN1(\mem0[87][0] ), .IN2(n703), .S(n7304), .Q(n17252) );
  AND2X1 U8630 ( .IN1(n7296), .IN2(n7116), .Q(n7304) );
  MUX21X1 U8631 ( .IN1(\mem0[86][7] ), .IN2(n857), .S(n7305), .Q(n17251) );
  MUX21X1 U8632 ( .IN1(\mem0[86][6] ), .IN2(n835), .S(n7305), .Q(n17250) );
  MUX21X1 U8633 ( .IN1(\mem0[86][5] ), .IN2(n813), .S(n7305), .Q(n17249) );
  MUX21X1 U8634 ( .IN1(\mem0[86][4] ), .IN2(n791), .S(n7305), .Q(n17248) );
  MUX21X1 U8635 ( .IN1(\mem0[86][3] ), .IN2(n769), .S(n7305), .Q(n17247) );
  MUX21X1 U8636 ( .IN1(\mem0[86][2] ), .IN2(n747), .S(n7305), .Q(n17246) );
  MUX21X1 U8637 ( .IN1(\mem0[86][1] ), .IN2(n725), .S(n7305), .Q(n17245) );
  MUX21X1 U8638 ( .IN1(\mem0[86][0] ), .IN2(n703), .S(n7305), .Q(n17244) );
  AND2X1 U8639 ( .IN1(n7296), .IN2(n7118), .Q(n7305) );
  MUX21X1 U8640 ( .IN1(\mem0[85][7] ), .IN2(n857), .S(n7306), .Q(n17243) );
  MUX21X1 U8641 ( .IN1(\mem0[85][6] ), .IN2(n835), .S(n7306), .Q(n17242) );
  MUX21X1 U8642 ( .IN1(\mem0[85][5] ), .IN2(n813), .S(n7306), .Q(n17241) );
  MUX21X1 U8643 ( .IN1(\mem0[85][4] ), .IN2(n791), .S(n7306), .Q(n17240) );
  MUX21X1 U8644 ( .IN1(\mem0[85][3] ), .IN2(n769), .S(n7306), .Q(n17239) );
  MUX21X1 U8645 ( .IN1(\mem0[85][2] ), .IN2(n747), .S(n7306), .Q(n17238) );
  MUX21X1 U8646 ( .IN1(\mem0[85][1] ), .IN2(n725), .S(n7306), .Q(n17237) );
  MUX21X1 U8647 ( .IN1(\mem0[85][0] ), .IN2(n703), .S(n7306), .Q(n17236) );
  AND2X1 U8648 ( .IN1(n7296), .IN2(n7120), .Q(n7306) );
  MUX21X1 U8649 ( .IN1(\mem0[84][7] ), .IN2(n857), .S(n7307), .Q(n17235) );
  MUX21X1 U8650 ( .IN1(\mem0[84][6] ), .IN2(n835), .S(n7307), .Q(n17234) );
  MUX21X1 U8651 ( .IN1(\mem0[84][5] ), .IN2(n813), .S(n7307), .Q(n17233) );
  MUX21X1 U8652 ( .IN1(\mem0[84][4] ), .IN2(n791), .S(n7307), .Q(n17232) );
  MUX21X1 U8653 ( .IN1(\mem0[84][3] ), .IN2(n769), .S(n7307), .Q(n17231) );
  MUX21X1 U8654 ( .IN1(\mem0[84][2] ), .IN2(n747), .S(n7307), .Q(n17230) );
  MUX21X1 U8655 ( .IN1(\mem0[84][1] ), .IN2(n725), .S(n7307), .Q(n17229) );
  MUX21X1 U8656 ( .IN1(\mem0[84][0] ), .IN2(n703), .S(n7307), .Q(n17228) );
  AND2X1 U8657 ( .IN1(n7296), .IN2(n7122), .Q(n7307) );
  MUX21X1 U8658 ( .IN1(\mem0[83][7] ), .IN2(n857), .S(n7308), .Q(n17227) );
  MUX21X1 U8659 ( .IN1(\mem0[83][6] ), .IN2(n835), .S(n7308), .Q(n17226) );
  MUX21X1 U8660 ( .IN1(\mem0[83][5] ), .IN2(n813), .S(n7308), .Q(n17225) );
  MUX21X1 U8661 ( .IN1(\mem0[83][4] ), .IN2(n791), .S(n7308), .Q(n17224) );
  MUX21X1 U8662 ( .IN1(\mem0[83][3] ), .IN2(n769), .S(n7308), .Q(n17223) );
  MUX21X1 U8663 ( .IN1(\mem0[83][2] ), .IN2(n747), .S(n7308), .Q(n17222) );
  MUX21X1 U8664 ( .IN1(\mem0[83][1] ), .IN2(n725), .S(n7308), .Q(n17221) );
  MUX21X1 U8665 ( .IN1(\mem0[83][0] ), .IN2(n703), .S(n7308), .Q(n17220) );
  AND2X1 U8666 ( .IN1(n7296), .IN2(n7124), .Q(n7308) );
  MUX21X1 U8667 ( .IN1(\mem0[82][7] ), .IN2(n857), .S(n7309), .Q(n17219) );
  MUX21X1 U8668 ( .IN1(\mem0[82][6] ), .IN2(n835), .S(n7309), .Q(n17218) );
  MUX21X1 U8669 ( .IN1(\mem0[82][5] ), .IN2(n813), .S(n7309), .Q(n17217) );
  MUX21X1 U8670 ( .IN1(\mem0[82][4] ), .IN2(n791), .S(n7309), .Q(n17216) );
  MUX21X1 U8671 ( .IN1(\mem0[82][3] ), .IN2(n769), .S(n7309), .Q(n17215) );
  MUX21X1 U8672 ( .IN1(\mem0[82][2] ), .IN2(n747), .S(n7309), .Q(n17214) );
  MUX21X1 U8673 ( .IN1(\mem0[82][1] ), .IN2(n725), .S(n7309), .Q(n17213) );
  MUX21X1 U8674 ( .IN1(\mem0[82][0] ), .IN2(n703), .S(n7309), .Q(n17212) );
  AND2X1 U8675 ( .IN1(n7296), .IN2(n7126), .Q(n7309) );
  MUX21X1 U8676 ( .IN1(\mem0[81][7] ), .IN2(n857), .S(n7310), .Q(n17211) );
  MUX21X1 U8677 ( .IN1(\mem0[81][6] ), .IN2(n835), .S(n7310), .Q(n17210) );
  MUX21X1 U8678 ( .IN1(\mem0[81][5] ), .IN2(n813), .S(n7310), .Q(n17209) );
  MUX21X1 U8679 ( .IN1(\mem0[81][4] ), .IN2(n791), .S(n7310), .Q(n17208) );
  MUX21X1 U8680 ( .IN1(\mem0[81][3] ), .IN2(n769), .S(n7310), .Q(n17207) );
  MUX21X1 U8681 ( .IN1(\mem0[81][2] ), .IN2(n747), .S(n7310), .Q(n17206) );
  MUX21X1 U8682 ( .IN1(\mem0[81][1] ), .IN2(n725), .S(n7310), .Q(n17205) );
  MUX21X1 U8683 ( .IN1(\mem0[81][0] ), .IN2(n703), .S(n7310), .Q(n17204) );
  AND2X1 U8684 ( .IN1(n7296), .IN2(n7128), .Q(n7310) );
  MUX21X1 U8685 ( .IN1(\mem0[80][7] ), .IN2(n857), .S(n7311), .Q(n17203) );
  MUX21X1 U8686 ( .IN1(\mem0[80][6] ), .IN2(n835), .S(n7311), .Q(n17202) );
  MUX21X1 U8687 ( .IN1(\mem0[80][5] ), .IN2(n813), .S(n7311), .Q(n17201) );
  MUX21X1 U8688 ( .IN1(\mem0[80][4] ), .IN2(n791), .S(n7311), .Q(n17200) );
  MUX21X1 U8689 ( .IN1(\mem0[80][3] ), .IN2(n769), .S(n7311), .Q(n17199) );
  MUX21X1 U8690 ( .IN1(\mem0[80][2] ), .IN2(n747), .S(n7311), .Q(n17198) );
  MUX21X1 U8691 ( .IN1(\mem0[80][1] ), .IN2(n725), .S(n7311), .Q(n17197) );
  MUX21X1 U8692 ( .IN1(\mem0[80][0] ), .IN2(n703), .S(n7311), .Q(n17196) );
  AND2X1 U8693 ( .IN1(n7296), .IN2(n7130), .Q(n7311) );
  AND2X1 U8694 ( .IN1(n7312), .IN2(n7132), .Q(n7296) );
  MUX21X1 U8695 ( .IN1(\mem0[79][7] ), .IN2(n857), .S(n7313), .Q(n17195) );
  MUX21X1 U8696 ( .IN1(\mem0[79][6] ), .IN2(n835), .S(n7313), .Q(n17194) );
  MUX21X1 U8697 ( .IN1(\mem0[79][5] ), .IN2(n813), .S(n7313), .Q(n17193) );
  MUX21X1 U8698 ( .IN1(\mem0[79][4] ), .IN2(n791), .S(n7313), .Q(n17192) );
  MUX21X1 U8699 ( .IN1(\mem0[79][3] ), .IN2(n769), .S(n7313), .Q(n17191) );
  MUX21X1 U8700 ( .IN1(\mem0[79][2] ), .IN2(n747), .S(n7313), .Q(n17190) );
  MUX21X1 U8701 ( .IN1(\mem0[79][1] ), .IN2(n725), .S(n7313), .Q(n17189) );
  MUX21X1 U8702 ( .IN1(\mem0[79][0] ), .IN2(n703), .S(n7313), .Q(n17188) );
  AND2X1 U8703 ( .IN1(n7314), .IN2(n7099), .Q(n7313) );
  MUX21X1 U8704 ( .IN1(\mem0[78][7] ), .IN2(n857), .S(n7315), .Q(n17187) );
  MUX21X1 U8705 ( .IN1(\mem0[78][6] ), .IN2(n835), .S(n7315), .Q(n17186) );
  MUX21X1 U8706 ( .IN1(\mem0[78][5] ), .IN2(n813), .S(n7315), .Q(n17185) );
  MUX21X1 U8707 ( .IN1(\mem0[78][4] ), .IN2(n791), .S(n7315), .Q(n17184) );
  MUX21X1 U8708 ( .IN1(\mem0[78][3] ), .IN2(n769), .S(n7315), .Q(n17183) );
  MUX21X1 U8709 ( .IN1(\mem0[78][2] ), .IN2(n747), .S(n7315), .Q(n17182) );
  MUX21X1 U8710 ( .IN1(\mem0[78][1] ), .IN2(n725), .S(n7315), .Q(n17181) );
  MUX21X1 U8711 ( .IN1(\mem0[78][0] ), .IN2(n703), .S(n7315), .Q(n17180) );
  AND2X1 U8712 ( .IN1(n7314), .IN2(n7102), .Q(n7315) );
  MUX21X1 U8713 ( .IN1(\mem0[77][7] ), .IN2(n857), .S(n7316), .Q(n17179) );
  MUX21X1 U8714 ( .IN1(\mem0[77][6] ), .IN2(n835), .S(n7316), .Q(n17178) );
  MUX21X1 U8715 ( .IN1(\mem0[77][5] ), .IN2(n813), .S(n7316), .Q(n17177) );
  MUX21X1 U8716 ( .IN1(\mem0[77][4] ), .IN2(n791), .S(n7316), .Q(n17176) );
  MUX21X1 U8717 ( .IN1(\mem0[77][3] ), .IN2(n769), .S(n7316), .Q(n17175) );
  MUX21X1 U8718 ( .IN1(\mem0[77][2] ), .IN2(n747), .S(n7316), .Q(n17174) );
  MUX21X1 U8719 ( .IN1(\mem0[77][1] ), .IN2(n725), .S(n7316), .Q(n17173) );
  MUX21X1 U8720 ( .IN1(\mem0[77][0] ), .IN2(n703), .S(n7316), .Q(n17172) );
  AND2X1 U8721 ( .IN1(n7314), .IN2(n7104), .Q(n7316) );
  MUX21X1 U8722 ( .IN1(\mem0[76][7] ), .IN2(n857), .S(n7317), .Q(n17171) );
  MUX21X1 U8723 ( .IN1(\mem0[76][6] ), .IN2(n835), .S(n7317), .Q(n17170) );
  MUX21X1 U8724 ( .IN1(\mem0[76][5] ), .IN2(n813), .S(n7317), .Q(n17169) );
  MUX21X1 U8725 ( .IN1(\mem0[76][4] ), .IN2(n791), .S(n7317), .Q(n17168) );
  MUX21X1 U8726 ( .IN1(\mem0[76][3] ), .IN2(n769), .S(n7317), .Q(n17167) );
  MUX21X1 U8727 ( .IN1(\mem0[76][2] ), .IN2(n747), .S(n7317), .Q(n17166) );
  MUX21X1 U8728 ( .IN1(\mem0[76][1] ), .IN2(n725), .S(n7317), .Q(n17165) );
  MUX21X1 U8729 ( .IN1(\mem0[76][0] ), .IN2(n703), .S(n7317), .Q(n17164) );
  AND2X1 U8730 ( .IN1(n7314), .IN2(n7106), .Q(n7317) );
  MUX21X1 U8731 ( .IN1(\mem0[75][7] ), .IN2(n858), .S(n7318), .Q(n17163) );
  MUX21X1 U8732 ( .IN1(\mem0[75][6] ), .IN2(n836), .S(n7318), .Q(n17162) );
  MUX21X1 U8733 ( .IN1(\mem0[75][5] ), .IN2(n814), .S(n7318), .Q(n17161) );
  MUX21X1 U8734 ( .IN1(\mem0[75][4] ), .IN2(n792), .S(n7318), .Q(n17160) );
  MUX21X1 U8735 ( .IN1(\mem0[75][3] ), .IN2(n770), .S(n7318), .Q(n17159) );
  MUX21X1 U8736 ( .IN1(\mem0[75][2] ), .IN2(n748), .S(n7318), .Q(n17158) );
  MUX21X1 U8737 ( .IN1(\mem0[75][1] ), .IN2(n726), .S(n7318), .Q(n17157) );
  MUX21X1 U8738 ( .IN1(\mem0[75][0] ), .IN2(n704), .S(n7318), .Q(n17156) );
  AND2X1 U8739 ( .IN1(n7314), .IN2(n7108), .Q(n7318) );
  MUX21X1 U8740 ( .IN1(\mem0[74][7] ), .IN2(n858), .S(n7319), .Q(n17155) );
  MUX21X1 U8741 ( .IN1(\mem0[74][6] ), .IN2(n836), .S(n7319), .Q(n17154) );
  MUX21X1 U8742 ( .IN1(\mem0[74][5] ), .IN2(n814), .S(n7319), .Q(n17153) );
  MUX21X1 U8743 ( .IN1(\mem0[74][4] ), .IN2(n792), .S(n7319), .Q(n17152) );
  MUX21X1 U8744 ( .IN1(\mem0[74][3] ), .IN2(n770), .S(n7319), .Q(n17151) );
  MUX21X1 U8745 ( .IN1(\mem0[74][2] ), .IN2(n748), .S(n7319), .Q(n17150) );
  MUX21X1 U8746 ( .IN1(\mem0[74][1] ), .IN2(n726), .S(n7319), .Q(n17149) );
  MUX21X1 U8747 ( .IN1(\mem0[74][0] ), .IN2(n704), .S(n7319), .Q(n17148) );
  AND2X1 U8748 ( .IN1(n7314), .IN2(n7110), .Q(n7319) );
  MUX21X1 U8749 ( .IN1(\mem0[73][7] ), .IN2(n858), .S(n7320), .Q(n17147) );
  MUX21X1 U8750 ( .IN1(\mem0[73][6] ), .IN2(n836), .S(n7320), .Q(n17146) );
  MUX21X1 U8751 ( .IN1(\mem0[73][5] ), .IN2(n814), .S(n7320), .Q(n17145) );
  MUX21X1 U8752 ( .IN1(\mem0[73][4] ), .IN2(n792), .S(n7320), .Q(n17144) );
  MUX21X1 U8753 ( .IN1(\mem0[73][3] ), .IN2(n770), .S(n7320), .Q(n17143) );
  MUX21X1 U8754 ( .IN1(\mem0[73][2] ), .IN2(n748), .S(n7320), .Q(n17142) );
  MUX21X1 U8755 ( .IN1(\mem0[73][1] ), .IN2(n726), .S(n7320), .Q(n17141) );
  MUX21X1 U8756 ( .IN1(\mem0[73][0] ), .IN2(n704), .S(n7320), .Q(n17140) );
  AND2X1 U8757 ( .IN1(n7314), .IN2(n7112), .Q(n7320) );
  MUX21X1 U8758 ( .IN1(\mem0[72][7] ), .IN2(n858), .S(n7321), .Q(n17139) );
  MUX21X1 U8759 ( .IN1(\mem0[72][6] ), .IN2(n836), .S(n7321), .Q(n17138) );
  MUX21X1 U8760 ( .IN1(\mem0[72][5] ), .IN2(n814), .S(n7321), .Q(n17137) );
  MUX21X1 U8761 ( .IN1(\mem0[72][4] ), .IN2(n792), .S(n7321), .Q(n17136) );
  MUX21X1 U8762 ( .IN1(\mem0[72][3] ), .IN2(n770), .S(n7321), .Q(n17135) );
  MUX21X1 U8763 ( .IN1(\mem0[72][2] ), .IN2(n748), .S(n7321), .Q(n17134) );
  MUX21X1 U8764 ( .IN1(\mem0[72][1] ), .IN2(n726), .S(n7321), .Q(n17133) );
  MUX21X1 U8765 ( .IN1(\mem0[72][0] ), .IN2(n704), .S(n7321), .Q(n17132) );
  AND2X1 U8766 ( .IN1(n7314), .IN2(n7114), .Q(n7321) );
  MUX21X1 U8767 ( .IN1(\mem0[71][7] ), .IN2(n858), .S(n7322), .Q(n17131) );
  MUX21X1 U8768 ( .IN1(\mem0[71][6] ), .IN2(n836), .S(n7322), .Q(n17130) );
  MUX21X1 U8769 ( .IN1(\mem0[71][5] ), .IN2(n814), .S(n7322), .Q(n17129) );
  MUX21X1 U8770 ( .IN1(\mem0[71][4] ), .IN2(n792), .S(n7322), .Q(n17128) );
  MUX21X1 U8771 ( .IN1(\mem0[71][3] ), .IN2(n770), .S(n7322), .Q(n17127) );
  MUX21X1 U8772 ( .IN1(\mem0[71][2] ), .IN2(n748), .S(n7322), .Q(n17126) );
  MUX21X1 U8773 ( .IN1(\mem0[71][1] ), .IN2(n726), .S(n7322), .Q(n17125) );
  MUX21X1 U8774 ( .IN1(\mem0[71][0] ), .IN2(n704), .S(n7322), .Q(n17124) );
  AND2X1 U8775 ( .IN1(n7314), .IN2(n7116), .Q(n7322) );
  MUX21X1 U8776 ( .IN1(\mem0[70][7] ), .IN2(n858), .S(n7323), .Q(n17123) );
  MUX21X1 U8777 ( .IN1(\mem0[70][6] ), .IN2(n836), .S(n7323), .Q(n17122) );
  MUX21X1 U8778 ( .IN1(\mem0[70][5] ), .IN2(n814), .S(n7323), .Q(n17121) );
  MUX21X1 U8779 ( .IN1(\mem0[70][4] ), .IN2(n792), .S(n7323), .Q(n17120) );
  MUX21X1 U8780 ( .IN1(\mem0[70][3] ), .IN2(n770), .S(n7323), .Q(n17119) );
  MUX21X1 U8781 ( .IN1(\mem0[70][2] ), .IN2(n748), .S(n7323), .Q(n17118) );
  MUX21X1 U8782 ( .IN1(\mem0[70][1] ), .IN2(n726), .S(n7323), .Q(n17117) );
  MUX21X1 U8783 ( .IN1(\mem0[70][0] ), .IN2(n704), .S(n7323), .Q(n17116) );
  AND2X1 U8784 ( .IN1(n7314), .IN2(n7118), .Q(n7323) );
  MUX21X1 U8785 ( .IN1(\mem0[69][7] ), .IN2(n858), .S(n7324), .Q(n17115) );
  MUX21X1 U8786 ( .IN1(\mem0[69][6] ), .IN2(n836), .S(n7324), .Q(n17114) );
  MUX21X1 U8787 ( .IN1(\mem0[69][5] ), .IN2(n814), .S(n7324), .Q(n17113) );
  MUX21X1 U8788 ( .IN1(\mem0[69][4] ), .IN2(n792), .S(n7324), .Q(n17112) );
  MUX21X1 U8789 ( .IN1(\mem0[69][3] ), .IN2(n770), .S(n7324), .Q(n17111) );
  MUX21X1 U8790 ( .IN1(\mem0[69][2] ), .IN2(n748), .S(n7324), .Q(n17110) );
  MUX21X1 U8791 ( .IN1(\mem0[69][1] ), .IN2(n726), .S(n7324), .Q(n17109) );
  MUX21X1 U8792 ( .IN1(\mem0[69][0] ), .IN2(n704), .S(n7324), .Q(n17108) );
  AND2X1 U8793 ( .IN1(n7314), .IN2(n7120), .Q(n7324) );
  MUX21X1 U8794 ( .IN1(\mem0[68][7] ), .IN2(n858), .S(n7325), .Q(n17107) );
  MUX21X1 U8795 ( .IN1(\mem0[68][6] ), .IN2(n836), .S(n7325), .Q(n17106) );
  MUX21X1 U8796 ( .IN1(\mem0[68][5] ), .IN2(n814), .S(n7325), .Q(n17105) );
  MUX21X1 U8797 ( .IN1(\mem0[68][4] ), .IN2(n792), .S(n7325), .Q(n17104) );
  MUX21X1 U8798 ( .IN1(\mem0[68][3] ), .IN2(n770), .S(n7325), .Q(n17103) );
  MUX21X1 U8799 ( .IN1(\mem0[68][2] ), .IN2(n748), .S(n7325), .Q(n17102) );
  MUX21X1 U8800 ( .IN1(\mem0[68][1] ), .IN2(n726), .S(n7325), .Q(n17101) );
  MUX21X1 U8801 ( .IN1(\mem0[68][0] ), .IN2(n704), .S(n7325), .Q(n17100) );
  AND2X1 U8802 ( .IN1(n7314), .IN2(n7122), .Q(n7325) );
  MUX21X1 U8803 ( .IN1(\mem0[67][7] ), .IN2(n858), .S(n7326), .Q(n17099) );
  MUX21X1 U8804 ( .IN1(\mem0[67][6] ), .IN2(n836), .S(n7326), .Q(n17098) );
  MUX21X1 U8805 ( .IN1(\mem0[67][5] ), .IN2(n814), .S(n7326), .Q(n17097) );
  MUX21X1 U8806 ( .IN1(\mem0[67][4] ), .IN2(n792), .S(n7326), .Q(n17096) );
  MUX21X1 U8807 ( .IN1(\mem0[67][3] ), .IN2(n770), .S(n7326), .Q(n17095) );
  MUX21X1 U8808 ( .IN1(\mem0[67][2] ), .IN2(n748), .S(n7326), .Q(n17094) );
  MUX21X1 U8809 ( .IN1(\mem0[67][1] ), .IN2(n726), .S(n7326), .Q(n17093) );
  MUX21X1 U8810 ( .IN1(\mem0[67][0] ), .IN2(n704), .S(n7326), .Q(n17092) );
  AND2X1 U8811 ( .IN1(n7314), .IN2(n7124), .Q(n7326) );
  MUX21X1 U8812 ( .IN1(\mem0[66][7] ), .IN2(n858), .S(n7327), .Q(n17091) );
  MUX21X1 U8813 ( .IN1(\mem0[66][6] ), .IN2(n836), .S(n7327), .Q(n17090) );
  MUX21X1 U8814 ( .IN1(\mem0[66][5] ), .IN2(n814), .S(n7327), .Q(n17089) );
  MUX21X1 U8815 ( .IN1(\mem0[66][4] ), .IN2(n792), .S(n7327), .Q(n17088) );
  MUX21X1 U8816 ( .IN1(\mem0[66][3] ), .IN2(n770), .S(n7327), .Q(n17087) );
  MUX21X1 U8817 ( .IN1(\mem0[66][2] ), .IN2(n748), .S(n7327), .Q(n17086) );
  MUX21X1 U8818 ( .IN1(\mem0[66][1] ), .IN2(n726), .S(n7327), .Q(n17085) );
  MUX21X1 U8819 ( .IN1(\mem0[66][0] ), .IN2(n704), .S(n7327), .Q(n17084) );
  AND2X1 U8820 ( .IN1(n7314), .IN2(n7126), .Q(n7327) );
  MUX21X1 U8821 ( .IN1(\mem0[65][7] ), .IN2(n858), .S(n7328), .Q(n17083) );
  MUX21X1 U8822 ( .IN1(\mem0[65][6] ), .IN2(n836), .S(n7328), .Q(n17082) );
  MUX21X1 U8823 ( .IN1(\mem0[65][5] ), .IN2(n814), .S(n7328), .Q(n17081) );
  MUX21X1 U8824 ( .IN1(\mem0[65][4] ), .IN2(n792), .S(n7328), .Q(n17080) );
  MUX21X1 U8825 ( .IN1(\mem0[65][3] ), .IN2(n770), .S(n7328), .Q(n17079) );
  MUX21X1 U8826 ( .IN1(\mem0[65][2] ), .IN2(n748), .S(n7328), .Q(n17078) );
  MUX21X1 U8827 ( .IN1(\mem0[65][1] ), .IN2(n726), .S(n7328), .Q(n17077) );
  MUX21X1 U8828 ( .IN1(\mem0[65][0] ), .IN2(n704), .S(n7328), .Q(n17076) );
  AND2X1 U8829 ( .IN1(n7314), .IN2(n7128), .Q(n7328) );
  MUX21X1 U8830 ( .IN1(\mem0[64][7] ), .IN2(n858), .S(n7329), .Q(n17075) );
  MUX21X1 U8831 ( .IN1(\mem0[64][6] ), .IN2(n836), .S(n7329), .Q(n17074) );
  MUX21X1 U8832 ( .IN1(\mem0[64][5] ), .IN2(n814), .S(n7329), .Q(n17073) );
  MUX21X1 U8833 ( .IN1(\mem0[64][4] ), .IN2(n792), .S(n7329), .Q(n17072) );
  MUX21X1 U8834 ( .IN1(\mem0[64][3] ), .IN2(n770), .S(n7329), .Q(n17071) );
  MUX21X1 U8835 ( .IN1(\mem0[64][2] ), .IN2(n748), .S(n7329), .Q(n17070) );
  MUX21X1 U8836 ( .IN1(\mem0[64][1] ), .IN2(n726), .S(n7329), .Q(n17069) );
  MUX21X1 U8837 ( .IN1(\mem0[64][0] ), .IN2(n704), .S(n7329), .Q(n17068) );
  AND2X1 U8838 ( .IN1(n7314), .IN2(n7130), .Q(n7329) );
  AND2X1 U8839 ( .IN1(n7330), .IN2(n7132), .Q(n7314) );
  MUX21X1 U8840 ( .IN1(\mem0[63][7] ), .IN2(n859), .S(n7331), .Q(n17067) );
  MUX21X1 U8841 ( .IN1(\mem0[63][6] ), .IN2(n837), .S(n7331), .Q(n17066) );
  MUX21X1 U8842 ( .IN1(\mem0[63][5] ), .IN2(n815), .S(n7331), .Q(n17065) );
  MUX21X1 U8843 ( .IN1(\mem0[63][4] ), .IN2(n793), .S(n7331), .Q(n17064) );
  MUX21X1 U8844 ( .IN1(\mem0[63][3] ), .IN2(n771), .S(n7331), .Q(n17063) );
  MUX21X1 U8845 ( .IN1(\mem0[63][2] ), .IN2(n749), .S(n7331), .Q(n17062) );
  MUX21X1 U8846 ( .IN1(\mem0[63][1] ), .IN2(n727), .S(n7331), .Q(n17061) );
  MUX21X1 U8847 ( .IN1(\mem0[63][0] ), .IN2(n705), .S(n7331), .Q(n17060) );
  AND2X1 U8848 ( .IN1(n7332), .IN2(n7099), .Q(n7331) );
  MUX21X1 U8849 ( .IN1(\mem0[62][7] ), .IN2(n859), .S(n7333), .Q(n17059) );
  MUX21X1 U8850 ( .IN1(\mem0[62][6] ), .IN2(n837), .S(n7333), .Q(n17058) );
  MUX21X1 U8851 ( .IN1(\mem0[62][5] ), .IN2(n815), .S(n7333), .Q(n17057) );
  MUX21X1 U8852 ( .IN1(\mem0[62][4] ), .IN2(n793), .S(n7333), .Q(n17056) );
  MUX21X1 U8853 ( .IN1(\mem0[62][3] ), .IN2(n771), .S(n7333), .Q(n17055) );
  MUX21X1 U8854 ( .IN1(\mem0[62][2] ), .IN2(n749), .S(n7333), .Q(n17054) );
  MUX21X1 U8855 ( .IN1(\mem0[62][1] ), .IN2(n727), .S(n7333), .Q(n17053) );
  MUX21X1 U8856 ( .IN1(\mem0[62][0] ), .IN2(n705), .S(n7333), .Q(n17052) );
  AND2X1 U8857 ( .IN1(n7332), .IN2(n7102), .Q(n7333) );
  MUX21X1 U8858 ( .IN1(\mem0[61][7] ), .IN2(n859), .S(n7334), .Q(n17051) );
  MUX21X1 U8859 ( .IN1(\mem0[61][6] ), .IN2(n837), .S(n7334), .Q(n17050) );
  MUX21X1 U8860 ( .IN1(\mem0[61][5] ), .IN2(n815), .S(n7334), .Q(n17049) );
  MUX21X1 U8861 ( .IN1(\mem0[61][4] ), .IN2(n793), .S(n7334), .Q(n17048) );
  MUX21X1 U8862 ( .IN1(\mem0[61][3] ), .IN2(n771), .S(n7334), .Q(n17047) );
  MUX21X1 U8863 ( .IN1(\mem0[61][2] ), .IN2(n749), .S(n7334), .Q(n17046) );
  MUX21X1 U8864 ( .IN1(\mem0[61][1] ), .IN2(n727), .S(n7334), .Q(n17045) );
  MUX21X1 U8865 ( .IN1(\mem0[61][0] ), .IN2(n705), .S(n7334), .Q(n17044) );
  AND2X1 U8866 ( .IN1(n7332), .IN2(n7104), .Q(n7334) );
  MUX21X1 U8867 ( .IN1(\mem0[60][7] ), .IN2(n859), .S(n7335), .Q(n17043) );
  MUX21X1 U8868 ( .IN1(\mem0[60][6] ), .IN2(n837), .S(n7335), .Q(n17042) );
  MUX21X1 U8869 ( .IN1(\mem0[60][5] ), .IN2(n815), .S(n7335), .Q(n17041) );
  MUX21X1 U8870 ( .IN1(\mem0[60][4] ), .IN2(n793), .S(n7335), .Q(n17040) );
  MUX21X1 U8871 ( .IN1(\mem0[60][3] ), .IN2(n771), .S(n7335), .Q(n17039) );
  MUX21X1 U8872 ( .IN1(\mem0[60][2] ), .IN2(n749), .S(n7335), .Q(n17038) );
  MUX21X1 U8873 ( .IN1(\mem0[60][1] ), .IN2(n727), .S(n7335), .Q(n17037) );
  MUX21X1 U8874 ( .IN1(\mem0[60][0] ), .IN2(n705), .S(n7335), .Q(n17036) );
  AND2X1 U8875 ( .IN1(n7332), .IN2(n7106), .Q(n7335) );
  MUX21X1 U8876 ( .IN1(\mem0[59][7] ), .IN2(n859), .S(n7336), .Q(n17035) );
  MUX21X1 U8877 ( .IN1(\mem0[59][6] ), .IN2(n837), .S(n7336), .Q(n17034) );
  MUX21X1 U8878 ( .IN1(\mem0[59][5] ), .IN2(n815), .S(n7336), .Q(n17033) );
  MUX21X1 U8879 ( .IN1(\mem0[59][4] ), .IN2(n793), .S(n7336), .Q(n17032) );
  MUX21X1 U8880 ( .IN1(\mem0[59][3] ), .IN2(n771), .S(n7336), .Q(n17031) );
  MUX21X1 U8881 ( .IN1(\mem0[59][2] ), .IN2(n749), .S(n7336), .Q(n17030) );
  MUX21X1 U8882 ( .IN1(\mem0[59][1] ), .IN2(n727), .S(n7336), .Q(n17029) );
  MUX21X1 U8883 ( .IN1(\mem0[59][0] ), .IN2(n705), .S(n7336), .Q(n17028) );
  AND2X1 U8884 ( .IN1(n7332), .IN2(n7108), .Q(n7336) );
  MUX21X1 U8885 ( .IN1(\mem0[58][7] ), .IN2(n859), .S(n7337), .Q(n17027) );
  MUX21X1 U8886 ( .IN1(\mem0[58][6] ), .IN2(n837), .S(n7337), .Q(n17026) );
  MUX21X1 U8887 ( .IN1(\mem0[58][5] ), .IN2(n815), .S(n7337), .Q(n17025) );
  MUX21X1 U8888 ( .IN1(\mem0[58][4] ), .IN2(n793), .S(n7337), .Q(n17024) );
  MUX21X1 U8889 ( .IN1(\mem0[58][3] ), .IN2(n771), .S(n7337), .Q(n17023) );
  MUX21X1 U8890 ( .IN1(\mem0[58][2] ), .IN2(n749), .S(n7337), .Q(n17022) );
  MUX21X1 U8891 ( .IN1(\mem0[58][1] ), .IN2(n727), .S(n7337), .Q(n17021) );
  MUX21X1 U8892 ( .IN1(\mem0[58][0] ), .IN2(n705), .S(n7337), .Q(n17020) );
  AND2X1 U8893 ( .IN1(n7332), .IN2(n7110), .Q(n7337) );
  MUX21X1 U8894 ( .IN1(\mem0[57][7] ), .IN2(n859), .S(n7338), .Q(n17019) );
  MUX21X1 U8895 ( .IN1(\mem0[57][6] ), .IN2(n837), .S(n7338), .Q(n17018) );
  MUX21X1 U8896 ( .IN1(\mem0[57][5] ), .IN2(n815), .S(n7338), .Q(n17017) );
  MUX21X1 U8897 ( .IN1(\mem0[57][4] ), .IN2(n793), .S(n7338), .Q(n17016) );
  MUX21X1 U8898 ( .IN1(\mem0[57][3] ), .IN2(n771), .S(n7338), .Q(n17015) );
  MUX21X1 U8899 ( .IN1(\mem0[57][2] ), .IN2(n749), .S(n7338), .Q(n17014) );
  MUX21X1 U8900 ( .IN1(\mem0[57][1] ), .IN2(n727), .S(n7338), .Q(n17013) );
  MUX21X1 U8901 ( .IN1(\mem0[57][0] ), .IN2(n705), .S(n7338), .Q(n17012) );
  AND2X1 U8902 ( .IN1(n7332), .IN2(n7112), .Q(n7338) );
  MUX21X1 U8903 ( .IN1(\mem0[56][7] ), .IN2(n859), .S(n7339), .Q(n17011) );
  MUX21X1 U8904 ( .IN1(\mem0[56][6] ), .IN2(n837), .S(n7339), .Q(n17010) );
  MUX21X1 U8905 ( .IN1(\mem0[56][5] ), .IN2(n815), .S(n7339), .Q(n17009) );
  MUX21X1 U8906 ( .IN1(\mem0[56][4] ), .IN2(n793), .S(n7339), .Q(n17008) );
  MUX21X1 U8907 ( .IN1(\mem0[56][3] ), .IN2(n771), .S(n7339), .Q(n17007) );
  MUX21X1 U8908 ( .IN1(\mem0[56][2] ), .IN2(n749), .S(n7339), .Q(n17006) );
  MUX21X1 U8909 ( .IN1(\mem0[56][1] ), .IN2(n727), .S(n7339), .Q(n17005) );
  MUX21X1 U8910 ( .IN1(\mem0[56][0] ), .IN2(n705), .S(n7339), .Q(n17004) );
  AND2X1 U8911 ( .IN1(n7332), .IN2(n7114), .Q(n7339) );
  MUX21X1 U8912 ( .IN1(\mem0[55][7] ), .IN2(n859), .S(n7340), .Q(n17003) );
  MUX21X1 U8913 ( .IN1(\mem0[55][6] ), .IN2(n837), .S(n7340), .Q(n17002) );
  MUX21X1 U8914 ( .IN1(\mem0[55][5] ), .IN2(n815), .S(n7340), .Q(n17001) );
  MUX21X1 U8915 ( .IN1(\mem0[55][4] ), .IN2(n793), .S(n7340), .Q(n17000) );
  MUX21X1 U8916 ( .IN1(\mem0[55][3] ), .IN2(n771), .S(n7340), .Q(n16999) );
  MUX21X1 U8917 ( .IN1(\mem0[55][2] ), .IN2(n749), .S(n7340), .Q(n16998) );
  MUX21X1 U8918 ( .IN1(\mem0[55][1] ), .IN2(n727), .S(n7340), .Q(n16997) );
  MUX21X1 U8919 ( .IN1(\mem0[55][0] ), .IN2(n705), .S(n7340), .Q(n16996) );
  AND2X1 U8920 ( .IN1(n7332), .IN2(n7116), .Q(n7340) );
  MUX21X1 U8921 ( .IN1(\mem0[54][7] ), .IN2(n859), .S(n7341), .Q(n16995) );
  MUX21X1 U8922 ( .IN1(\mem0[54][6] ), .IN2(n837), .S(n7341), .Q(n16994) );
  MUX21X1 U8923 ( .IN1(\mem0[54][5] ), .IN2(n815), .S(n7341), .Q(n16993) );
  MUX21X1 U8924 ( .IN1(\mem0[54][4] ), .IN2(n793), .S(n7341), .Q(n16992) );
  MUX21X1 U8925 ( .IN1(\mem0[54][3] ), .IN2(n771), .S(n7341), .Q(n16991) );
  MUX21X1 U8926 ( .IN1(\mem0[54][2] ), .IN2(n749), .S(n7341), .Q(n16990) );
  MUX21X1 U8927 ( .IN1(\mem0[54][1] ), .IN2(n727), .S(n7341), .Q(n16989) );
  MUX21X1 U8928 ( .IN1(\mem0[54][0] ), .IN2(n705), .S(n7341), .Q(n16988) );
  AND2X1 U8929 ( .IN1(n7332), .IN2(n7118), .Q(n7341) );
  MUX21X1 U8930 ( .IN1(\mem0[53][7] ), .IN2(n859), .S(n7342), .Q(n16987) );
  MUX21X1 U8931 ( .IN1(\mem0[53][6] ), .IN2(n837), .S(n7342), .Q(n16986) );
  MUX21X1 U8932 ( .IN1(\mem0[53][5] ), .IN2(n815), .S(n7342), .Q(n16985) );
  MUX21X1 U8933 ( .IN1(\mem0[53][4] ), .IN2(n793), .S(n7342), .Q(n16984) );
  MUX21X1 U8934 ( .IN1(\mem0[53][3] ), .IN2(n771), .S(n7342), .Q(n16983) );
  MUX21X1 U8935 ( .IN1(\mem0[53][2] ), .IN2(n749), .S(n7342), .Q(n16982) );
  MUX21X1 U8936 ( .IN1(\mem0[53][1] ), .IN2(n727), .S(n7342), .Q(n16981) );
  MUX21X1 U8937 ( .IN1(\mem0[53][0] ), .IN2(n705), .S(n7342), .Q(n16980) );
  AND2X1 U8938 ( .IN1(n7332), .IN2(n7120), .Q(n7342) );
  MUX21X1 U8939 ( .IN1(\mem0[52][7] ), .IN2(n859), .S(n7343), .Q(n16979) );
  MUX21X1 U8940 ( .IN1(\mem0[52][6] ), .IN2(n837), .S(n7343), .Q(n16978) );
  MUX21X1 U8941 ( .IN1(\mem0[52][5] ), .IN2(n815), .S(n7343), .Q(n16977) );
  MUX21X1 U8942 ( .IN1(\mem0[52][4] ), .IN2(n793), .S(n7343), .Q(n16976) );
  MUX21X1 U8943 ( .IN1(\mem0[52][3] ), .IN2(n771), .S(n7343), .Q(n16975) );
  MUX21X1 U8944 ( .IN1(\mem0[52][2] ), .IN2(n749), .S(n7343), .Q(n16974) );
  MUX21X1 U8945 ( .IN1(\mem0[52][1] ), .IN2(n727), .S(n7343), .Q(n16973) );
  MUX21X1 U8946 ( .IN1(\mem0[52][0] ), .IN2(n705), .S(n7343), .Q(n16972) );
  AND2X1 U8947 ( .IN1(n7332), .IN2(n7122), .Q(n7343) );
  MUX21X1 U8948 ( .IN1(\mem0[51][7] ), .IN2(n860), .S(n7344), .Q(n16971) );
  MUX21X1 U8949 ( .IN1(\mem0[51][6] ), .IN2(n838), .S(n7344), .Q(n16970) );
  MUX21X1 U8950 ( .IN1(\mem0[51][5] ), .IN2(n816), .S(n7344), .Q(n16969) );
  MUX21X1 U8951 ( .IN1(\mem0[51][4] ), .IN2(n794), .S(n7344), .Q(n16968) );
  MUX21X1 U8952 ( .IN1(\mem0[51][3] ), .IN2(n772), .S(n7344), .Q(n16967) );
  MUX21X1 U8953 ( .IN1(\mem0[51][2] ), .IN2(n750), .S(n7344), .Q(n16966) );
  MUX21X1 U8954 ( .IN1(\mem0[51][1] ), .IN2(n728), .S(n7344), .Q(n16965) );
  MUX21X1 U8955 ( .IN1(\mem0[51][0] ), .IN2(n706), .S(n7344), .Q(n16964) );
  AND2X1 U8956 ( .IN1(n7332), .IN2(n7124), .Q(n7344) );
  MUX21X1 U8957 ( .IN1(\mem0[50][7] ), .IN2(n860), .S(n7345), .Q(n16963) );
  MUX21X1 U8958 ( .IN1(\mem0[50][6] ), .IN2(n838), .S(n7345), .Q(n16962) );
  MUX21X1 U8959 ( .IN1(\mem0[50][5] ), .IN2(n816), .S(n7345), .Q(n16961) );
  MUX21X1 U8960 ( .IN1(\mem0[50][4] ), .IN2(n794), .S(n7345), .Q(n16960) );
  MUX21X1 U8961 ( .IN1(\mem0[50][3] ), .IN2(n772), .S(n7345), .Q(n16959) );
  MUX21X1 U8962 ( .IN1(\mem0[50][2] ), .IN2(n750), .S(n7345), .Q(n16958) );
  MUX21X1 U8963 ( .IN1(\mem0[50][1] ), .IN2(n728), .S(n7345), .Q(n16957) );
  MUX21X1 U8964 ( .IN1(\mem0[50][0] ), .IN2(n706), .S(n7345), .Q(n16956) );
  AND2X1 U8965 ( .IN1(n7332), .IN2(n7126), .Q(n7345) );
  MUX21X1 U8966 ( .IN1(\mem0[49][7] ), .IN2(n860), .S(n7346), .Q(n16955) );
  MUX21X1 U8967 ( .IN1(\mem0[49][6] ), .IN2(n838), .S(n7346), .Q(n16954) );
  MUX21X1 U8968 ( .IN1(\mem0[49][5] ), .IN2(n816), .S(n7346), .Q(n16953) );
  MUX21X1 U8969 ( .IN1(\mem0[49][4] ), .IN2(n794), .S(n7346), .Q(n16952) );
  MUX21X1 U8970 ( .IN1(\mem0[49][3] ), .IN2(n772), .S(n7346), .Q(n16951) );
  MUX21X1 U8971 ( .IN1(\mem0[49][2] ), .IN2(n750), .S(n7346), .Q(n16950) );
  MUX21X1 U8972 ( .IN1(\mem0[49][1] ), .IN2(n728), .S(n7346), .Q(n16949) );
  MUX21X1 U8973 ( .IN1(\mem0[49][0] ), .IN2(n706), .S(n7346), .Q(n16948) );
  AND2X1 U8974 ( .IN1(n7332), .IN2(n7128), .Q(n7346) );
  MUX21X1 U8975 ( .IN1(\mem0[48][7] ), .IN2(n860), .S(n7347), .Q(n16947) );
  MUX21X1 U8976 ( .IN1(\mem0[48][6] ), .IN2(n838), .S(n7347), .Q(n16946) );
  MUX21X1 U8977 ( .IN1(\mem0[48][5] ), .IN2(n816), .S(n7347), .Q(n16945) );
  MUX21X1 U8978 ( .IN1(\mem0[48][4] ), .IN2(n794), .S(n7347), .Q(n16944) );
  MUX21X1 U8979 ( .IN1(\mem0[48][3] ), .IN2(n772), .S(n7347), .Q(n16943) );
  MUX21X1 U8980 ( .IN1(\mem0[48][2] ), .IN2(n750), .S(n7347), .Q(n16942) );
  MUX21X1 U8981 ( .IN1(\mem0[48][1] ), .IN2(n728), .S(n7347), .Q(n16941) );
  MUX21X1 U8982 ( .IN1(\mem0[48][0] ), .IN2(n706), .S(n7347), .Q(n16940) );
  AND2X1 U8983 ( .IN1(n7332), .IN2(n7130), .Q(n7347) );
  AND2X1 U8984 ( .IN1(n7348), .IN2(n7132), .Q(n7332) );
  MUX21X1 U8985 ( .IN1(\mem0[47][7] ), .IN2(n860), .S(n7349), .Q(n16939) );
  MUX21X1 U8986 ( .IN1(\mem0[47][6] ), .IN2(n838), .S(n7349), .Q(n16938) );
  MUX21X1 U8987 ( .IN1(\mem0[47][5] ), .IN2(n816), .S(n7349), .Q(n16937) );
  MUX21X1 U8988 ( .IN1(\mem0[47][4] ), .IN2(n794), .S(n7349), .Q(n16936) );
  MUX21X1 U8989 ( .IN1(\mem0[47][3] ), .IN2(n772), .S(n7349), .Q(n16935) );
  MUX21X1 U8990 ( .IN1(\mem0[47][2] ), .IN2(n750), .S(n7349), .Q(n16934) );
  MUX21X1 U8991 ( .IN1(\mem0[47][1] ), .IN2(n728), .S(n7349), .Q(n16933) );
  MUX21X1 U8992 ( .IN1(\mem0[47][0] ), .IN2(n706), .S(n7349), .Q(n16932) );
  AND2X1 U8993 ( .IN1(n7350), .IN2(n7099), .Q(n7349) );
  MUX21X1 U8994 ( .IN1(\mem0[46][7] ), .IN2(n860), .S(n7351), .Q(n16931) );
  MUX21X1 U8995 ( .IN1(\mem0[46][6] ), .IN2(n838), .S(n7351), .Q(n16930) );
  MUX21X1 U8996 ( .IN1(\mem0[46][5] ), .IN2(n816), .S(n7351), .Q(n16929) );
  MUX21X1 U8997 ( .IN1(\mem0[46][4] ), .IN2(n794), .S(n7351), .Q(n16928) );
  MUX21X1 U8998 ( .IN1(\mem0[46][3] ), .IN2(n772), .S(n7351), .Q(n16927) );
  MUX21X1 U8999 ( .IN1(\mem0[46][2] ), .IN2(n750), .S(n7351), .Q(n16926) );
  MUX21X1 U9000 ( .IN1(\mem0[46][1] ), .IN2(n728), .S(n7351), .Q(n16925) );
  MUX21X1 U9001 ( .IN1(\mem0[46][0] ), .IN2(n706), .S(n7351), .Q(n16924) );
  AND2X1 U9002 ( .IN1(n7350), .IN2(n7102), .Q(n7351) );
  MUX21X1 U9003 ( .IN1(\mem0[45][7] ), .IN2(n860), .S(n7352), .Q(n16923) );
  MUX21X1 U9004 ( .IN1(\mem0[45][6] ), .IN2(n838), .S(n7352), .Q(n16922) );
  MUX21X1 U9005 ( .IN1(\mem0[45][5] ), .IN2(n816), .S(n7352), .Q(n16921) );
  MUX21X1 U9006 ( .IN1(\mem0[45][4] ), .IN2(n794), .S(n7352), .Q(n16920) );
  MUX21X1 U9007 ( .IN1(\mem0[45][3] ), .IN2(n772), .S(n7352), .Q(n16919) );
  MUX21X1 U9008 ( .IN1(\mem0[45][2] ), .IN2(n750), .S(n7352), .Q(n16918) );
  MUX21X1 U9009 ( .IN1(\mem0[45][1] ), .IN2(n728), .S(n7352), .Q(n16917) );
  MUX21X1 U9010 ( .IN1(\mem0[45][0] ), .IN2(n706), .S(n7352), .Q(n16916) );
  AND2X1 U9011 ( .IN1(n7350), .IN2(n7104), .Q(n7352) );
  MUX21X1 U9012 ( .IN1(\mem0[44][7] ), .IN2(n860), .S(n7353), .Q(n16915) );
  MUX21X1 U9013 ( .IN1(\mem0[44][6] ), .IN2(n838), .S(n7353), .Q(n16914) );
  MUX21X1 U9014 ( .IN1(\mem0[44][5] ), .IN2(n816), .S(n7353), .Q(n16913) );
  MUX21X1 U9015 ( .IN1(\mem0[44][4] ), .IN2(n794), .S(n7353), .Q(n16912) );
  MUX21X1 U9016 ( .IN1(\mem0[44][3] ), .IN2(n772), .S(n7353), .Q(n16911) );
  MUX21X1 U9017 ( .IN1(\mem0[44][2] ), .IN2(n750), .S(n7353), .Q(n16910) );
  MUX21X1 U9018 ( .IN1(\mem0[44][1] ), .IN2(n728), .S(n7353), .Q(n16909) );
  MUX21X1 U9019 ( .IN1(\mem0[44][0] ), .IN2(n706), .S(n7353), .Q(n16908) );
  AND2X1 U9020 ( .IN1(n7350), .IN2(n7106), .Q(n7353) );
  MUX21X1 U9021 ( .IN1(\mem0[43][7] ), .IN2(n860), .S(n7354), .Q(n16907) );
  MUX21X1 U9022 ( .IN1(\mem0[43][6] ), .IN2(n838), .S(n7354), .Q(n16906) );
  MUX21X1 U9023 ( .IN1(\mem0[43][5] ), .IN2(n816), .S(n7354), .Q(n16905) );
  MUX21X1 U9024 ( .IN1(\mem0[43][4] ), .IN2(n794), .S(n7354), .Q(n16904) );
  MUX21X1 U9025 ( .IN1(\mem0[43][3] ), .IN2(n772), .S(n7354), .Q(n16903) );
  MUX21X1 U9026 ( .IN1(\mem0[43][2] ), .IN2(n750), .S(n7354), .Q(n16902) );
  MUX21X1 U9027 ( .IN1(\mem0[43][1] ), .IN2(n728), .S(n7354), .Q(n16901) );
  MUX21X1 U9028 ( .IN1(\mem0[43][0] ), .IN2(n706), .S(n7354), .Q(n16900) );
  AND2X1 U9029 ( .IN1(n7350), .IN2(n7108), .Q(n7354) );
  MUX21X1 U9030 ( .IN1(\mem0[42][7] ), .IN2(n860), .S(n7355), .Q(n16899) );
  MUX21X1 U9031 ( .IN1(\mem0[42][6] ), .IN2(n838), .S(n7355), .Q(n16898) );
  MUX21X1 U9032 ( .IN1(\mem0[42][5] ), .IN2(n816), .S(n7355), .Q(n16897) );
  MUX21X1 U9033 ( .IN1(\mem0[42][4] ), .IN2(n794), .S(n7355), .Q(n16896) );
  MUX21X1 U9034 ( .IN1(\mem0[42][3] ), .IN2(n772), .S(n7355), .Q(n16895) );
  MUX21X1 U9035 ( .IN1(\mem0[42][2] ), .IN2(n750), .S(n7355), .Q(n16894) );
  MUX21X1 U9036 ( .IN1(\mem0[42][1] ), .IN2(n728), .S(n7355), .Q(n16893) );
  MUX21X1 U9037 ( .IN1(\mem0[42][0] ), .IN2(n706), .S(n7355), .Q(n16892) );
  AND2X1 U9038 ( .IN1(n7350), .IN2(n7110), .Q(n7355) );
  MUX21X1 U9039 ( .IN1(\mem0[41][7] ), .IN2(n860), .S(n7356), .Q(n16891) );
  MUX21X1 U9040 ( .IN1(\mem0[41][6] ), .IN2(n838), .S(n7356), .Q(n16890) );
  MUX21X1 U9041 ( .IN1(\mem0[41][5] ), .IN2(n816), .S(n7356), .Q(n16889) );
  MUX21X1 U9042 ( .IN1(\mem0[41][4] ), .IN2(n794), .S(n7356), .Q(n16888) );
  MUX21X1 U9043 ( .IN1(\mem0[41][3] ), .IN2(n772), .S(n7356), .Q(n16887) );
  MUX21X1 U9044 ( .IN1(\mem0[41][2] ), .IN2(n750), .S(n7356), .Q(n16886) );
  MUX21X1 U9045 ( .IN1(\mem0[41][1] ), .IN2(n728), .S(n7356), .Q(n16885) );
  MUX21X1 U9046 ( .IN1(\mem0[41][0] ), .IN2(n706), .S(n7356), .Q(n16884) );
  AND2X1 U9047 ( .IN1(n7350), .IN2(n7112), .Q(n7356) );
  MUX21X1 U9048 ( .IN1(\mem0[40][7] ), .IN2(n860), .S(n7357), .Q(n16883) );
  MUX21X1 U9049 ( .IN1(\mem0[40][6] ), .IN2(n838), .S(n7357), .Q(n16882) );
  MUX21X1 U9050 ( .IN1(\mem0[40][5] ), .IN2(n816), .S(n7357), .Q(n16881) );
  MUX21X1 U9051 ( .IN1(\mem0[40][4] ), .IN2(n794), .S(n7357), .Q(n16880) );
  MUX21X1 U9052 ( .IN1(\mem0[40][3] ), .IN2(n772), .S(n7357), .Q(n16879) );
  MUX21X1 U9053 ( .IN1(\mem0[40][2] ), .IN2(n750), .S(n7357), .Q(n16878) );
  MUX21X1 U9054 ( .IN1(\mem0[40][1] ), .IN2(n728), .S(n7357), .Q(n16877) );
  MUX21X1 U9055 ( .IN1(\mem0[40][0] ), .IN2(n706), .S(n7357), .Q(n16876) );
  AND2X1 U9056 ( .IN1(n7350), .IN2(n7114), .Q(n7357) );
  MUX21X1 U9057 ( .IN1(\mem0[39][7] ), .IN2(n861), .S(n7358), .Q(n16875) );
  MUX21X1 U9058 ( .IN1(\mem0[39][6] ), .IN2(n839), .S(n7358), .Q(n16874) );
  MUX21X1 U9059 ( .IN1(\mem0[39][5] ), .IN2(n817), .S(n7358), .Q(n16873) );
  MUX21X1 U9060 ( .IN1(\mem0[39][4] ), .IN2(n795), .S(n7358), .Q(n16872) );
  MUX21X1 U9061 ( .IN1(\mem0[39][3] ), .IN2(n773), .S(n7358), .Q(n16871) );
  MUX21X1 U9062 ( .IN1(\mem0[39][2] ), .IN2(n751), .S(n7358), .Q(n16870) );
  MUX21X1 U9063 ( .IN1(\mem0[39][1] ), .IN2(n729), .S(n7358), .Q(n16869) );
  MUX21X1 U9064 ( .IN1(\mem0[39][0] ), .IN2(n707), .S(n7358), .Q(n16868) );
  AND2X1 U9065 ( .IN1(n7350), .IN2(n7116), .Q(n7358) );
  MUX21X1 U9066 ( .IN1(\mem0[38][7] ), .IN2(n861), .S(n7359), .Q(n16867) );
  MUX21X1 U9067 ( .IN1(\mem0[38][6] ), .IN2(n839), .S(n7359), .Q(n16866) );
  MUX21X1 U9068 ( .IN1(\mem0[38][5] ), .IN2(n817), .S(n7359), .Q(n16865) );
  MUX21X1 U9069 ( .IN1(\mem0[38][4] ), .IN2(n795), .S(n7359), .Q(n16864) );
  MUX21X1 U9070 ( .IN1(\mem0[38][3] ), .IN2(n773), .S(n7359), .Q(n16863) );
  MUX21X1 U9071 ( .IN1(\mem0[38][2] ), .IN2(n751), .S(n7359), .Q(n16862) );
  MUX21X1 U9072 ( .IN1(\mem0[38][1] ), .IN2(n729), .S(n7359), .Q(n16861) );
  MUX21X1 U9073 ( .IN1(\mem0[38][0] ), .IN2(n707), .S(n7359), .Q(n16860) );
  AND2X1 U9074 ( .IN1(n7350), .IN2(n7118), .Q(n7359) );
  MUX21X1 U9075 ( .IN1(\mem0[37][7] ), .IN2(n861), .S(n7360), .Q(n16859) );
  MUX21X1 U9076 ( .IN1(\mem0[37][6] ), .IN2(n839), .S(n7360), .Q(n16858) );
  MUX21X1 U9077 ( .IN1(\mem0[37][5] ), .IN2(n817), .S(n7360), .Q(n16857) );
  MUX21X1 U9078 ( .IN1(\mem0[37][4] ), .IN2(n795), .S(n7360), .Q(n16856) );
  MUX21X1 U9079 ( .IN1(\mem0[37][3] ), .IN2(n773), .S(n7360), .Q(n16855) );
  MUX21X1 U9080 ( .IN1(\mem0[37][2] ), .IN2(n751), .S(n7360), .Q(n16854) );
  MUX21X1 U9081 ( .IN1(\mem0[37][1] ), .IN2(n729), .S(n7360), .Q(n16853) );
  MUX21X1 U9082 ( .IN1(\mem0[37][0] ), .IN2(n707), .S(n7360), .Q(n16852) );
  AND2X1 U9083 ( .IN1(n7350), .IN2(n7120), .Q(n7360) );
  MUX21X1 U9084 ( .IN1(\mem0[36][7] ), .IN2(n861), .S(n7361), .Q(n16851) );
  MUX21X1 U9085 ( .IN1(\mem0[36][6] ), .IN2(n839), .S(n7361), .Q(n16850) );
  MUX21X1 U9086 ( .IN1(\mem0[36][5] ), .IN2(n817), .S(n7361), .Q(n16849) );
  MUX21X1 U9087 ( .IN1(\mem0[36][4] ), .IN2(n795), .S(n7361), .Q(n16848) );
  MUX21X1 U9088 ( .IN1(\mem0[36][3] ), .IN2(n773), .S(n7361), .Q(n16847) );
  MUX21X1 U9089 ( .IN1(\mem0[36][2] ), .IN2(n751), .S(n7361), .Q(n16846) );
  MUX21X1 U9090 ( .IN1(\mem0[36][1] ), .IN2(n729), .S(n7361), .Q(n16845) );
  MUX21X1 U9091 ( .IN1(\mem0[36][0] ), .IN2(n707), .S(n7361), .Q(n16844) );
  AND2X1 U9092 ( .IN1(n7350), .IN2(n7122), .Q(n7361) );
  MUX21X1 U9093 ( .IN1(\mem0[35][7] ), .IN2(n861), .S(n7362), .Q(n16843) );
  MUX21X1 U9094 ( .IN1(\mem0[35][6] ), .IN2(n839), .S(n7362), .Q(n16842) );
  MUX21X1 U9095 ( .IN1(\mem0[35][5] ), .IN2(n817), .S(n7362), .Q(n16841) );
  MUX21X1 U9096 ( .IN1(\mem0[35][4] ), .IN2(n795), .S(n7362), .Q(n16840) );
  MUX21X1 U9097 ( .IN1(\mem0[35][3] ), .IN2(n773), .S(n7362), .Q(n16839) );
  MUX21X1 U9098 ( .IN1(\mem0[35][2] ), .IN2(n751), .S(n7362), .Q(n16838) );
  MUX21X1 U9099 ( .IN1(\mem0[35][1] ), .IN2(n729), .S(n7362), .Q(n16837) );
  MUX21X1 U9100 ( .IN1(\mem0[35][0] ), .IN2(n707), .S(n7362), .Q(n16836) );
  AND2X1 U9101 ( .IN1(n7350), .IN2(n7124), .Q(n7362) );
  MUX21X1 U9102 ( .IN1(\mem0[34][7] ), .IN2(n861), .S(n7363), .Q(n16835) );
  MUX21X1 U9103 ( .IN1(\mem0[34][6] ), .IN2(n839), .S(n7363), .Q(n16834) );
  MUX21X1 U9104 ( .IN1(\mem0[34][5] ), .IN2(n817), .S(n7363), .Q(n16833) );
  MUX21X1 U9105 ( .IN1(\mem0[34][4] ), .IN2(n795), .S(n7363), .Q(n16832) );
  MUX21X1 U9106 ( .IN1(\mem0[34][3] ), .IN2(n773), .S(n7363), .Q(n16831) );
  MUX21X1 U9107 ( .IN1(\mem0[34][2] ), .IN2(n751), .S(n7363), .Q(n16830) );
  MUX21X1 U9108 ( .IN1(\mem0[34][1] ), .IN2(n729), .S(n7363), .Q(n16829) );
  MUX21X1 U9109 ( .IN1(\mem0[34][0] ), .IN2(n707), .S(n7363), .Q(n16828) );
  AND2X1 U9110 ( .IN1(n7350), .IN2(n7126), .Q(n7363) );
  MUX21X1 U9111 ( .IN1(\mem0[33][7] ), .IN2(n861), .S(n7364), .Q(n16827) );
  MUX21X1 U9112 ( .IN1(\mem0[33][6] ), .IN2(n839), .S(n7364), .Q(n16826) );
  MUX21X1 U9113 ( .IN1(\mem0[33][5] ), .IN2(n817), .S(n7364), .Q(n16825) );
  MUX21X1 U9114 ( .IN1(\mem0[33][4] ), .IN2(n795), .S(n7364), .Q(n16824) );
  MUX21X1 U9115 ( .IN1(\mem0[33][3] ), .IN2(n773), .S(n7364), .Q(n16823) );
  MUX21X1 U9116 ( .IN1(\mem0[33][2] ), .IN2(n751), .S(n7364), .Q(n16822) );
  MUX21X1 U9117 ( .IN1(\mem0[33][1] ), .IN2(n729), .S(n7364), .Q(n16821) );
  MUX21X1 U9118 ( .IN1(\mem0[33][0] ), .IN2(n707), .S(n7364), .Q(n16820) );
  AND2X1 U9119 ( .IN1(n7350), .IN2(n7128), .Q(n7364) );
  MUX21X1 U9120 ( .IN1(\mem0[32][7] ), .IN2(n861), .S(n7365), .Q(n16819) );
  MUX21X1 U9121 ( .IN1(\mem0[32][6] ), .IN2(n839), .S(n7365), .Q(n16818) );
  MUX21X1 U9122 ( .IN1(\mem0[32][5] ), .IN2(n817), .S(n7365), .Q(n16817) );
  MUX21X1 U9123 ( .IN1(\mem0[32][4] ), .IN2(n795), .S(n7365), .Q(n16816) );
  MUX21X1 U9124 ( .IN1(\mem0[32][3] ), .IN2(n773), .S(n7365), .Q(n16815) );
  MUX21X1 U9125 ( .IN1(\mem0[32][2] ), .IN2(n751), .S(n7365), .Q(n16814) );
  MUX21X1 U9126 ( .IN1(\mem0[32][1] ), .IN2(n729), .S(n7365), .Q(n16813) );
  MUX21X1 U9127 ( .IN1(\mem0[32][0] ), .IN2(n707), .S(n7365), .Q(n16812) );
  AND2X1 U9128 ( .IN1(n7350), .IN2(n7130), .Q(n7365) );
  AND2X1 U9129 ( .IN1(n7366), .IN2(n7132), .Q(n7350) );
  MUX21X1 U9130 ( .IN1(\mem0[31][7] ), .IN2(n861), .S(n7367), .Q(n16811) );
  MUX21X1 U9131 ( .IN1(\mem0[31][6] ), .IN2(n839), .S(n7367), .Q(n16810) );
  MUX21X1 U9132 ( .IN1(\mem0[31][5] ), .IN2(n817), .S(n7367), .Q(n16809) );
  MUX21X1 U9133 ( .IN1(\mem0[31][4] ), .IN2(n795), .S(n7367), .Q(n16808) );
  MUX21X1 U9134 ( .IN1(\mem0[31][3] ), .IN2(n773), .S(n7367), .Q(n16807) );
  MUX21X1 U9135 ( .IN1(\mem0[31][2] ), .IN2(n751), .S(n7367), .Q(n16806) );
  MUX21X1 U9136 ( .IN1(\mem0[31][1] ), .IN2(n729), .S(n7367), .Q(n16805) );
  MUX21X1 U9137 ( .IN1(\mem0[31][0] ), .IN2(n707), .S(n7367), .Q(n16804) );
  AND2X1 U9138 ( .IN1(n7368), .IN2(n7099), .Q(n7367) );
  MUX21X1 U9139 ( .IN1(\mem0[30][7] ), .IN2(n861), .S(n7369), .Q(n16803) );
  MUX21X1 U9140 ( .IN1(\mem0[30][6] ), .IN2(n839), .S(n7369), .Q(n16802) );
  MUX21X1 U9141 ( .IN1(\mem0[30][5] ), .IN2(n817), .S(n7369), .Q(n16801) );
  MUX21X1 U9142 ( .IN1(\mem0[30][4] ), .IN2(n795), .S(n7369), .Q(n16800) );
  MUX21X1 U9143 ( .IN1(\mem0[30][3] ), .IN2(n773), .S(n7369), .Q(n16799) );
  MUX21X1 U9144 ( .IN1(\mem0[30][2] ), .IN2(n751), .S(n7369), .Q(n16798) );
  MUX21X1 U9145 ( .IN1(\mem0[30][1] ), .IN2(n729), .S(n7369), .Q(n16797) );
  MUX21X1 U9146 ( .IN1(\mem0[30][0] ), .IN2(n707), .S(n7369), .Q(n16796) );
  AND2X1 U9147 ( .IN1(n7368), .IN2(n7102), .Q(n7369) );
  MUX21X1 U9148 ( .IN1(\mem0[29][7] ), .IN2(n861), .S(n7370), .Q(n16795) );
  MUX21X1 U9149 ( .IN1(\mem0[29][6] ), .IN2(n839), .S(n7370), .Q(n16794) );
  MUX21X1 U9150 ( .IN1(\mem0[29][5] ), .IN2(n817), .S(n7370), .Q(n16793) );
  MUX21X1 U9151 ( .IN1(\mem0[29][4] ), .IN2(n795), .S(n7370), .Q(n16792) );
  MUX21X1 U9152 ( .IN1(\mem0[29][3] ), .IN2(n773), .S(n7370), .Q(n16791) );
  MUX21X1 U9153 ( .IN1(\mem0[29][2] ), .IN2(n751), .S(n7370), .Q(n16790) );
  MUX21X1 U9154 ( .IN1(\mem0[29][1] ), .IN2(n729), .S(n7370), .Q(n16789) );
  MUX21X1 U9155 ( .IN1(\mem0[29][0] ), .IN2(n707), .S(n7370), .Q(n16788) );
  AND2X1 U9156 ( .IN1(n7368), .IN2(n7104), .Q(n7370) );
  MUX21X1 U9157 ( .IN1(\mem0[28][7] ), .IN2(n861), .S(n7371), .Q(n16787) );
  MUX21X1 U9158 ( .IN1(\mem0[28][6] ), .IN2(n839), .S(n7371), .Q(n16786) );
  MUX21X1 U9159 ( .IN1(\mem0[28][5] ), .IN2(n817), .S(n7371), .Q(n16785) );
  MUX21X1 U9160 ( .IN1(\mem0[28][4] ), .IN2(n795), .S(n7371), .Q(n16784) );
  MUX21X1 U9161 ( .IN1(\mem0[28][3] ), .IN2(n773), .S(n7371), .Q(n16783) );
  MUX21X1 U9162 ( .IN1(\mem0[28][2] ), .IN2(n751), .S(n7371), .Q(n16782) );
  MUX21X1 U9163 ( .IN1(\mem0[28][1] ), .IN2(n729), .S(n7371), .Q(n16781) );
  MUX21X1 U9164 ( .IN1(\mem0[28][0] ), .IN2(n707), .S(n7371), .Q(n16780) );
  AND2X1 U9165 ( .IN1(n7368), .IN2(n7106), .Q(n7371) );
  MUX21X1 U9166 ( .IN1(\mem0[27][7] ), .IN2(n862), .S(n7372), .Q(n16779) );
  MUX21X1 U9167 ( .IN1(\mem0[27][6] ), .IN2(n840), .S(n7372), .Q(n16778) );
  MUX21X1 U9168 ( .IN1(\mem0[27][5] ), .IN2(n818), .S(n7372), .Q(n16777) );
  MUX21X1 U9169 ( .IN1(\mem0[27][4] ), .IN2(n796), .S(n7372), .Q(n16776) );
  MUX21X1 U9170 ( .IN1(\mem0[27][3] ), .IN2(n774), .S(n7372), .Q(n16775) );
  MUX21X1 U9171 ( .IN1(\mem0[27][2] ), .IN2(n752), .S(n7372), .Q(n16774) );
  MUX21X1 U9172 ( .IN1(\mem0[27][1] ), .IN2(n730), .S(n7372), .Q(n16773) );
  MUX21X1 U9173 ( .IN1(\mem0[27][0] ), .IN2(n708), .S(n7372), .Q(n16772) );
  AND2X1 U9174 ( .IN1(n7368), .IN2(n7108), .Q(n7372) );
  MUX21X1 U9175 ( .IN1(\mem0[26][7] ), .IN2(n862), .S(n7373), .Q(n16771) );
  MUX21X1 U9176 ( .IN1(\mem0[26][6] ), .IN2(n840), .S(n7373), .Q(n16770) );
  MUX21X1 U9177 ( .IN1(\mem0[26][5] ), .IN2(n818), .S(n7373), .Q(n16769) );
  MUX21X1 U9178 ( .IN1(\mem0[26][4] ), .IN2(n796), .S(n7373), .Q(n16768) );
  MUX21X1 U9179 ( .IN1(\mem0[26][3] ), .IN2(n774), .S(n7373), .Q(n16767) );
  MUX21X1 U9180 ( .IN1(\mem0[26][2] ), .IN2(n752), .S(n7373), .Q(n16766) );
  MUX21X1 U9181 ( .IN1(\mem0[26][1] ), .IN2(n730), .S(n7373), .Q(n16765) );
  MUX21X1 U9182 ( .IN1(\mem0[26][0] ), .IN2(n708), .S(n7373), .Q(n16764) );
  AND2X1 U9183 ( .IN1(n7368), .IN2(n7110), .Q(n7373) );
  MUX21X1 U9184 ( .IN1(\mem0[25][7] ), .IN2(n862), .S(n7374), .Q(n16763) );
  MUX21X1 U9185 ( .IN1(\mem0[25][6] ), .IN2(n840), .S(n7374), .Q(n16762) );
  MUX21X1 U9186 ( .IN1(\mem0[25][5] ), .IN2(n818), .S(n7374), .Q(n16761) );
  MUX21X1 U9187 ( .IN1(\mem0[25][4] ), .IN2(n796), .S(n7374), .Q(n16760) );
  MUX21X1 U9188 ( .IN1(\mem0[25][3] ), .IN2(n774), .S(n7374), .Q(n16759) );
  MUX21X1 U9189 ( .IN1(\mem0[25][2] ), .IN2(n752), .S(n7374), .Q(n16758) );
  MUX21X1 U9190 ( .IN1(\mem0[25][1] ), .IN2(n730), .S(n7374), .Q(n16757) );
  MUX21X1 U9191 ( .IN1(\mem0[25][0] ), .IN2(n708), .S(n7374), .Q(n16756) );
  AND2X1 U9192 ( .IN1(n7368), .IN2(n7112), .Q(n7374) );
  MUX21X1 U9193 ( .IN1(\mem0[24][7] ), .IN2(n862), .S(n7375), .Q(n16755) );
  MUX21X1 U9194 ( .IN1(\mem0[24][6] ), .IN2(n840), .S(n7375), .Q(n16754) );
  MUX21X1 U9195 ( .IN1(\mem0[24][5] ), .IN2(n818), .S(n7375), .Q(n16753) );
  MUX21X1 U9196 ( .IN1(\mem0[24][4] ), .IN2(n796), .S(n7375), .Q(n16752) );
  MUX21X1 U9197 ( .IN1(\mem0[24][3] ), .IN2(n774), .S(n7375), .Q(n16751) );
  MUX21X1 U9198 ( .IN1(\mem0[24][2] ), .IN2(n752), .S(n7375), .Q(n16750) );
  MUX21X1 U9199 ( .IN1(\mem0[24][1] ), .IN2(n730), .S(n7375), .Q(n16749) );
  MUX21X1 U9200 ( .IN1(\mem0[24][0] ), .IN2(n708), .S(n7375), .Q(n16748) );
  AND2X1 U9201 ( .IN1(n7368), .IN2(n7114), .Q(n7375) );
  MUX21X1 U9202 ( .IN1(\mem0[23][7] ), .IN2(n862), .S(n7376), .Q(n16747) );
  MUX21X1 U9203 ( .IN1(\mem0[23][6] ), .IN2(n840), .S(n7376), .Q(n16746) );
  MUX21X1 U9204 ( .IN1(\mem0[23][5] ), .IN2(n818), .S(n7376), .Q(n16745) );
  MUX21X1 U9205 ( .IN1(\mem0[23][4] ), .IN2(n796), .S(n7376), .Q(n16744) );
  MUX21X1 U9206 ( .IN1(\mem0[23][3] ), .IN2(n774), .S(n7376), .Q(n16743) );
  MUX21X1 U9207 ( .IN1(\mem0[23][2] ), .IN2(n752), .S(n7376), .Q(n16742) );
  MUX21X1 U9208 ( .IN1(\mem0[23][1] ), .IN2(n730), .S(n7376), .Q(n16741) );
  MUX21X1 U9209 ( .IN1(\mem0[23][0] ), .IN2(n708), .S(n7376), .Q(n16740) );
  AND2X1 U9210 ( .IN1(n7368), .IN2(n7116), .Q(n7376) );
  MUX21X1 U9211 ( .IN1(\mem0[22][7] ), .IN2(n862), .S(n7377), .Q(n16739) );
  MUX21X1 U9212 ( .IN1(\mem0[22][6] ), .IN2(n840), .S(n7377), .Q(n16738) );
  MUX21X1 U9213 ( .IN1(\mem0[22][5] ), .IN2(n818), .S(n7377), .Q(n16737) );
  MUX21X1 U9214 ( .IN1(\mem0[22][4] ), .IN2(n796), .S(n7377), .Q(n16736) );
  MUX21X1 U9215 ( .IN1(\mem0[22][3] ), .IN2(n774), .S(n7377), .Q(n16735) );
  MUX21X1 U9216 ( .IN1(\mem0[22][2] ), .IN2(n752), .S(n7377), .Q(n16734) );
  MUX21X1 U9217 ( .IN1(\mem0[22][1] ), .IN2(n730), .S(n7377), .Q(n16733) );
  MUX21X1 U9218 ( .IN1(\mem0[22][0] ), .IN2(n708), .S(n7377), .Q(n16732) );
  AND2X1 U9219 ( .IN1(n7368), .IN2(n7118), .Q(n7377) );
  MUX21X1 U9220 ( .IN1(\mem0[21][7] ), .IN2(n862), .S(n7378), .Q(n16731) );
  MUX21X1 U9221 ( .IN1(\mem0[21][6] ), .IN2(n840), .S(n7378), .Q(n16730) );
  MUX21X1 U9222 ( .IN1(\mem0[21][5] ), .IN2(n818), .S(n7378), .Q(n16729) );
  MUX21X1 U9223 ( .IN1(\mem0[21][4] ), .IN2(n796), .S(n7378), .Q(n16728) );
  MUX21X1 U9224 ( .IN1(\mem0[21][3] ), .IN2(n774), .S(n7378), .Q(n16727) );
  MUX21X1 U9225 ( .IN1(\mem0[21][2] ), .IN2(n752), .S(n7378), .Q(n16726) );
  MUX21X1 U9226 ( .IN1(\mem0[21][1] ), .IN2(n730), .S(n7378), .Q(n16725) );
  MUX21X1 U9227 ( .IN1(\mem0[21][0] ), .IN2(n708), .S(n7378), .Q(n16724) );
  AND2X1 U9228 ( .IN1(n7368), .IN2(n7120), .Q(n7378) );
  MUX21X1 U9229 ( .IN1(\mem0[20][7] ), .IN2(n862), .S(n7379), .Q(n16723) );
  MUX21X1 U9230 ( .IN1(\mem0[20][6] ), .IN2(n840), .S(n7379), .Q(n16722) );
  MUX21X1 U9231 ( .IN1(\mem0[20][5] ), .IN2(n818), .S(n7379), .Q(n16721) );
  MUX21X1 U9232 ( .IN1(\mem0[20][4] ), .IN2(n796), .S(n7379), .Q(n16720) );
  MUX21X1 U9233 ( .IN1(\mem0[20][3] ), .IN2(n774), .S(n7379), .Q(n16719) );
  MUX21X1 U9234 ( .IN1(\mem0[20][2] ), .IN2(n752), .S(n7379), .Q(n16718) );
  MUX21X1 U9235 ( .IN1(\mem0[20][1] ), .IN2(n730), .S(n7379), .Q(n16717) );
  MUX21X1 U9236 ( .IN1(\mem0[20][0] ), .IN2(n708), .S(n7379), .Q(n16716) );
  AND2X1 U9237 ( .IN1(n7368), .IN2(n7122), .Q(n7379) );
  MUX21X1 U9238 ( .IN1(\mem0[19][7] ), .IN2(n862), .S(n7380), .Q(n16715) );
  MUX21X1 U9239 ( .IN1(\mem0[19][6] ), .IN2(n840), .S(n7380), .Q(n16714) );
  MUX21X1 U9240 ( .IN1(\mem0[19][5] ), .IN2(n818), .S(n7380), .Q(n16713) );
  MUX21X1 U9241 ( .IN1(\mem0[19][4] ), .IN2(n796), .S(n7380), .Q(n16712) );
  MUX21X1 U9242 ( .IN1(\mem0[19][3] ), .IN2(n774), .S(n7380), .Q(n16711) );
  MUX21X1 U9243 ( .IN1(\mem0[19][2] ), .IN2(n752), .S(n7380), .Q(n16710) );
  MUX21X1 U9244 ( .IN1(\mem0[19][1] ), .IN2(n730), .S(n7380), .Q(n16709) );
  MUX21X1 U9245 ( .IN1(\mem0[19][0] ), .IN2(n708), .S(n7380), .Q(n16708) );
  AND2X1 U9246 ( .IN1(n7368), .IN2(n7124), .Q(n7380) );
  MUX21X1 U9247 ( .IN1(\mem0[18][7] ), .IN2(n862), .S(n7381), .Q(n16707) );
  MUX21X1 U9248 ( .IN1(\mem0[18][6] ), .IN2(n840), .S(n7381), .Q(n16706) );
  MUX21X1 U9249 ( .IN1(\mem0[18][5] ), .IN2(n818), .S(n7381), .Q(n16705) );
  MUX21X1 U9250 ( .IN1(\mem0[18][4] ), .IN2(n796), .S(n7381), .Q(n16704) );
  MUX21X1 U9251 ( .IN1(\mem0[18][3] ), .IN2(n774), .S(n7381), .Q(n16703) );
  MUX21X1 U9252 ( .IN1(\mem0[18][2] ), .IN2(n752), .S(n7381), .Q(n16702) );
  MUX21X1 U9253 ( .IN1(\mem0[18][1] ), .IN2(n730), .S(n7381), .Q(n16701) );
  MUX21X1 U9254 ( .IN1(\mem0[18][0] ), .IN2(n708), .S(n7381), .Q(n16700) );
  AND2X1 U9255 ( .IN1(n7368), .IN2(n7126), .Q(n7381) );
  MUX21X1 U9256 ( .IN1(\mem0[17][7] ), .IN2(n862), .S(n7382), .Q(n16699) );
  MUX21X1 U9257 ( .IN1(\mem0[17][6] ), .IN2(n840), .S(n7382), .Q(n16698) );
  MUX21X1 U9258 ( .IN1(\mem0[17][5] ), .IN2(n818), .S(n7382), .Q(n16697) );
  MUX21X1 U9259 ( .IN1(\mem0[17][4] ), .IN2(n796), .S(n7382), .Q(n16696) );
  MUX21X1 U9260 ( .IN1(\mem0[17][3] ), .IN2(n774), .S(n7382), .Q(n16695) );
  MUX21X1 U9261 ( .IN1(\mem0[17][2] ), .IN2(n752), .S(n7382), .Q(n16694) );
  MUX21X1 U9262 ( .IN1(\mem0[17][1] ), .IN2(n730), .S(n7382), .Q(n16693) );
  MUX21X1 U9263 ( .IN1(\mem0[17][0] ), .IN2(n708), .S(n7382), .Q(n16692) );
  AND2X1 U9264 ( .IN1(n7368), .IN2(n7128), .Q(n7382) );
  MUX21X1 U9265 ( .IN1(\mem0[16][7] ), .IN2(n862), .S(n7383), .Q(n16691) );
  MUX21X1 U9266 ( .IN1(\mem0[16][6] ), .IN2(n840), .S(n7383), .Q(n16690) );
  MUX21X1 U9267 ( .IN1(\mem0[16][5] ), .IN2(n818), .S(n7383), .Q(n16689) );
  MUX21X1 U9268 ( .IN1(\mem0[16][4] ), .IN2(n796), .S(n7383), .Q(n16688) );
  MUX21X1 U9269 ( .IN1(\mem0[16][3] ), .IN2(n774), .S(n7383), .Q(n16687) );
  MUX21X1 U9270 ( .IN1(\mem0[16][2] ), .IN2(n752), .S(n7383), .Q(n16686) );
  MUX21X1 U9271 ( .IN1(\mem0[16][1] ), .IN2(n730), .S(n7383), .Q(n16685) );
  MUX21X1 U9272 ( .IN1(\mem0[16][0] ), .IN2(n708), .S(n7383), .Q(n16684) );
  AND2X1 U9273 ( .IN1(n7368), .IN2(n7130), .Q(n7383) );
  AND2X1 U9274 ( .IN1(n7384), .IN2(n7132), .Q(n7368) );
  MUX21X1 U9275 ( .IN1(\mem0[15][7] ), .IN2(n863), .S(n7385), .Q(n16683) );
  MUX21X1 U9276 ( .IN1(\mem0[15][6] ), .IN2(n841), .S(n7385), .Q(n16682) );
  MUX21X1 U9277 ( .IN1(\mem0[15][5] ), .IN2(n819), .S(n7385), .Q(n16681) );
  MUX21X1 U9278 ( .IN1(\mem0[15][4] ), .IN2(n797), .S(n7385), .Q(n16680) );
  MUX21X1 U9279 ( .IN1(\mem0[15][3] ), .IN2(n775), .S(n7385), .Q(n16679) );
  MUX21X1 U9280 ( .IN1(\mem0[15][2] ), .IN2(n753), .S(n7385), .Q(n16678) );
  MUX21X1 U9281 ( .IN1(\mem0[15][1] ), .IN2(n731), .S(n7385), .Q(n16677) );
  MUX21X1 U9282 ( .IN1(\mem0[15][0] ), .IN2(n709), .S(n7385), .Q(n16676) );
  AND2X1 U9283 ( .IN1(n7386), .IN2(n7099), .Q(n7385) );
  MUX21X1 U9284 ( .IN1(\mem0[14][7] ), .IN2(n863), .S(n7387), .Q(n16675) );
  MUX21X1 U9285 ( .IN1(\mem0[14][6] ), .IN2(n841), .S(n7387), .Q(n16674) );
  MUX21X1 U9286 ( .IN1(\mem0[14][5] ), .IN2(n819), .S(n7387), .Q(n16673) );
  MUX21X1 U9287 ( .IN1(\mem0[14][4] ), .IN2(n797), .S(n7387), .Q(n16672) );
  MUX21X1 U9288 ( .IN1(\mem0[14][3] ), .IN2(n775), .S(n7387), .Q(n16671) );
  MUX21X1 U9289 ( .IN1(\mem0[14][2] ), .IN2(n753), .S(n7387), .Q(n16670) );
  MUX21X1 U9290 ( .IN1(\mem0[14][1] ), .IN2(n731), .S(n7387), .Q(n16669) );
  MUX21X1 U9291 ( .IN1(\mem0[14][0] ), .IN2(n709), .S(n7387), .Q(n16668) );
  AND2X1 U9292 ( .IN1(n7386), .IN2(n7102), .Q(n7387) );
  MUX21X1 U9293 ( .IN1(\mem0[13][7] ), .IN2(n863), .S(n7388), .Q(n16667) );
  MUX21X1 U9294 ( .IN1(\mem0[13][6] ), .IN2(n841), .S(n7388), .Q(n16666) );
  MUX21X1 U9295 ( .IN1(\mem0[13][5] ), .IN2(n819), .S(n7388), .Q(n16665) );
  MUX21X1 U9296 ( .IN1(\mem0[13][4] ), .IN2(n797), .S(n7388), .Q(n16664) );
  MUX21X1 U9297 ( .IN1(\mem0[13][3] ), .IN2(n775), .S(n7388), .Q(n16663) );
  MUX21X1 U9298 ( .IN1(\mem0[13][2] ), .IN2(n753), .S(n7388), .Q(n16662) );
  MUX21X1 U9299 ( .IN1(\mem0[13][1] ), .IN2(n731), .S(n7388), .Q(n16661) );
  MUX21X1 U9300 ( .IN1(\mem0[13][0] ), .IN2(n709), .S(n7388), .Q(n16660) );
  AND2X1 U9301 ( .IN1(n7386), .IN2(n7104), .Q(n7388) );
  MUX21X1 U9302 ( .IN1(\mem0[12][7] ), .IN2(n863), .S(n7389), .Q(n16659) );
  MUX21X1 U9303 ( .IN1(\mem0[12][6] ), .IN2(n841), .S(n7389), .Q(n16658) );
  MUX21X1 U9304 ( .IN1(\mem0[12][5] ), .IN2(n819), .S(n7389), .Q(n16657) );
  MUX21X1 U9305 ( .IN1(\mem0[12][4] ), .IN2(n797), .S(n7389), .Q(n16656) );
  MUX21X1 U9306 ( .IN1(\mem0[12][3] ), .IN2(n775), .S(n7389), .Q(n16655) );
  MUX21X1 U9307 ( .IN1(\mem0[12][2] ), .IN2(n753), .S(n7389), .Q(n16654) );
  MUX21X1 U9308 ( .IN1(\mem0[12][1] ), .IN2(n731), .S(n7389), .Q(n16653) );
  MUX21X1 U9309 ( .IN1(\mem0[12][0] ), .IN2(n709), .S(n7389), .Q(n16652) );
  AND2X1 U9310 ( .IN1(n7386), .IN2(n7106), .Q(n7389) );
  MUX21X1 U9311 ( .IN1(\mem0[11][7] ), .IN2(n863), .S(n7390), .Q(n16651) );
  MUX21X1 U9312 ( .IN1(\mem0[11][6] ), .IN2(n841), .S(n7390), .Q(n16650) );
  MUX21X1 U9313 ( .IN1(\mem0[11][5] ), .IN2(n819), .S(n7390), .Q(n16649) );
  MUX21X1 U9314 ( .IN1(\mem0[11][4] ), .IN2(n797), .S(n7390), .Q(n16648) );
  MUX21X1 U9315 ( .IN1(\mem0[11][3] ), .IN2(n775), .S(n7390), .Q(n16647) );
  MUX21X1 U9316 ( .IN1(\mem0[11][2] ), .IN2(n753), .S(n7390), .Q(n16646) );
  MUX21X1 U9317 ( .IN1(\mem0[11][1] ), .IN2(n731), .S(n7390), .Q(n16645) );
  MUX21X1 U9318 ( .IN1(\mem0[11][0] ), .IN2(n709), .S(n7390), .Q(n16644) );
  AND2X1 U9319 ( .IN1(n7386), .IN2(n7108), .Q(n7390) );
  MUX21X1 U9320 ( .IN1(\mem0[10][7] ), .IN2(n863), .S(n7391), .Q(n16643) );
  MUX21X1 U9321 ( .IN1(\mem0[10][6] ), .IN2(n841), .S(n7391), .Q(n16642) );
  MUX21X1 U9322 ( .IN1(\mem0[10][5] ), .IN2(n819), .S(n7391), .Q(n16641) );
  MUX21X1 U9323 ( .IN1(\mem0[10][4] ), .IN2(n797), .S(n7391), .Q(n16640) );
  MUX21X1 U9324 ( .IN1(\mem0[10][3] ), .IN2(n775), .S(n7391), .Q(n16639) );
  MUX21X1 U9325 ( .IN1(\mem0[10][2] ), .IN2(n753), .S(n7391), .Q(n16638) );
  MUX21X1 U9326 ( .IN1(\mem0[10][1] ), .IN2(n731), .S(n7391), .Q(n16637) );
  MUX21X1 U9327 ( .IN1(\mem0[10][0] ), .IN2(n709), .S(n7391), .Q(n16636) );
  AND2X1 U9328 ( .IN1(n7386), .IN2(n7110), .Q(n7391) );
  MUX21X1 U9329 ( .IN1(\mem0[9][7] ), .IN2(n863), .S(n7392), .Q(n16635) );
  MUX21X1 U9330 ( .IN1(\mem0[9][6] ), .IN2(n841), .S(n7392), .Q(n16634) );
  MUX21X1 U9331 ( .IN1(\mem0[9][5] ), .IN2(n819), .S(n7392), .Q(n16633) );
  MUX21X1 U9332 ( .IN1(\mem0[9][4] ), .IN2(n797), .S(n7392), .Q(n16632) );
  MUX21X1 U9333 ( .IN1(\mem0[9][3] ), .IN2(n775), .S(n7392), .Q(n16631) );
  MUX21X1 U9334 ( .IN1(\mem0[9][2] ), .IN2(n753), .S(n7392), .Q(n16630) );
  MUX21X1 U9335 ( .IN1(\mem0[9][1] ), .IN2(n731), .S(n7392), .Q(n16629) );
  MUX21X1 U9336 ( .IN1(\mem0[9][0] ), .IN2(n709), .S(n7392), .Q(n16628) );
  AND2X1 U9337 ( .IN1(n7386), .IN2(n7112), .Q(n7392) );
  MUX21X1 U9338 ( .IN1(\mem0[8][7] ), .IN2(n863), .S(n7393), .Q(n16627) );
  MUX21X1 U9339 ( .IN1(\mem0[8][6] ), .IN2(n841), .S(n7393), .Q(n16626) );
  MUX21X1 U9340 ( .IN1(\mem0[8][5] ), .IN2(n819), .S(n7393), .Q(n16625) );
  MUX21X1 U9341 ( .IN1(\mem0[8][4] ), .IN2(n797), .S(n7393), .Q(n16624) );
  MUX21X1 U9342 ( .IN1(\mem0[8][3] ), .IN2(n775), .S(n7393), .Q(n16623) );
  MUX21X1 U9343 ( .IN1(\mem0[8][2] ), .IN2(n753), .S(n7393), .Q(n16622) );
  MUX21X1 U9344 ( .IN1(\mem0[8][1] ), .IN2(n731), .S(n7393), .Q(n16621) );
  MUX21X1 U9345 ( .IN1(\mem0[8][0] ), .IN2(n709), .S(n7393), .Q(n16620) );
  AND2X1 U9346 ( .IN1(n7386), .IN2(n7114), .Q(n7393) );
  MUX21X1 U9347 ( .IN1(\mem0[7][7] ), .IN2(n863), .S(n7394), .Q(n16619) );
  MUX21X1 U9348 ( .IN1(\mem0[7][6] ), .IN2(n841), .S(n7394), .Q(n16618) );
  MUX21X1 U9349 ( .IN1(\mem0[7][5] ), .IN2(n819), .S(n7394), .Q(n16617) );
  MUX21X1 U9350 ( .IN1(\mem0[7][4] ), .IN2(n797), .S(n7394), .Q(n16616) );
  MUX21X1 U9351 ( .IN1(\mem0[7][3] ), .IN2(n775), .S(n7394), .Q(n16615) );
  MUX21X1 U9352 ( .IN1(\mem0[7][2] ), .IN2(n753), .S(n7394), .Q(n16614) );
  MUX21X1 U9353 ( .IN1(\mem0[7][1] ), .IN2(n731), .S(n7394), .Q(n16613) );
  MUX21X1 U9354 ( .IN1(\mem0[7][0] ), .IN2(n709), .S(n7394), .Q(n16612) );
  AND2X1 U9355 ( .IN1(n7386), .IN2(n7116), .Q(n7394) );
  MUX21X1 U9356 ( .IN1(\mem0[6][7] ), .IN2(n863), .S(n7395), .Q(n16611) );
  MUX21X1 U9357 ( .IN1(\mem0[6][6] ), .IN2(n841), .S(n7395), .Q(n16610) );
  MUX21X1 U9358 ( .IN1(\mem0[6][5] ), .IN2(n819), .S(n7395), .Q(n16609) );
  MUX21X1 U9359 ( .IN1(\mem0[6][4] ), .IN2(n797), .S(n7395), .Q(n16608) );
  MUX21X1 U9360 ( .IN1(\mem0[6][3] ), .IN2(n775), .S(n7395), .Q(n16607) );
  MUX21X1 U9361 ( .IN1(\mem0[6][2] ), .IN2(n753), .S(n7395), .Q(n16606) );
  MUX21X1 U9362 ( .IN1(\mem0[6][1] ), .IN2(n731), .S(n7395), .Q(n16605) );
  MUX21X1 U9363 ( .IN1(\mem0[6][0] ), .IN2(n709), .S(n7395), .Q(n16604) );
  AND2X1 U9364 ( .IN1(n7386), .IN2(n7118), .Q(n7395) );
  MUX21X1 U9365 ( .IN1(\mem0[5][7] ), .IN2(n863), .S(n7396), .Q(n16603) );
  MUX21X1 U9366 ( .IN1(\mem0[5][6] ), .IN2(n841), .S(n7396), .Q(n16602) );
  MUX21X1 U9367 ( .IN1(\mem0[5][5] ), .IN2(n819), .S(n7396), .Q(n16601) );
  MUX21X1 U9368 ( .IN1(\mem0[5][4] ), .IN2(n797), .S(n7396), .Q(n16600) );
  MUX21X1 U9369 ( .IN1(\mem0[5][3] ), .IN2(n775), .S(n7396), .Q(n16599) );
  MUX21X1 U9370 ( .IN1(\mem0[5][2] ), .IN2(n753), .S(n7396), .Q(n16598) );
  MUX21X1 U9371 ( .IN1(\mem0[5][1] ), .IN2(n731), .S(n7396), .Q(n16597) );
  MUX21X1 U9372 ( .IN1(\mem0[5][0] ), .IN2(n709), .S(n7396), .Q(n16596) );
  AND2X1 U9373 ( .IN1(n7386), .IN2(n7120), .Q(n7396) );
  MUX21X1 U9374 ( .IN1(\mem0[4][7] ), .IN2(n863), .S(n7397), .Q(n16595) );
  MUX21X1 U9375 ( .IN1(\mem0[4][6] ), .IN2(n841), .S(n7397), .Q(n16594) );
  MUX21X1 U9376 ( .IN1(\mem0[4][5] ), .IN2(n819), .S(n7397), .Q(n16593) );
  MUX21X1 U9377 ( .IN1(\mem0[4][4] ), .IN2(n797), .S(n7397), .Q(n16592) );
  MUX21X1 U9378 ( .IN1(\mem0[4][3] ), .IN2(n775), .S(n7397), .Q(n16591) );
  MUX21X1 U9379 ( .IN1(\mem0[4][2] ), .IN2(n753), .S(n7397), .Q(n16590) );
  MUX21X1 U9380 ( .IN1(\mem0[4][1] ), .IN2(n731), .S(n7397), .Q(n16589) );
  MUX21X1 U9381 ( .IN1(\mem0[4][0] ), .IN2(n709), .S(n7397), .Q(n16588) );
  AND2X1 U9382 ( .IN1(n7386), .IN2(n7122), .Q(n7397) );
  MUX21X1 U9383 ( .IN1(\mem0[3][7] ), .IN2(n864), .S(n7398), .Q(n16587) );
  MUX21X1 U9384 ( .IN1(\mem0[3][6] ), .IN2(n842), .S(n7398), .Q(n16586) );
  MUX21X1 U9385 ( .IN1(\mem0[3][5] ), .IN2(n820), .S(n7398), .Q(n16585) );
  MUX21X1 U9386 ( .IN1(\mem0[3][4] ), .IN2(n798), .S(n7398), .Q(n16584) );
  MUX21X1 U9387 ( .IN1(\mem0[3][3] ), .IN2(n776), .S(n7398), .Q(n16583) );
  MUX21X1 U9388 ( .IN1(\mem0[3][2] ), .IN2(n754), .S(n7398), .Q(n16582) );
  MUX21X1 U9389 ( .IN1(\mem0[3][1] ), .IN2(n732), .S(n7398), .Q(n16581) );
  MUX21X1 U9390 ( .IN1(\mem0[3][0] ), .IN2(n710), .S(n7398), .Q(n16580) );
  AND2X1 U9391 ( .IN1(n7386), .IN2(n7124), .Q(n7398) );
  MUX21X1 U9392 ( .IN1(\mem0[2][7] ), .IN2(n864), .S(n7399), .Q(n16579) );
  MUX21X1 U9393 ( .IN1(\mem0[2][6] ), .IN2(n842), .S(n7399), .Q(n16578) );
  MUX21X1 U9394 ( .IN1(\mem0[2][5] ), .IN2(n820), .S(n7399), .Q(n16577) );
  MUX21X1 U9395 ( .IN1(\mem0[2][4] ), .IN2(n798), .S(n7399), .Q(n16576) );
  MUX21X1 U9396 ( .IN1(\mem0[2][3] ), .IN2(n776), .S(n7399), .Q(n16575) );
  MUX21X1 U9397 ( .IN1(\mem0[2][2] ), .IN2(n754), .S(n7399), .Q(n16574) );
  MUX21X1 U9398 ( .IN1(\mem0[2][1] ), .IN2(n732), .S(n7399), .Q(n16573) );
  MUX21X1 U9399 ( .IN1(\mem0[2][0] ), .IN2(n710), .S(n7399), .Q(n16572) );
  AND2X1 U9400 ( .IN1(n7386), .IN2(n7126), .Q(n7399) );
  MUX21X1 U9401 ( .IN1(\mem0[1][7] ), .IN2(n864), .S(n7400), .Q(n16571) );
  MUX21X1 U9402 ( .IN1(\mem0[1][6] ), .IN2(n842), .S(n7400), .Q(n16570) );
  MUX21X1 U9403 ( .IN1(\mem0[1][5] ), .IN2(n820), .S(n7400), .Q(n16569) );
  MUX21X1 U9404 ( .IN1(\mem0[1][4] ), .IN2(n798), .S(n7400), .Q(n16568) );
  MUX21X1 U9405 ( .IN1(\mem0[1][3] ), .IN2(n776), .S(n7400), .Q(n16567) );
  MUX21X1 U9406 ( .IN1(\mem0[1][2] ), .IN2(n754), .S(n7400), .Q(n16566) );
  MUX21X1 U9407 ( .IN1(\mem0[1][1] ), .IN2(n732), .S(n7400), .Q(n16565) );
  MUX21X1 U9408 ( .IN1(\mem0[1][0] ), .IN2(n710), .S(n7400), .Q(n16564) );
  AND2X1 U9409 ( .IN1(n7386), .IN2(n7128), .Q(n7400) );
  MUX21X1 U9410 ( .IN1(\mem0[0][7] ), .IN2(n864), .S(n7401), .Q(n16563) );
  MUX21X1 U9411 ( .IN1(\mem0[0][6] ), .IN2(n842), .S(n7401), .Q(n16562) );
  MUX21X1 U9412 ( .IN1(\mem0[0][5] ), .IN2(n820), .S(n7401), .Q(n16561) );
  MUX21X1 U9413 ( .IN1(\mem0[0][4] ), .IN2(n798), .S(n7401), .Q(n16560) );
  MUX21X1 U9414 ( .IN1(\mem0[0][3] ), .IN2(n776), .S(n7401), .Q(n16559) );
  MUX21X1 U9415 ( .IN1(\mem0[0][2] ), .IN2(n754), .S(n7401), .Q(n16558) );
  MUX21X1 U9416 ( .IN1(\mem0[0][1] ), .IN2(n732), .S(n7401), .Q(n16557) );
  MUX21X1 U9417 ( .IN1(\mem0[0][0] ), .IN2(n710), .S(n7401), .Q(n16556) );
  AND2X1 U9418 ( .IN1(n7386), .IN2(n7130), .Q(n7401) );
  AND2X1 U9419 ( .IN1(n7402), .IN2(n7132), .Q(n7386) );
  AND2X1 U9420 ( .IN1(we[0]), .IN2(ce), .Q(n7132) );
  MUX21X1 U9421 ( .IN1(\mem1[255][15] ), .IN2(n1019), .S(n7403), .Q(n16555) );
  MUX21X1 U9422 ( .IN1(\mem1[255][14] ), .IN2(n997), .S(n7403), .Q(n16554) );
  MUX21X1 U9423 ( .IN1(\mem1[255][13] ), .IN2(n975), .S(n7403), .Q(n16553) );
  MUX21X1 U9424 ( .IN1(\mem1[255][12] ), .IN2(n953), .S(n7403), .Q(n16552) );
  MUX21X1 U9425 ( .IN1(\mem1[255][11] ), .IN2(n931), .S(n7403), .Q(n16551) );
  MUX21X1 U9426 ( .IN1(\mem1[255][10] ), .IN2(n909), .S(n7403), .Q(n16550) );
  MUX21X1 U9427 ( .IN1(\mem1[255][9] ), .IN2(n887), .S(n7403), .Q(n16549) );
  MUX21X1 U9428 ( .IN1(\mem1[255][8] ), .IN2(n865), .S(n7403), .Q(n16548) );
  AND2X1 U9429 ( .IN1(n7404), .IN2(n7099), .Q(n7403) );
  MUX21X1 U9430 ( .IN1(\mem1[254][15] ), .IN2(n1019), .S(n7405), .Q(n16547) );
  MUX21X1 U9431 ( .IN1(\mem1[254][14] ), .IN2(n997), .S(n7405), .Q(n16546) );
  MUX21X1 U9432 ( .IN1(\mem1[254][13] ), .IN2(n975), .S(n7405), .Q(n16545) );
  MUX21X1 U9433 ( .IN1(\mem1[254][12] ), .IN2(n953), .S(n7405), .Q(n16544) );
  MUX21X1 U9434 ( .IN1(\mem1[254][11] ), .IN2(n931), .S(n7405), .Q(n16543) );
  MUX21X1 U9435 ( .IN1(\mem1[254][10] ), .IN2(n909), .S(n7405), .Q(n16542) );
  MUX21X1 U9436 ( .IN1(\mem1[254][9] ), .IN2(n887), .S(n7405), .Q(n16541) );
  MUX21X1 U9437 ( .IN1(\mem1[254][8] ), .IN2(n865), .S(n7405), .Q(n16540) );
  AND2X1 U9438 ( .IN1(n7404), .IN2(n7102), .Q(n7405) );
  MUX21X1 U9439 ( .IN1(\mem1[253][15] ), .IN2(n1019), .S(n7406), .Q(n16539) );
  MUX21X1 U9440 ( .IN1(\mem1[253][14] ), .IN2(n997), .S(n7406), .Q(n16538) );
  MUX21X1 U9441 ( .IN1(\mem1[253][13] ), .IN2(n975), .S(n7406), .Q(n16537) );
  MUX21X1 U9442 ( .IN1(\mem1[253][12] ), .IN2(n953), .S(n7406), .Q(n16536) );
  MUX21X1 U9443 ( .IN1(\mem1[253][11] ), .IN2(n931), .S(n7406), .Q(n16535) );
  MUX21X1 U9444 ( .IN1(\mem1[253][10] ), .IN2(n909), .S(n7406), .Q(n16534) );
  MUX21X1 U9445 ( .IN1(\mem1[253][9] ), .IN2(n887), .S(n7406), .Q(n16533) );
  MUX21X1 U9446 ( .IN1(\mem1[253][8] ), .IN2(n865), .S(n7406), .Q(n16532) );
  AND2X1 U9447 ( .IN1(n7404), .IN2(n7104), .Q(n7406) );
  MUX21X1 U9448 ( .IN1(\mem1[252][15] ), .IN2(n1019), .S(n7407), .Q(n16531) );
  MUX21X1 U9449 ( .IN1(\mem1[252][14] ), .IN2(n997), .S(n7407), .Q(n16530) );
  MUX21X1 U9450 ( .IN1(\mem1[252][13] ), .IN2(n975), .S(n7407), .Q(n16529) );
  MUX21X1 U9451 ( .IN1(\mem1[252][12] ), .IN2(n953), .S(n7407), .Q(n16528) );
  MUX21X1 U9452 ( .IN1(\mem1[252][11] ), .IN2(n931), .S(n7407), .Q(n16527) );
  MUX21X1 U9453 ( .IN1(\mem1[252][10] ), .IN2(n909), .S(n7407), .Q(n16526) );
  MUX21X1 U9454 ( .IN1(\mem1[252][9] ), .IN2(n887), .S(n7407), .Q(n16525) );
  MUX21X1 U9455 ( .IN1(\mem1[252][8] ), .IN2(n865), .S(n7407), .Q(n16524) );
  AND2X1 U9456 ( .IN1(n7404), .IN2(n7106), .Q(n7407) );
  MUX21X1 U9457 ( .IN1(\mem1[251][15] ), .IN2(n1019), .S(n7408), .Q(n16523) );
  MUX21X1 U9458 ( .IN1(\mem1[251][14] ), .IN2(n997), .S(n7408), .Q(n16522) );
  MUX21X1 U9459 ( .IN1(\mem1[251][13] ), .IN2(n975), .S(n7408), .Q(n16521) );
  MUX21X1 U9460 ( .IN1(\mem1[251][12] ), .IN2(n953), .S(n7408), .Q(n16520) );
  MUX21X1 U9461 ( .IN1(\mem1[251][11] ), .IN2(n931), .S(n7408), .Q(n16519) );
  MUX21X1 U9462 ( .IN1(\mem1[251][10] ), .IN2(n909), .S(n7408), .Q(n16518) );
  MUX21X1 U9463 ( .IN1(\mem1[251][9] ), .IN2(n887), .S(n7408), .Q(n16517) );
  MUX21X1 U9464 ( .IN1(\mem1[251][8] ), .IN2(n865), .S(n7408), .Q(n16516) );
  AND2X1 U9465 ( .IN1(n7404), .IN2(n7108), .Q(n7408) );
  MUX21X1 U9466 ( .IN1(\mem1[250][15] ), .IN2(n1019), .S(n7409), .Q(n16515) );
  MUX21X1 U9467 ( .IN1(\mem1[250][14] ), .IN2(n997), .S(n7409), .Q(n16514) );
  MUX21X1 U9468 ( .IN1(\mem1[250][13] ), .IN2(n975), .S(n7409), .Q(n16513) );
  MUX21X1 U9469 ( .IN1(\mem1[250][12] ), .IN2(n953), .S(n7409), .Q(n16512) );
  MUX21X1 U9470 ( .IN1(\mem1[250][11] ), .IN2(n931), .S(n7409), .Q(n16511) );
  MUX21X1 U9471 ( .IN1(\mem1[250][10] ), .IN2(n909), .S(n7409), .Q(n16510) );
  MUX21X1 U9472 ( .IN1(\mem1[250][9] ), .IN2(n887), .S(n7409), .Q(n16509) );
  MUX21X1 U9473 ( .IN1(\mem1[250][8] ), .IN2(n865), .S(n7409), .Q(n16508) );
  AND2X1 U9474 ( .IN1(n7404), .IN2(n7110), .Q(n7409) );
  MUX21X1 U9475 ( .IN1(\mem1[249][15] ), .IN2(n1019), .S(n7410), .Q(n16507) );
  MUX21X1 U9476 ( .IN1(\mem1[249][14] ), .IN2(n997), .S(n7410), .Q(n16506) );
  MUX21X1 U9477 ( .IN1(\mem1[249][13] ), .IN2(n975), .S(n7410), .Q(n16505) );
  MUX21X1 U9478 ( .IN1(\mem1[249][12] ), .IN2(n953), .S(n7410), .Q(n16504) );
  MUX21X1 U9479 ( .IN1(\mem1[249][11] ), .IN2(n931), .S(n7410), .Q(n16503) );
  MUX21X1 U9480 ( .IN1(\mem1[249][10] ), .IN2(n909), .S(n7410), .Q(n16502) );
  MUX21X1 U9481 ( .IN1(\mem1[249][9] ), .IN2(n887), .S(n7410), .Q(n16501) );
  MUX21X1 U9482 ( .IN1(\mem1[249][8] ), .IN2(n865), .S(n7410), .Q(n16500) );
  AND2X1 U9483 ( .IN1(n7404), .IN2(n7112), .Q(n7410) );
  MUX21X1 U9484 ( .IN1(\mem1[248][15] ), .IN2(n1019), .S(n7411), .Q(n16499) );
  MUX21X1 U9485 ( .IN1(\mem1[248][14] ), .IN2(n997), .S(n7411), .Q(n16498) );
  MUX21X1 U9486 ( .IN1(\mem1[248][13] ), .IN2(n975), .S(n7411), .Q(n16497) );
  MUX21X1 U9487 ( .IN1(\mem1[248][12] ), .IN2(n953), .S(n7411), .Q(n16496) );
  MUX21X1 U9488 ( .IN1(\mem1[248][11] ), .IN2(n931), .S(n7411), .Q(n16495) );
  MUX21X1 U9489 ( .IN1(\mem1[248][10] ), .IN2(n909), .S(n7411), .Q(n16494) );
  MUX21X1 U9490 ( .IN1(\mem1[248][9] ), .IN2(n887), .S(n7411), .Q(n16493) );
  MUX21X1 U9491 ( .IN1(\mem1[248][8] ), .IN2(n865), .S(n7411), .Q(n16492) );
  AND2X1 U9492 ( .IN1(n7404), .IN2(n7114), .Q(n7411) );
  MUX21X1 U9493 ( .IN1(\mem1[247][15] ), .IN2(n1019), .S(n7412), .Q(n16491) );
  MUX21X1 U9494 ( .IN1(\mem1[247][14] ), .IN2(n997), .S(n7412), .Q(n16490) );
  MUX21X1 U9495 ( .IN1(\mem1[247][13] ), .IN2(n975), .S(n7412), .Q(n16489) );
  MUX21X1 U9496 ( .IN1(\mem1[247][12] ), .IN2(n953), .S(n7412), .Q(n16488) );
  MUX21X1 U9497 ( .IN1(\mem1[247][11] ), .IN2(n931), .S(n7412), .Q(n16487) );
  MUX21X1 U9498 ( .IN1(\mem1[247][10] ), .IN2(n909), .S(n7412), .Q(n16486) );
  MUX21X1 U9499 ( .IN1(\mem1[247][9] ), .IN2(n887), .S(n7412), .Q(n16485) );
  MUX21X1 U9500 ( .IN1(\mem1[247][8] ), .IN2(n865), .S(n7412), .Q(n16484) );
  AND2X1 U9501 ( .IN1(n7404), .IN2(n7116), .Q(n7412) );
  MUX21X1 U9502 ( .IN1(\mem1[246][15] ), .IN2(n1019), .S(n7413), .Q(n16483) );
  MUX21X1 U9503 ( .IN1(\mem1[246][14] ), .IN2(n997), .S(n7413), .Q(n16482) );
  MUX21X1 U9504 ( .IN1(\mem1[246][13] ), .IN2(n975), .S(n7413), .Q(n16481) );
  MUX21X1 U9505 ( .IN1(\mem1[246][12] ), .IN2(n953), .S(n7413), .Q(n16480) );
  MUX21X1 U9506 ( .IN1(\mem1[246][11] ), .IN2(n931), .S(n7413), .Q(n16479) );
  MUX21X1 U9507 ( .IN1(\mem1[246][10] ), .IN2(n909), .S(n7413), .Q(n16478) );
  MUX21X1 U9508 ( .IN1(\mem1[246][9] ), .IN2(n887), .S(n7413), .Q(n16477) );
  MUX21X1 U9509 ( .IN1(\mem1[246][8] ), .IN2(n865), .S(n7413), .Q(n16476) );
  AND2X1 U9510 ( .IN1(n7404), .IN2(n7118), .Q(n7413) );
  MUX21X1 U9511 ( .IN1(\mem1[245][15] ), .IN2(n1019), .S(n7414), .Q(n16475) );
  MUX21X1 U9512 ( .IN1(\mem1[245][14] ), .IN2(n997), .S(n7414), .Q(n16474) );
  MUX21X1 U9513 ( .IN1(\mem1[245][13] ), .IN2(n975), .S(n7414), .Q(n16473) );
  MUX21X1 U9514 ( .IN1(\mem1[245][12] ), .IN2(n953), .S(n7414), .Q(n16472) );
  MUX21X1 U9515 ( .IN1(\mem1[245][11] ), .IN2(n931), .S(n7414), .Q(n16471) );
  MUX21X1 U9516 ( .IN1(\mem1[245][10] ), .IN2(n909), .S(n7414), .Q(n16470) );
  MUX21X1 U9517 ( .IN1(\mem1[245][9] ), .IN2(n887), .S(n7414), .Q(n16469) );
  MUX21X1 U9518 ( .IN1(\mem1[245][8] ), .IN2(n865), .S(n7414), .Q(n16468) );
  AND2X1 U9519 ( .IN1(n7404), .IN2(n7120), .Q(n7414) );
  MUX21X1 U9520 ( .IN1(\mem1[244][15] ), .IN2(n1019), .S(n7415), .Q(n16467) );
  MUX21X1 U9521 ( .IN1(\mem1[244][14] ), .IN2(n997), .S(n7415), .Q(n16466) );
  MUX21X1 U9522 ( .IN1(\mem1[244][13] ), .IN2(n975), .S(n7415), .Q(n16465) );
  MUX21X1 U9523 ( .IN1(\mem1[244][12] ), .IN2(n953), .S(n7415), .Q(n16464) );
  MUX21X1 U9524 ( .IN1(\mem1[244][11] ), .IN2(n931), .S(n7415), .Q(n16463) );
  MUX21X1 U9525 ( .IN1(\mem1[244][10] ), .IN2(n909), .S(n7415), .Q(n16462) );
  MUX21X1 U9526 ( .IN1(\mem1[244][9] ), .IN2(n887), .S(n7415), .Q(n16461) );
  MUX21X1 U9527 ( .IN1(\mem1[244][8] ), .IN2(n865), .S(n7415), .Q(n16460) );
  AND2X1 U9528 ( .IN1(n7404), .IN2(n7122), .Q(n7415) );
  MUX21X1 U9529 ( .IN1(\mem1[243][15] ), .IN2(n1020), .S(n7416), .Q(n16459) );
  MUX21X1 U9530 ( .IN1(\mem1[243][14] ), .IN2(n998), .S(n7416), .Q(n16458) );
  MUX21X1 U9531 ( .IN1(\mem1[243][13] ), .IN2(n976), .S(n7416), .Q(n16457) );
  MUX21X1 U9532 ( .IN1(\mem1[243][12] ), .IN2(n954), .S(n7416), .Q(n16456) );
  MUX21X1 U9533 ( .IN1(\mem1[243][11] ), .IN2(n932), .S(n7416), .Q(n16455) );
  MUX21X1 U9534 ( .IN1(\mem1[243][10] ), .IN2(n910), .S(n7416), .Q(n16454) );
  MUX21X1 U9535 ( .IN1(\mem1[243][9] ), .IN2(n888), .S(n7416), .Q(n16453) );
  MUX21X1 U9536 ( .IN1(\mem1[243][8] ), .IN2(n866), .S(n7416), .Q(n16452) );
  AND2X1 U9537 ( .IN1(n7404), .IN2(n7124), .Q(n7416) );
  MUX21X1 U9538 ( .IN1(\mem1[242][15] ), .IN2(n1020), .S(n7417), .Q(n16451) );
  MUX21X1 U9539 ( .IN1(\mem1[242][14] ), .IN2(n998), .S(n7417), .Q(n16450) );
  MUX21X1 U9540 ( .IN1(\mem1[242][13] ), .IN2(n976), .S(n7417), .Q(n16449) );
  MUX21X1 U9541 ( .IN1(\mem1[242][12] ), .IN2(n954), .S(n7417), .Q(n16448) );
  MUX21X1 U9542 ( .IN1(\mem1[242][11] ), .IN2(n932), .S(n7417), .Q(n16447) );
  MUX21X1 U9543 ( .IN1(\mem1[242][10] ), .IN2(n910), .S(n7417), .Q(n16446) );
  MUX21X1 U9544 ( .IN1(\mem1[242][9] ), .IN2(n888), .S(n7417), .Q(n16445) );
  MUX21X1 U9545 ( .IN1(\mem1[242][8] ), .IN2(n866), .S(n7417), .Q(n16444) );
  AND2X1 U9546 ( .IN1(n7404), .IN2(n7126), .Q(n7417) );
  MUX21X1 U9547 ( .IN1(\mem1[241][15] ), .IN2(n1020), .S(n7418), .Q(n16443) );
  MUX21X1 U9548 ( .IN1(\mem1[241][14] ), .IN2(n998), .S(n7418), .Q(n16442) );
  MUX21X1 U9549 ( .IN1(\mem1[241][13] ), .IN2(n976), .S(n7418), .Q(n16441) );
  MUX21X1 U9550 ( .IN1(\mem1[241][12] ), .IN2(n954), .S(n7418), .Q(n16440) );
  MUX21X1 U9551 ( .IN1(\mem1[241][11] ), .IN2(n932), .S(n7418), .Q(n16439) );
  MUX21X1 U9552 ( .IN1(\mem1[241][10] ), .IN2(n910), .S(n7418), .Q(n16438) );
  MUX21X1 U9553 ( .IN1(\mem1[241][9] ), .IN2(n888), .S(n7418), .Q(n16437) );
  MUX21X1 U9554 ( .IN1(\mem1[241][8] ), .IN2(n866), .S(n7418), .Q(n16436) );
  AND2X1 U9555 ( .IN1(n7404), .IN2(n7128), .Q(n7418) );
  MUX21X1 U9556 ( .IN1(\mem1[240][15] ), .IN2(n1020), .S(n7419), .Q(n16435) );
  MUX21X1 U9557 ( .IN1(\mem1[240][14] ), .IN2(n998), .S(n7419), .Q(n16434) );
  MUX21X1 U9558 ( .IN1(\mem1[240][13] ), .IN2(n976), .S(n7419), .Q(n16433) );
  MUX21X1 U9559 ( .IN1(\mem1[240][12] ), .IN2(n954), .S(n7419), .Q(n16432) );
  MUX21X1 U9560 ( .IN1(\mem1[240][11] ), .IN2(n932), .S(n7419), .Q(n16431) );
  MUX21X1 U9561 ( .IN1(\mem1[240][10] ), .IN2(n910), .S(n7419), .Q(n16430) );
  MUX21X1 U9562 ( .IN1(\mem1[240][9] ), .IN2(n888), .S(n7419), .Q(n16429) );
  MUX21X1 U9563 ( .IN1(\mem1[240][8] ), .IN2(n866), .S(n7419), .Q(n16428) );
  AND2X1 U9564 ( .IN1(n7404), .IN2(n7130), .Q(n7419) );
  AND2X1 U9565 ( .IN1(n7420), .IN2(n7131), .Q(n7404) );
  MUX21X1 U9566 ( .IN1(\mem1[239][15] ), .IN2(n1020), .S(n7421), .Q(n16427) );
  MUX21X1 U9567 ( .IN1(\mem1[239][14] ), .IN2(n998), .S(n7421), .Q(n16426) );
  MUX21X1 U9568 ( .IN1(\mem1[239][13] ), .IN2(n976), .S(n7421), .Q(n16425) );
  MUX21X1 U9569 ( .IN1(\mem1[239][12] ), .IN2(n954), .S(n7421), .Q(n16424) );
  MUX21X1 U9570 ( .IN1(\mem1[239][11] ), .IN2(n932), .S(n7421), .Q(n16423) );
  MUX21X1 U9571 ( .IN1(\mem1[239][10] ), .IN2(n910), .S(n7421), .Q(n16422) );
  MUX21X1 U9572 ( .IN1(\mem1[239][9] ), .IN2(n888), .S(n7421), .Q(n16421) );
  MUX21X1 U9573 ( .IN1(\mem1[239][8] ), .IN2(n866), .S(n7421), .Q(n16420) );
  AND2X1 U9574 ( .IN1(n7422), .IN2(n7099), .Q(n7421) );
  MUX21X1 U9575 ( .IN1(\mem1[238][15] ), .IN2(n1020), .S(n7423), .Q(n16419) );
  MUX21X1 U9576 ( .IN1(\mem1[238][14] ), .IN2(n998), .S(n7423), .Q(n16418) );
  MUX21X1 U9577 ( .IN1(\mem1[238][13] ), .IN2(n976), .S(n7423), .Q(n16417) );
  MUX21X1 U9578 ( .IN1(\mem1[238][12] ), .IN2(n954), .S(n7423), .Q(n16416) );
  MUX21X1 U9579 ( .IN1(\mem1[238][11] ), .IN2(n932), .S(n7423), .Q(n16415) );
  MUX21X1 U9580 ( .IN1(\mem1[238][10] ), .IN2(n910), .S(n7423), .Q(n16414) );
  MUX21X1 U9581 ( .IN1(\mem1[238][9] ), .IN2(n888), .S(n7423), .Q(n16413) );
  MUX21X1 U9582 ( .IN1(\mem1[238][8] ), .IN2(n866), .S(n7423), .Q(n16412) );
  AND2X1 U9583 ( .IN1(n7422), .IN2(n7102), .Q(n7423) );
  MUX21X1 U9584 ( .IN1(\mem1[237][15] ), .IN2(n1020), .S(n7424), .Q(n16411) );
  MUX21X1 U9585 ( .IN1(\mem1[237][14] ), .IN2(n998), .S(n7424), .Q(n16410) );
  MUX21X1 U9586 ( .IN1(\mem1[237][13] ), .IN2(n976), .S(n7424), .Q(n16409) );
  MUX21X1 U9587 ( .IN1(\mem1[237][12] ), .IN2(n954), .S(n7424), .Q(n16408) );
  MUX21X1 U9588 ( .IN1(\mem1[237][11] ), .IN2(n932), .S(n7424), .Q(n16407) );
  MUX21X1 U9589 ( .IN1(\mem1[237][10] ), .IN2(n910), .S(n7424), .Q(n16406) );
  MUX21X1 U9590 ( .IN1(\mem1[237][9] ), .IN2(n888), .S(n7424), .Q(n16405) );
  MUX21X1 U9591 ( .IN1(\mem1[237][8] ), .IN2(n866), .S(n7424), .Q(n16404) );
  AND2X1 U9592 ( .IN1(n7422), .IN2(n7104), .Q(n7424) );
  MUX21X1 U9593 ( .IN1(\mem1[236][15] ), .IN2(n1020), .S(n7425), .Q(n16403) );
  MUX21X1 U9594 ( .IN1(\mem1[236][14] ), .IN2(n998), .S(n7425), .Q(n16402) );
  MUX21X1 U9595 ( .IN1(\mem1[236][13] ), .IN2(n976), .S(n7425), .Q(n16401) );
  MUX21X1 U9596 ( .IN1(\mem1[236][12] ), .IN2(n954), .S(n7425), .Q(n16400) );
  MUX21X1 U9597 ( .IN1(\mem1[236][11] ), .IN2(n932), .S(n7425), .Q(n16399) );
  MUX21X1 U9598 ( .IN1(\mem1[236][10] ), .IN2(n910), .S(n7425), .Q(n16398) );
  MUX21X1 U9599 ( .IN1(\mem1[236][9] ), .IN2(n888), .S(n7425), .Q(n16397) );
  MUX21X1 U9600 ( .IN1(\mem1[236][8] ), .IN2(n866), .S(n7425), .Q(n16396) );
  AND2X1 U9601 ( .IN1(n7422), .IN2(n7106), .Q(n7425) );
  MUX21X1 U9602 ( .IN1(\mem1[235][15] ), .IN2(n1020), .S(n7426), .Q(n16395) );
  MUX21X1 U9603 ( .IN1(\mem1[235][14] ), .IN2(n998), .S(n7426), .Q(n16394) );
  MUX21X1 U9604 ( .IN1(\mem1[235][13] ), .IN2(n976), .S(n7426), .Q(n16393) );
  MUX21X1 U9605 ( .IN1(\mem1[235][12] ), .IN2(n954), .S(n7426), .Q(n16392) );
  MUX21X1 U9606 ( .IN1(\mem1[235][11] ), .IN2(n932), .S(n7426), .Q(n16391) );
  MUX21X1 U9607 ( .IN1(\mem1[235][10] ), .IN2(n910), .S(n7426), .Q(n16390) );
  MUX21X1 U9608 ( .IN1(\mem1[235][9] ), .IN2(n888), .S(n7426), .Q(n16389) );
  MUX21X1 U9609 ( .IN1(\mem1[235][8] ), .IN2(n866), .S(n7426), .Q(n16388) );
  AND2X1 U9610 ( .IN1(n7422), .IN2(n7108), .Q(n7426) );
  MUX21X1 U9611 ( .IN1(\mem1[234][15] ), .IN2(n1020), .S(n7427), .Q(n16387) );
  MUX21X1 U9612 ( .IN1(\mem1[234][14] ), .IN2(n998), .S(n7427), .Q(n16386) );
  MUX21X1 U9613 ( .IN1(\mem1[234][13] ), .IN2(n976), .S(n7427), .Q(n16385) );
  MUX21X1 U9614 ( .IN1(\mem1[234][12] ), .IN2(n954), .S(n7427), .Q(n16384) );
  MUX21X1 U9615 ( .IN1(\mem1[234][11] ), .IN2(n932), .S(n7427), .Q(n16383) );
  MUX21X1 U9616 ( .IN1(\mem1[234][10] ), .IN2(n910), .S(n7427), .Q(n16382) );
  MUX21X1 U9617 ( .IN1(\mem1[234][9] ), .IN2(n888), .S(n7427), .Q(n16381) );
  MUX21X1 U9618 ( .IN1(\mem1[234][8] ), .IN2(n866), .S(n7427), .Q(n16380) );
  AND2X1 U9619 ( .IN1(n7422), .IN2(n7110), .Q(n7427) );
  MUX21X1 U9620 ( .IN1(\mem1[233][15] ), .IN2(n1020), .S(n7428), .Q(n16379) );
  MUX21X1 U9621 ( .IN1(\mem1[233][14] ), .IN2(n998), .S(n7428), .Q(n16378) );
  MUX21X1 U9622 ( .IN1(\mem1[233][13] ), .IN2(n976), .S(n7428), .Q(n16377) );
  MUX21X1 U9623 ( .IN1(\mem1[233][12] ), .IN2(n954), .S(n7428), .Q(n16376) );
  MUX21X1 U9624 ( .IN1(\mem1[233][11] ), .IN2(n932), .S(n7428), .Q(n16375) );
  MUX21X1 U9625 ( .IN1(\mem1[233][10] ), .IN2(n910), .S(n7428), .Q(n16374) );
  MUX21X1 U9626 ( .IN1(\mem1[233][9] ), .IN2(n888), .S(n7428), .Q(n16373) );
  MUX21X1 U9627 ( .IN1(\mem1[233][8] ), .IN2(n866), .S(n7428), .Q(n16372) );
  AND2X1 U9628 ( .IN1(n7422), .IN2(n7112), .Q(n7428) );
  MUX21X1 U9629 ( .IN1(\mem1[232][15] ), .IN2(n1020), .S(n7429), .Q(n16371) );
  MUX21X1 U9630 ( .IN1(\mem1[232][14] ), .IN2(n998), .S(n7429), .Q(n16370) );
  MUX21X1 U9631 ( .IN1(\mem1[232][13] ), .IN2(n976), .S(n7429), .Q(n16369) );
  MUX21X1 U9632 ( .IN1(\mem1[232][12] ), .IN2(n954), .S(n7429), .Q(n16368) );
  MUX21X1 U9633 ( .IN1(\mem1[232][11] ), .IN2(n932), .S(n7429), .Q(n16367) );
  MUX21X1 U9634 ( .IN1(\mem1[232][10] ), .IN2(n910), .S(n7429), .Q(n16366) );
  MUX21X1 U9635 ( .IN1(\mem1[232][9] ), .IN2(n888), .S(n7429), .Q(n16365) );
  MUX21X1 U9636 ( .IN1(\mem1[232][8] ), .IN2(n866), .S(n7429), .Q(n16364) );
  AND2X1 U9637 ( .IN1(n7422), .IN2(n7114), .Q(n7429) );
  MUX21X1 U9638 ( .IN1(\mem1[231][15] ), .IN2(n1021), .S(n7430), .Q(n16363) );
  MUX21X1 U9639 ( .IN1(\mem1[231][14] ), .IN2(n999), .S(n7430), .Q(n16362) );
  MUX21X1 U9640 ( .IN1(\mem1[231][13] ), .IN2(n977), .S(n7430), .Q(n16361) );
  MUX21X1 U9641 ( .IN1(\mem1[231][12] ), .IN2(n955), .S(n7430), .Q(n16360) );
  MUX21X1 U9642 ( .IN1(\mem1[231][11] ), .IN2(n933), .S(n7430), .Q(n16359) );
  MUX21X1 U9643 ( .IN1(\mem1[231][10] ), .IN2(n911), .S(n7430), .Q(n16358) );
  MUX21X1 U9644 ( .IN1(\mem1[231][9] ), .IN2(n889), .S(n7430), .Q(n16357) );
  MUX21X1 U9645 ( .IN1(\mem1[231][8] ), .IN2(n867), .S(n7430), .Q(n16356) );
  AND2X1 U9646 ( .IN1(n7422), .IN2(n7116), .Q(n7430) );
  MUX21X1 U9647 ( .IN1(\mem1[230][15] ), .IN2(n1021), .S(n7431), .Q(n16355) );
  MUX21X1 U9648 ( .IN1(\mem1[230][14] ), .IN2(n999), .S(n7431), .Q(n16354) );
  MUX21X1 U9649 ( .IN1(\mem1[230][13] ), .IN2(n977), .S(n7431), .Q(n16353) );
  MUX21X1 U9650 ( .IN1(\mem1[230][12] ), .IN2(n955), .S(n7431), .Q(n16352) );
  MUX21X1 U9651 ( .IN1(\mem1[230][11] ), .IN2(n933), .S(n7431), .Q(n16351) );
  MUX21X1 U9652 ( .IN1(\mem1[230][10] ), .IN2(n911), .S(n7431), .Q(n16350) );
  MUX21X1 U9653 ( .IN1(\mem1[230][9] ), .IN2(n889), .S(n7431), .Q(n16349) );
  MUX21X1 U9654 ( .IN1(\mem1[230][8] ), .IN2(n867), .S(n7431), .Q(n16348) );
  AND2X1 U9655 ( .IN1(n7422), .IN2(n7118), .Q(n7431) );
  MUX21X1 U9656 ( .IN1(\mem1[229][15] ), .IN2(n1021), .S(n7432), .Q(n16347) );
  MUX21X1 U9657 ( .IN1(\mem1[229][14] ), .IN2(n999), .S(n7432), .Q(n16346) );
  MUX21X1 U9658 ( .IN1(\mem1[229][13] ), .IN2(n977), .S(n7432), .Q(n16345) );
  MUX21X1 U9659 ( .IN1(\mem1[229][12] ), .IN2(n955), .S(n7432), .Q(n16344) );
  MUX21X1 U9660 ( .IN1(\mem1[229][11] ), .IN2(n933), .S(n7432), .Q(n16343) );
  MUX21X1 U9661 ( .IN1(\mem1[229][10] ), .IN2(n911), .S(n7432), .Q(n16342) );
  MUX21X1 U9662 ( .IN1(\mem1[229][9] ), .IN2(n889), .S(n7432), .Q(n16341) );
  MUX21X1 U9663 ( .IN1(\mem1[229][8] ), .IN2(n867), .S(n7432), .Q(n16340) );
  AND2X1 U9664 ( .IN1(n7422), .IN2(n7120), .Q(n7432) );
  MUX21X1 U9665 ( .IN1(\mem1[228][15] ), .IN2(n1021), .S(n7433), .Q(n16339) );
  MUX21X1 U9666 ( .IN1(\mem1[228][14] ), .IN2(n999), .S(n7433), .Q(n16338) );
  MUX21X1 U9667 ( .IN1(\mem1[228][13] ), .IN2(n977), .S(n7433), .Q(n16337) );
  MUX21X1 U9668 ( .IN1(\mem1[228][12] ), .IN2(n955), .S(n7433), .Q(n16336) );
  MUX21X1 U9669 ( .IN1(\mem1[228][11] ), .IN2(n933), .S(n7433), .Q(n16335) );
  MUX21X1 U9670 ( .IN1(\mem1[228][10] ), .IN2(n911), .S(n7433), .Q(n16334) );
  MUX21X1 U9671 ( .IN1(\mem1[228][9] ), .IN2(n889), .S(n7433), .Q(n16333) );
  MUX21X1 U9672 ( .IN1(\mem1[228][8] ), .IN2(n867), .S(n7433), .Q(n16332) );
  AND2X1 U9673 ( .IN1(n7422), .IN2(n7122), .Q(n7433) );
  MUX21X1 U9674 ( .IN1(\mem1[227][15] ), .IN2(n1021), .S(n7434), .Q(n16331) );
  MUX21X1 U9675 ( .IN1(\mem1[227][14] ), .IN2(n999), .S(n7434), .Q(n16330) );
  MUX21X1 U9676 ( .IN1(\mem1[227][13] ), .IN2(n977), .S(n7434), .Q(n16329) );
  MUX21X1 U9677 ( .IN1(\mem1[227][12] ), .IN2(n955), .S(n7434), .Q(n16328) );
  MUX21X1 U9678 ( .IN1(\mem1[227][11] ), .IN2(n933), .S(n7434), .Q(n16327) );
  MUX21X1 U9679 ( .IN1(\mem1[227][10] ), .IN2(n911), .S(n7434), .Q(n16326) );
  MUX21X1 U9680 ( .IN1(\mem1[227][9] ), .IN2(n889), .S(n7434), .Q(n16325) );
  MUX21X1 U9681 ( .IN1(\mem1[227][8] ), .IN2(n867), .S(n7434), .Q(n16324) );
  AND2X1 U9682 ( .IN1(n7422), .IN2(n7124), .Q(n7434) );
  MUX21X1 U9683 ( .IN1(\mem1[226][15] ), .IN2(n1021), .S(n7435), .Q(n16323) );
  MUX21X1 U9684 ( .IN1(\mem1[226][14] ), .IN2(n999), .S(n7435), .Q(n16322) );
  MUX21X1 U9685 ( .IN1(\mem1[226][13] ), .IN2(n977), .S(n7435), .Q(n16321) );
  MUX21X1 U9686 ( .IN1(\mem1[226][12] ), .IN2(n955), .S(n7435), .Q(n16320) );
  MUX21X1 U9687 ( .IN1(\mem1[226][11] ), .IN2(n933), .S(n7435), .Q(n16319) );
  MUX21X1 U9688 ( .IN1(\mem1[226][10] ), .IN2(n911), .S(n7435), .Q(n16318) );
  MUX21X1 U9689 ( .IN1(\mem1[226][9] ), .IN2(n889), .S(n7435), .Q(n16317) );
  MUX21X1 U9690 ( .IN1(\mem1[226][8] ), .IN2(n867), .S(n7435), .Q(n16316) );
  AND2X1 U9691 ( .IN1(n7422), .IN2(n7126), .Q(n7435) );
  MUX21X1 U9692 ( .IN1(\mem1[225][15] ), .IN2(n1021), .S(n7436), .Q(n16315) );
  MUX21X1 U9693 ( .IN1(\mem1[225][14] ), .IN2(n999), .S(n7436), .Q(n16314) );
  MUX21X1 U9694 ( .IN1(\mem1[225][13] ), .IN2(n977), .S(n7436), .Q(n16313) );
  MUX21X1 U9695 ( .IN1(\mem1[225][12] ), .IN2(n955), .S(n7436), .Q(n16312) );
  MUX21X1 U9696 ( .IN1(\mem1[225][11] ), .IN2(n933), .S(n7436), .Q(n16311) );
  MUX21X1 U9697 ( .IN1(\mem1[225][10] ), .IN2(n911), .S(n7436), .Q(n16310) );
  MUX21X1 U9698 ( .IN1(\mem1[225][9] ), .IN2(n889), .S(n7436), .Q(n16309) );
  MUX21X1 U9699 ( .IN1(\mem1[225][8] ), .IN2(n867), .S(n7436), .Q(n16308) );
  AND2X1 U9700 ( .IN1(n7422), .IN2(n7128), .Q(n7436) );
  MUX21X1 U9701 ( .IN1(\mem1[224][15] ), .IN2(n1021), .S(n7437), .Q(n16307) );
  MUX21X1 U9702 ( .IN1(\mem1[224][14] ), .IN2(n999), .S(n7437), .Q(n16306) );
  MUX21X1 U9703 ( .IN1(\mem1[224][13] ), .IN2(n977), .S(n7437), .Q(n16305) );
  MUX21X1 U9704 ( .IN1(\mem1[224][12] ), .IN2(n955), .S(n7437), .Q(n16304) );
  MUX21X1 U9705 ( .IN1(\mem1[224][11] ), .IN2(n933), .S(n7437), .Q(n16303) );
  MUX21X1 U9706 ( .IN1(\mem1[224][10] ), .IN2(n911), .S(n7437), .Q(n16302) );
  MUX21X1 U9707 ( .IN1(\mem1[224][9] ), .IN2(n889), .S(n7437), .Q(n16301) );
  MUX21X1 U9708 ( .IN1(\mem1[224][8] ), .IN2(n867), .S(n7437), .Q(n16300) );
  AND2X1 U9709 ( .IN1(n7422), .IN2(n7130), .Q(n7437) );
  AND2X1 U9710 ( .IN1(n7420), .IN2(n7150), .Q(n7422) );
  MUX21X1 U9711 ( .IN1(\mem1[223][15] ), .IN2(n1021), .S(n7438), .Q(n16299) );
  MUX21X1 U9712 ( .IN1(\mem1[223][14] ), .IN2(n999), .S(n7438), .Q(n16298) );
  MUX21X1 U9713 ( .IN1(\mem1[223][13] ), .IN2(n977), .S(n7438), .Q(n16297) );
  MUX21X1 U9714 ( .IN1(\mem1[223][12] ), .IN2(n955), .S(n7438), .Q(n16296) );
  MUX21X1 U9715 ( .IN1(\mem1[223][11] ), .IN2(n933), .S(n7438), .Q(n16295) );
  MUX21X1 U9716 ( .IN1(\mem1[223][10] ), .IN2(n911), .S(n7438), .Q(n16294) );
  MUX21X1 U9717 ( .IN1(\mem1[223][9] ), .IN2(n889), .S(n7438), .Q(n16293) );
  MUX21X1 U9718 ( .IN1(\mem1[223][8] ), .IN2(n867), .S(n7438), .Q(n16292) );
  AND2X1 U9719 ( .IN1(n7439), .IN2(n7099), .Q(n7438) );
  MUX21X1 U9720 ( .IN1(\mem1[222][15] ), .IN2(n1021), .S(n7440), .Q(n16291) );
  MUX21X1 U9721 ( .IN1(\mem1[222][14] ), .IN2(n999), .S(n7440), .Q(n16290) );
  MUX21X1 U9722 ( .IN1(\mem1[222][13] ), .IN2(n977), .S(n7440), .Q(n16289) );
  MUX21X1 U9723 ( .IN1(\mem1[222][12] ), .IN2(n955), .S(n7440), .Q(n16288) );
  MUX21X1 U9724 ( .IN1(\mem1[222][11] ), .IN2(n933), .S(n7440), .Q(n16287) );
  MUX21X1 U9725 ( .IN1(\mem1[222][10] ), .IN2(n911), .S(n7440), .Q(n16286) );
  MUX21X1 U9726 ( .IN1(\mem1[222][9] ), .IN2(n889), .S(n7440), .Q(n16285) );
  MUX21X1 U9727 ( .IN1(\mem1[222][8] ), .IN2(n867), .S(n7440), .Q(n16284) );
  AND2X1 U9728 ( .IN1(n7439), .IN2(n7102), .Q(n7440) );
  MUX21X1 U9729 ( .IN1(\mem1[221][15] ), .IN2(n1021), .S(n7441), .Q(n16283) );
  MUX21X1 U9730 ( .IN1(\mem1[221][14] ), .IN2(n999), .S(n7441), .Q(n16282) );
  MUX21X1 U9731 ( .IN1(\mem1[221][13] ), .IN2(n977), .S(n7441), .Q(n16281) );
  MUX21X1 U9732 ( .IN1(\mem1[221][12] ), .IN2(n955), .S(n7441), .Q(n16280) );
  MUX21X1 U9733 ( .IN1(\mem1[221][11] ), .IN2(n933), .S(n7441), .Q(n16279) );
  MUX21X1 U9734 ( .IN1(\mem1[221][10] ), .IN2(n911), .S(n7441), .Q(n16278) );
  MUX21X1 U9735 ( .IN1(\mem1[221][9] ), .IN2(n889), .S(n7441), .Q(n16277) );
  MUX21X1 U9736 ( .IN1(\mem1[221][8] ), .IN2(n867), .S(n7441), .Q(n16276) );
  AND2X1 U9737 ( .IN1(n7439), .IN2(n7104), .Q(n7441) );
  MUX21X1 U9738 ( .IN1(\mem1[220][15] ), .IN2(n1021), .S(n7442), .Q(n16275) );
  MUX21X1 U9739 ( .IN1(\mem1[220][14] ), .IN2(n999), .S(n7442), .Q(n16274) );
  MUX21X1 U9740 ( .IN1(\mem1[220][13] ), .IN2(n977), .S(n7442), .Q(n16273) );
  MUX21X1 U9741 ( .IN1(\mem1[220][12] ), .IN2(n955), .S(n7442), .Q(n16272) );
  MUX21X1 U9742 ( .IN1(\mem1[220][11] ), .IN2(n933), .S(n7442), .Q(n16271) );
  MUX21X1 U9743 ( .IN1(\mem1[220][10] ), .IN2(n911), .S(n7442), .Q(n16270) );
  MUX21X1 U9744 ( .IN1(\mem1[220][9] ), .IN2(n889), .S(n7442), .Q(n16269) );
  MUX21X1 U9745 ( .IN1(\mem1[220][8] ), .IN2(n867), .S(n7442), .Q(n16268) );
  AND2X1 U9746 ( .IN1(n7439), .IN2(n7106), .Q(n7442) );
  MUX21X1 U9747 ( .IN1(\mem1[219][15] ), .IN2(n1022), .S(n7443), .Q(n16267) );
  MUX21X1 U9748 ( .IN1(\mem1[219][14] ), .IN2(n1000), .S(n7443), .Q(n16266) );
  MUX21X1 U9749 ( .IN1(\mem1[219][13] ), .IN2(n978), .S(n7443), .Q(n16265) );
  MUX21X1 U9750 ( .IN1(\mem1[219][12] ), .IN2(n956), .S(n7443), .Q(n16264) );
  MUX21X1 U9751 ( .IN1(\mem1[219][11] ), .IN2(n934), .S(n7443), .Q(n16263) );
  MUX21X1 U9752 ( .IN1(\mem1[219][10] ), .IN2(n912), .S(n7443), .Q(n16262) );
  MUX21X1 U9753 ( .IN1(\mem1[219][9] ), .IN2(n890), .S(n7443), .Q(n16261) );
  MUX21X1 U9754 ( .IN1(\mem1[219][8] ), .IN2(n868), .S(n7443), .Q(n16260) );
  AND2X1 U9755 ( .IN1(n7439), .IN2(n7108), .Q(n7443) );
  MUX21X1 U9756 ( .IN1(\mem1[218][15] ), .IN2(n1022), .S(n7444), .Q(n16259) );
  MUX21X1 U9757 ( .IN1(\mem1[218][14] ), .IN2(n1000), .S(n7444), .Q(n16258) );
  MUX21X1 U9758 ( .IN1(\mem1[218][13] ), .IN2(n978), .S(n7444), .Q(n16257) );
  MUX21X1 U9759 ( .IN1(\mem1[218][12] ), .IN2(n956), .S(n7444), .Q(n16256) );
  MUX21X1 U9760 ( .IN1(\mem1[218][11] ), .IN2(n934), .S(n7444), .Q(n16255) );
  MUX21X1 U9761 ( .IN1(\mem1[218][10] ), .IN2(n912), .S(n7444), .Q(n16254) );
  MUX21X1 U9762 ( .IN1(\mem1[218][9] ), .IN2(n890), .S(n7444), .Q(n16253) );
  MUX21X1 U9763 ( .IN1(\mem1[218][8] ), .IN2(n868), .S(n7444), .Q(n16252) );
  AND2X1 U9764 ( .IN1(n7439), .IN2(n7110), .Q(n7444) );
  MUX21X1 U9765 ( .IN1(\mem1[217][15] ), .IN2(n1022), .S(n7445), .Q(n16251) );
  MUX21X1 U9766 ( .IN1(\mem1[217][14] ), .IN2(n1000), .S(n7445), .Q(n16250) );
  MUX21X1 U9767 ( .IN1(\mem1[217][13] ), .IN2(n978), .S(n7445), .Q(n16249) );
  MUX21X1 U9768 ( .IN1(\mem1[217][12] ), .IN2(n956), .S(n7445), .Q(n16248) );
  MUX21X1 U9769 ( .IN1(\mem1[217][11] ), .IN2(n934), .S(n7445), .Q(n16247) );
  MUX21X1 U9770 ( .IN1(\mem1[217][10] ), .IN2(n912), .S(n7445), .Q(n16246) );
  MUX21X1 U9771 ( .IN1(\mem1[217][9] ), .IN2(n890), .S(n7445), .Q(n16245) );
  MUX21X1 U9772 ( .IN1(\mem1[217][8] ), .IN2(n868), .S(n7445), .Q(n16244) );
  AND2X1 U9773 ( .IN1(n7439), .IN2(n7112), .Q(n7445) );
  MUX21X1 U9774 ( .IN1(\mem1[216][15] ), .IN2(n1022), .S(n7446), .Q(n16243) );
  MUX21X1 U9775 ( .IN1(\mem1[216][14] ), .IN2(n1000), .S(n7446), .Q(n16242) );
  MUX21X1 U9776 ( .IN1(\mem1[216][13] ), .IN2(n978), .S(n7446), .Q(n16241) );
  MUX21X1 U9777 ( .IN1(\mem1[216][12] ), .IN2(n956), .S(n7446), .Q(n16240) );
  MUX21X1 U9778 ( .IN1(\mem1[216][11] ), .IN2(n934), .S(n7446), .Q(n16239) );
  MUX21X1 U9779 ( .IN1(\mem1[216][10] ), .IN2(n912), .S(n7446), .Q(n16238) );
  MUX21X1 U9780 ( .IN1(\mem1[216][9] ), .IN2(n890), .S(n7446), .Q(n16237) );
  MUX21X1 U9781 ( .IN1(\mem1[216][8] ), .IN2(n868), .S(n7446), .Q(n16236) );
  AND2X1 U9782 ( .IN1(n7439), .IN2(n7114), .Q(n7446) );
  MUX21X1 U9783 ( .IN1(\mem1[215][15] ), .IN2(n1022), .S(n7447), .Q(n16235) );
  MUX21X1 U9784 ( .IN1(\mem1[215][14] ), .IN2(n1000), .S(n7447), .Q(n16234) );
  MUX21X1 U9785 ( .IN1(\mem1[215][13] ), .IN2(n978), .S(n7447), .Q(n16233) );
  MUX21X1 U9786 ( .IN1(\mem1[215][12] ), .IN2(n956), .S(n7447), .Q(n16232) );
  MUX21X1 U9787 ( .IN1(\mem1[215][11] ), .IN2(n934), .S(n7447), .Q(n16231) );
  MUX21X1 U9788 ( .IN1(\mem1[215][10] ), .IN2(n912), .S(n7447), .Q(n16230) );
  MUX21X1 U9789 ( .IN1(\mem1[215][9] ), .IN2(n890), .S(n7447), .Q(n16229) );
  MUX21X1 U9790 ( .IN1(\mem1[215][8] ), .IN2(n868), .S(n7447), .Q(n16228) );
  AND2X1 U9791 ( .IN1(n7439), .IN2(n7116), .Q(n7447) );
  MUX21X1 U9792 ( .IN1(\mem1[214][15] ), .IN2(n1022), .S(n7448), .Q(n16227) );
  MUX21X1 U9793 ( .IN1(\mem1[214][14] ), .IN2(n1000), .S(n7448), .Q(n16226) );
  MUX21X1 U9794 ( .IN1(\mem1[214][13] ), .IN2(n978), .S(n7448), .Q(n16225) );
  MUX21X1 U9795 ( .IN1(\mem1[214][12] ), .IN2(n956), .S(n7448), .Q(n16224) );
  MUX21X1 U9796 ( .IN1(\mem1[214][11] ), .IN2(n934), .S(n7448), .Q(n16223) );
  MUX21X1 U9797 ( .IN1(\mem1[214][10] ), .IN2(n912), .S(n7448), .Q(n16222) );
  MUX21X1 U9798 ( .IN1(\mem1[214][9] ), .IN2(n890), .S(n7448), .Q(n16221) );
  MUX21X1 U9799 ( .IN1(\mem1[214][8] ), .IN2(n868), .S(n7448), .Q(n16220) );
  AND2X1 U9800 ( .IN1(n7439), .IN2(n7118), .Q(n7448) );
  MUX21X1 U9801 ( .IN1(\mem1[213][15] ), .IN2(n1022), .S(n7449), .Q(n16219) );
  MUX21X1 U9802 ( .IN1(\mem1[213][14] ), .IN2(n1000), .S(n7449), .Q(n16218) );
  MUX21X1 U9803 ( .IN1(\mem1[213][13] ), .IN2(n978), .S(n7449), .Q(n16217) );
  MUX21X1 U9804 ( .IN1(\mem1[213][12] ), .IN2(n956), .S(n7449), .Q(n16216) );
  MUX21X1 U9805 ( .IN1(\mem1[213][11] ), .IN2(n934), .S(n7449), .Q(n16215) );
  MUX21X1 U9806 ( .IN1(\mem1[213][10] ), .IN2(n912), .S(n7449), .Q(n16214) );
  MUX21X1 U9807 ( .IN1(\mem1[213][9] ), .IN2(n890), .S(n7449), .Q(n16213) );
  MUX21X1 U9808 ( .IN1(\mem1[213][8] ), .IN2(n868), .S(n7449), .Q(n16212) );
  AND2X1 U9809 ( .IN1(n7439), .IN2(n7120), .Q(n7449) );
  MUX21X1 U9810 ( .IN1(\mem1[212][15] ), .IN2(n1022), .S(n7450), .Q(n16211) );
  MUX21X1 U9811 ( .IN1(\mem1[212][14] ), .IN2(n1000), .S(n7450), .Q(n16210) );
  MUX21X1 U9812 ( .IN1(\mem1[212][13] ), .IN2(n978), .S(n7450), .Q(n16209) );
  MUX21X1 U9813 ( .IN1(\mem1[212][12] ), .IN2(n956), .S(n7450), .Q(n16208) );
  MUX21X1 U9814 ( .IN1(\mem1[212][11] ), .IN2(n934), .S(n7450), .Q(n16207) );
  MUX21X1 U9815 ( .IN1(\mem1[212][10] ), .IN2(n912), .S(n7450), .Q(n16206) );
  MUX21X1 U9816 ( .IN1(\mem1[212][9] ), .IN2(n890), .S(n7450), .Q(n16205) );
  MUX21X1 U9817 ( .IN1(\mem1[212][8] ), .IN2(n868), .S(n7450), .Q(n16204) );
  AND2X1 U9818 ( .IN1(n7439), .IN2(n7122), .Q(n7450) );
  MUX21X1 U9819 ( .IN1(\mem1[211][15] ), .IN2(n1022), .S(n7451), .Q(n16203) );
  MUX21X1 U9820 ( .IN1(\mem1[211][14] ), .IN2(n1000), .S(n7451), .Q(n16202) );
  MUX21X1 U9821 ( .IN1(\mem1[211][13] ), .IN2(n978), .S(n7451), .Q(n16201) );
  MUX21X1 U9822 ( .IN1(\mem1[211][12] ), .IN2(n956), .S(n7451), .Q(n16200) );
  MUX21X1 U9823 ( .IN1(\mem1[211][11] ), .IN2(n934), .S(n7451), .Q(n16199) );
  MUX21X1 U9824 ( .IN1(\mem1[211][10] ), .IN2(n912), .S(n7451), .Q(n16198) );
  MUX21X1 U9825 ( .IN1(\mem1[211][9] ), .IN2(n890), .S(n7451), .Q(n16197) );
  MUX21X1 U9826 ( .IN1(\mem1[211][8] ), .IN2(n868), .S(n7451), .Q(n16196) );
  AND2X1 U9827 ( .IN1(n7439), .IN2(n7124), .Q(n7451) );
  MUX21X1 U9828 ( .IN1(\mem1[210][15] ), .IN2(n1022), .S(n7452), .Q(n16195) );
  MUX21X1 U9829 ( .IN1(\mem1[210][14] ), .IN2(n1000), .S(n7452), .Q(n16194) );
  MUX21X1 U9830 ( .IN1(\mem1[210][13] ), .IN2(n978), .S(n7452), .Q(n16193) );
  MUX21X1 U9831 ( .IN1(\mem1[210][12] ), .IN2(n956), .S(n7452), .Q(n16192) );
  MUX21X1 U9832 ( .IN1(\mem1[210][11] ), .IN2(n934), .S(n7452), .Q(n16191) );
  MUX21X1 U9833 ( .IN1(\mem1[210][10] ), .IN2(n912), .S(n7452), .Q(n16190) );
  MUX21X1 U9834 ( .IN1(\mem1[210][9] ), .IN2(n890), .S(n7452), .Q(n16189) );
  MUX21X1 U9835 ( .IN1(\mem1[210][8] ), .IN2(n868), .S(n7452), .Q(n16188) );
  AND2X1 U9836 ( .IN1(n7439), .IN2(n7126), .Q(n7452) );
  MUX21X1 U9837 ( .IN1(\mem1[209][15] ), .IN2(n1022), .S(n7453), .Q(n16187) );
  MUX21X1 U9838 ( .IN1(\mem1[209][14] ), .IN2(n1000), .S(n7453), .Q(n16186) );
  MUX21X1 U9839 ( .IN1(\mem1[209][13] ), .IN2(n978), .S(n7453), .Q(n16185) );
  MUX21X1 U9840 ( .IN1(\mem1[209][12] ), .IN2(n956), .S(n7453), .Q(n16184) );
  MUX21X1 U9841 ( .IN1(\mem1[209][11] ), .IN2(n934), .S(n7453), .Q(n16183) );
  MUX21X1 U9842 ( .IN1(\mem1[209][10] ), .IN2(n912), .S(n7453), .Q(n16182) );
  MUX21X1 U9843 ( .IN1(\mem1[209][9] ), .IN2(n890), .S(n7453), .Q(n16181) );
  MUX21X1 U9844 ( .IN1(\mem1[209][8] ), .IN2(n868), .S(n7453), .Q(n16180) );
  AND2X1 U9845 ( .IN1(n7439), .IN2(n7128), .Q(n7453) );
  MUX21X1 U9846 ( .IN1(\mem1[208][15] ), .IN2(n1022), .S(n7454), .Q(n16179) );
  MUX21X1 U9847 ( .IN1(\mem1[208][14] ), .IN2(n1000), .S(n7454), .Q(n16178) );
  MUX21X1 U9848 ( .IN1(\mem1[208][13] ), .IN2(n978), .S(n7454), .Q(n16177) );
  MUX21X1 U9849 ( .IN1(\mem1[208][12] ), .IN2(n956), .S(n7454), .Q(n16176) );
  MUX21X1 U9850 ( .IN1(\mem1[208][11] ), .IN2(n934), .S(n7454), .Q(n16175) );
  MUX21X1 U9851 ( .IN1(\mem1[208][10] ), .IN2(n912), .S(n7454), .Q(n16174) );
  MUX21X1 U9852 ( .IN1(\mem1[208][9] ), .IN2(n890), .S(n7454), .Q(n16173) );
  MUX21X1 U9853 ( .IN1(\mem1[208][8] ), .IN2(n868), .S(n7454), .Q(n16172) );
  AND2X1 U9854 ( .IN1(n7439), .IN2(n7130), .Q(n7454) );
  AND2X1 U9855 ( .IN1(n7420), .IN2(n7168), .Q(n7439) );
  MUX21X1 U9856 ( .IN1(\mem1[207][15] ), .IN2(n1023), .S(n7455), .Q(n16171) );
  MUX21X1 U9857 ( .IN1(\mem1[207][14] ), .IN2(n1001), .S(n7455), .Q(n16170) );
  MUX21X1 U9858 ( .IN1(\mem1[207][13] ), .IN2(n979), .S(n7455), .Q(n16169) );
  MUX21X1 U9859 ( .IN1(\mem1[207][12] ), .IN2(n957), .S(n7455), .Q(n16168) );
  MUX21X1 U9860 ( .IN1(\mem1[207][11] ), .IN2(n935), .S(n7455), .Q(n16167) );
  MUX21X1 U9861 ( .IN1(\mem1[207][10] ), .IN2(n913), .S(n7455), .Q(n16166) );
  MUX21X1 U9862 ( .IN1(\mem1[207][9] ), .IN2(n891), .S(n7455), .Q(n16165) );
  MUX21X1 U9863 ( .IN1(\mem1[207][8] ), .IN2(n869), .S(n7455), .Q(n16164) );
  AND2X1 U9864 ( .IN1(n7456), .IN2(n7099), .Q(n7455) );
  MUX21X1 U9865 ( .IN1(\mem1[206][15] ), .IN2(n1023), .S(n7457), .Q(n16163) );
  MUX21X1 U9866 ( .IN1(\mem1[206][14] ), .IN2(n1001), .S(n7457), .Q(n16162) );
  MUX21X1 U9867 ( .IN1(\mem1[206][13] ), .IN2(n979), .S(n7457), .Q(n16161) );
  MUX21X1 U9868 ( .IN1(\mem1[206][12] ), .IN2(n957), .S(n7457), .Q(n16160) );
  MUX21X1 U9869 ( .IN1(\mem1[206][11] ), .IN2(n935), .S(n7457), .Q(n16159) );
  MUX21X1 U9870 ( .IN1(\mem1[206][10] ), .IN2(n913), .S(n7457), .Q(n16158) );
  MUX21X1 U9871 ( .IN1(\mem1[206][9] ), .IN2(n891), .S(n7457), .Q(n16157) );
  MUX21X1 U9872 ( .IN1(\mem1[206][8] ), .IN2(n869), .S(n7457), .Q(n16156) );
  AND2X1 U9873 ( .IN1(n7456), .IN2(n7102), .Q(n7457) );
  MUX21X1 U9874 ( .IN1(\mem1[205][15] ), .IN2(n1023), .S(n7458), .Q(n16155) );
  MUX21X1 U9875 ( .IN1(\mem1[205][14] ), .IN2(n1001), .S(n7458), .Q(n16154) );
  MUX21X1 U9876 ( .IN1(\mem1[205][13] ), .IN2(n979), .S(n7458), .Q(n16153) );
  MUX21X1 U9877 ( .IN1(\mem1[205][12] ), .IN2(n957), .S(n7458), .Q(n16152) );
  MUX21X1 U9878 ( .IN1(\mem1[205][11] ), .IN2(n935), .S(n7458), .Q(n16151) );
  MUX21X1 U9879 ( .IN1(\mem1[205][10] ), .IN2(n913), .S(n7458), .Q(n16150) );
  MUX21X1 U9880 ( .IN1(\mem1[205][9] ), .IN2(n891), .S(n7458), .Q(n16149) );
  MUX21X1 U9881 ( .IN1(\mem1[205][8] ), .IN2(n869), .S(n7458), .Q(n16148) );
  AND2X1 U9882 ( .IN1(n7456), .IN2(n7104), .Q(n7458) );
  MUX21X1 U9883 ( .IN1(\mem1[204][15] ), .IN2(n1023), .S(n7459), .Q(n16147) );
  MUX21X1 U9884 ( .IN1(\mem1[204][14] ), .IN2(n1001), .S(n7459), .Q(n16146) );
  MUX21X1 U9885 ( .IN1(\mem1[204][13] ), .IN2(n979), .S(n7459), .Q(n16145) );
  MUX21X1 U9886 ( .IN1(\mem1[204][12] ), .IN2(n957), .S(n7459), .Q(n16144) );
  MUX21X1 U9887 ( .IN1(\mem1[204][11] ), .IN2(n935), .S(n7459), .Q(n16143) );
  MUX21X1 U9888 ( .IN1(\mem1[204][10] ), .IN2(n913), .S(n7459), .Q(n16142) );
  MUX21X1 U9889 ( .IN1(\mem1[204][9] ), .IN2(n891), .S(n7459), .Q(n16141) );
  MUX21X1 U9890 ( .IN1(\mem1[204][8] ), .IN2(n869), .S(n7459), .Q(n16140) );
  AND2X1 U9891 ( .IN1(n7456), .IN2(n7106), .Q(n7459) );
  MUX21X1 U9892 ( .IN1(\mem1[203][15] ), .IN2(n1023), .S(n7460), .Q(n16139) );
  MUX21X1 U9893 ( .IN1(\mem1[203][14] ), .IN2(n1001), .S(n7460), .Q(n16138) );
  MUX21X1 U9894 ( .IN1(\mem1[203][13] ), .IN2(n979), .S(n7460), .Q(n16137) );
  MUX21X1 U9895 ( .IN1(\mem1[203][12] ), .IN2(n957), .S(n7460), .Q(n16136) );
  MUX21X1 U9896 ( .IN1(\mem1[203][11] ), .IN2(n935), .S(n7460), .Q(n16135) );
  MUX21X1 U9897 ( .IN1(\mem1[203][10] ), .IN2(n913), .S(n7460), .Q(n16134) );
  MUX21X1 U9898 ( .IN1(\mem1[203][9] ), .IN2(n891), .S(n7460), .Q(n16133) );
  MUX21X1 U9899 ( .IN1(\mem1[203][8] ), .IN2(n869), .S(n7460), .Q(n16132) );
  AND2X1 U9900 ( .IN1(n7456), .IN2(n7108), .Q(n7460) );
  MUX21X1 U9901 ( .IN1(\mem1[202][15] ), .IN2(n1023), .S(n7461), .Q(n16131) );
  MUX21X1 U9902 ( .IN1(\mem1[202][14] ), .IN2(n1001), .S(n7461), .Q(n16130) );
  MUX21X1 U9903 ( .IN1(\mem1[202][13] ), .IN2(n979), .S(n7461), .Q(n16129) );
  MUX21X1 U9904 ( .IN1(\mem1[202][12] ), .IN2(n957), .S(n7461), .Q(n16128) );
  MUX21X1 U9905 ( .IN1(\mem1[202][11] ), .IN2(n935), .S(n7461), .Q(n16127) );
  MUX21X1 U9906 ( .IN1(\mem1[202][10] ), .IN2(n913), .S(n7461), .Q(n16126) );
  MUX21X1 U9907 ( .IN1(\mem1[202][9] ), .IN2(n891), .S(n7461), .Q(n16125) );
  MUX21X1 U9908 ( .IN1(\mem1[202][8] ), .IN2(n869), .S(n7461), .Q(n16124) );
  AND2X1 U9909 ( .IN1(n7456), .IN2(n7110), .Q(n7461) );
  MUX21X1 U9910 ( .IN1(\mem1[201][15] ), .IN2(n1023), .S(n7462), .Q(n16123) );
  MUX21X1 U9911 ( .IN1(\mem1[201][14] ), .IN2(n1001), .S(n7462), .Q(n16122) );
  MUX21X1 U9912 ( .IN1(\mem1[201][13] ), .IN2(n979), .S(n7462), .Q(n16121) );
  MUX21X1 U9913 ( .IN1(\mem1[201][12] ), .IN2(n957), .S(n7462), .Q(n16120) );
  MUX21X1 U9914 ( .IN1(\mem1[201][11] ), .IN2(n935), .S(n7462), .Q(n16119) );
  MUX21X1 U9915 ( .IN1(\mem1[201][10] ), .IN2(n913), .S(n7462), .Q(n16118) );
  MUX21X1 U9916 ( .IN1(\mem1[201][9] ), .IN2(n891), .S(n7462), .Q(n16117) );
  MUX21X1 U9917 ( .IN1(\mem1[201][8] ), .IN2(n869), .S(n7462), .Q(n16116) );
  AND2X1 U9918 ( .IN1(n7456), .IN2(n7112), .Q(n7462) );
  MUX21X1 U9919 ( .IN1(\mem1[200][15] ), .IN2(n1023), .S(n7463), .Q(n16115) );
  MUX21X1 U9920 ( .IN1(\mem1[200][14] ), .IN2(n1001), .S(n7463), .Q(n16114) );
  MUX21X1 U9921 ( .IN1(\mem1[200][13] ), .IN2(n979), .S(n7463), .Q(n16113) );
  MUX21X1 U9922 ( .IN1(\mem1[200][12] ), .IN2(n957), .S(n7463), .Q(n16112) );
  MUX21X1 U9923 ( .IN1(\mem1[200][11] ), .IN2(n935), .S(n7463), .Q(n16111) );
  MUX21X1 U9924 ( .IN1(\mem1[200][10] ), .IN2(n913), .S(n7463), .Q(n16110) );
  MUX21X1 U9925 ( .IN1(\mem1[200][9] ), .IN2(n891), .S(n7463), .Q(n16109) );
  MUX21X1 U9926 ( .IN1(\mem1[200][8] ), .IN2(n869), .S(n7463), .Q(n16108) );
  AND2X1 U9927 ( .IN1(n7456), .IN2(n7114), .Q(n7463) );
  MUX21X1 U9928 ( .IN1(\mem1[199][15] ), .IN2(n1023), .S(n7464), .Q(n16107) );
  MUX21X1 U9929 ( .IN1(\mem1[199][14] ), .IN2(n1001), .S(n7464), .Q(n16106) );
  MUX21X1 U9930 ( .IN1(\mem1[199][13] ), .IN2(n979), .S(n7464), .Q(n16105) );
  MUX21X1 U9931 ( .IN1(\mem1[199][12] ), .IN2(n957), .S(n7464), .Q(n16104) );
  MUX21X1 U9932 ( .IN1(\mem1[199][11] ), .IN2(n935), .S(n7464), .Q(n16103) );
  MUX21X1 U9933 ( .IN1(\mem1[199][10] ), .IN2(n913), .S(n7464), .Q(n16102) );
  MUX21X1 U9934 ( .IN1(\mem1[199][9] ), .IN2(n891), .S(n7464), .Q(n16101) );
  MUX21X1 U9935 ( .IN1(\mem1[199][8] ), .IN2(n869), .S(n7464), .Q(n16100) );
  AND2X1 U9936 ( .IN1(n7456), .IN2(n7116), .Q(n7464) );
  MUX21X1 U9937 ( .IN1(\mem1[198][15] ), .IN2(n1023), .S(n7465), .Q(n16099) );
  MUX21X1 U9938 ( .IN1(\mem1[198][14] ), .IN2(n1001), .S(n7465), .Q(n16098) );
  MUX21X1 U9939 ( .IN1(\mem1[198][13] ), .IN2(n979), .S(n7465), .Q(n16097) );
  MUX21X1 U9940 ( .IN1(\mem1[198][12] ), .IN2(n957), .S(n7465), .Q(n16096) );
  MUX21X1 U9941 ( .IN1(\mem1[198][11] ), .IN2(n935), .S(n7465), .Q(n16095) );
  MUX21X1 U9942 ( .IN1(\mem1[198][10] ), .IN2(n913), .S(n7465), .Q(n16094) );
  MUX21X1 U9943 ( .IN1(\mem1[198][9] ), .IN2(n891), .S(n7465), .Q(n16093) );
  MUX21X1 U9944 ( .IN1(\mem1[198][8] ), .IN2(n869), .S(n7465), .Q(n16092) );
  AND2X1 U9945 ( .IN1(n7456), .IN2(n7118), .Q(n7465) );
  MUX21X1 U9946 ( .IN1(\mem1[197][15] ), .IN2(n1023), .S(n7466), .Q(n16091) );
  MUX21X1 U9947 ( .IN1(\mem1[197][14] ), .IN2(n1001), .S(n7466), .Q(n16090) );
  MUX21X1 U9948 ( .IN1(\mem1[197][13] ), .IN2(n979), .S(n7466), .Q(n16089) );
  MUX21X1 U9949 ( .IN1(\mem1[197][12] ), .IN2(n957), .S(n7466), .Q(n16088) );
  MUX21X1 U9950 ( .IN1(\mem1[197][11] ), .IN2(n935), .S(n7466), .Q(n16087) );
  MUX21X1 U9951 ( .IN1(\mem1[197][10] ), .IN2(n913), .S(n7466), .Q(n16086) );
  MUX21X1 U9952 ( .IN1(\mem1[197][9] ), .IN2(n891), .S(n7466), .Q(n16085) );
  MUX21X1 U9953 ( .IN1(\mem1[197][8] ), .IN2(n869), .S(n7466), .Q(n16084) );
  AND2X1 U9954 ( .IN1(n7456), .IN2(n7120), .Q(n7466) );
  MUX21X1 U9955 ( .IN1(\mem1[196][15] ), .IN2(n1023), .S(n7467), .Q(n16083) );
  MUX21X1 U9956 ( .IN1(\mem1[196][14] ), .IN2(n1001), .S(n7467), .Q(n16082) );
  MUX21X1 U9957 ( .IN1(\mem1[196][13] ), .IN2(n979), .S(n7467), .Q(n16081) );
  MUX21X1 U9958 ( .IN1(\mem1[196][12] ), .IN2(n957), .S(n7467), .Q(n16080) );
  MUX21X1 U9959 ( .IN1(\mem1[196][11] ), .IN2(n935), .S(n7467), .Q(n16079) );
  MUX21X1 U9960 ( .IN1(\mem1[196][10] ), .IN2(n913), .S(n7467), .Q(n16078) );
  MUX21X1 U9961 ( .IN1(\mem1[196][9] ), .IN2(n891), .S(n7467), .Q(n16077) );
  MUX21X1 U9962 ( .IN1(\mem1[196][8] ), .IN2(n869), .S(n7467), .Q(n16076) );
  AND2X1 U9963 ( .IN1(n7456), .IN2(n7122), .Q(n7467) );
  MUX21X1 U9964 ( .IN1(\mem1[195][15] ), .IN2(n1024), .S(n7468), .Q(n16075) );
  MUX21X1 U9965 ( .IN1(\mem1[195][14] ), .IN2(n1002), .S(n7468), .Q(n16074) );
  MUX21X1 U9966 ( .IN1(\mem1[195][13] ), .IN2(n980), .S(n7468), .Q(n16073) );
  MUX21X1 U9967 ( .IN1(\mem1[195][12] ), .IN2(n958), .S(n7468), .Q(n16072) );
  MUX21X1 U9968 ( .IN1(\mem1[195][11] ), .IN2(n936), .S(n7468), .Q(n16071) );
  MUX21X1 U9969 ( .IN1(\mem1[195][10] ), .IN2(n914), .S(n7468), .Q(n16070) );
  MUX21X1 U9970 ( .IN1(\mem1[195][9] ), .IN2(n892), .S(n7468), .Q(n16069) );
  MUX21X1 U9971 ( .IN1(\mem1[195][8] ), .IN2(n870), .S(n7468), .Q(n16068) );
  AND2X1 U9972 ( .IN1(n7456), .IN2(n7124), .Q(n7468) );
  MUX21X1 U9973 ( .IN1(\mem1[194][15] ), .IN2(n1024), .S(n7469), .Q(n16067) );
  MUX21X1 U9974 ( .IN1(\mem1[194][14] ), .IN2(n1002), .S(n7469), .Q(n16066) );
  MUX21X1 U9975 ( .IN1(\mem1[194][13] ), .IN2(n980), .S(n7469), .Q(n16065) );
  MUX21X1 U9976 ( .IN1(\mem1[194][12] ), .IN2(n958), .S(n7469), .Q(n16064) );
  MUX21X1 U9977 ( .IN1(\mem1[194][11] ), .IN2(n936), .S(n7469), .Q(n16063) );
  MUX21X1 U9978 ( .IN1(\mem1[194][10] ), .IN2(n914), .S(n7469), .Q(n16062) );
  MUX21X1 U9979 ( .IN1(\mem1[194][9] ), .IN2(n892), .S(n7469), .Q(n16061) );
  MUX21X1 U9980 ( .IN1(\mem1[194][8] ), .IN2(n870), .S(n7469), .Q(n16060) );
  AND2X1 U9981 ( .IN1(n7456), .IN2(n7126), .Q(n7469) );
  MUX21X1 U9982 ( .IN1(\mem1[193][15] ), .IN2(n1024), .S(n7470), .Q(n16059) );
  MUX21X1 U9983 ( .IN1(\mem1[193][14] ), .IN2(n1002), .S(n7470), .Q(n16058) );
  MUX21X1 U9984 ( .IN1(\mem1[193][13] ), .IN2(n980), .S(n7470), .Q(n16057) );
  MUX21X1 U9985 ( .IN1(\mem1[193][12] ), .IN2(n958), .S(n7470), .Q(n16056) );
  MUX21X1 U9986 ( .IN1(\mem1[193][11] ), .IN2(n936), .S(n7470), .Q(n16055) );
  MUX21X1 U9987 ( .IN1(\mem1[193][10] ), .IN2(n914), .S(n7470), .Q(n16054) );
  MUX21X1 U9988 ( .IN1(\mem1[193][9] ), .IN2(n892), .S(n7470), .Q(n16053) );
  MUX21X1 U9989 ( .IN1(\mem1[193][8] ), .IN2(n870), .S(n7470), .Q(n16052) );
  AND2X1 U9990 ( .IN1(n7456), .IN2(n7128), .Q(n7470) );
  MUX21X1 U9991 ( .IN1(\mem1[192][15] ), .IN2(n1024), .S(n7471), .Q(n16051) );
  MUX21X1 U9992 ( .IN1(\mem1[192][14] ), .IN2(n1002), .S(n7471), .Q(n16050) );
  MUX21X1 U9993 ( .IN1(\mem1[192][13] ), .IN2(n980), .S(n7471), .Q(n16049) );
  MUX21X1 U9994 ( .IN1(\mem1[192][12] ), .IN2(n958), .S(n7471), .Q(n16048) );
  MUX21X1 U9995 ( .IN1(\mem1[192][11] ), .IN2(n936), .S(n7471), .Q(n16047) );
  MUX21X1 U9996 ( .IN1(\mem1[192][10] ), .IN2(n914), .S(n7471), .Q(n16046) );
  MUX21X1 U9997 ( .IN1(\mem1[192][9] ), .IN2(n892), .S(n7471), .Q(n16045) );
  MUX21X1 U9998 ( .IN1(\mem1[192][8] ), .IN2(n870), .S(n7471), .Q(n16044) );
  AND2X1 U9999 ( .IN1(n7456), .IN2(n7130), .Q(n7471) );
  AND2X1 U10000 ( .IN1(n7420), .IN2(n7186), .Q(n7456) );
  MUX21X1 U10001 ( .IN1(\mem1[191][15] ), .IN2(n1024), .S(n7472), .Q(n16043)
         );
  MUX21X1 U10002 ( .IN1(\mem1[191][14] ), .IN2(n1002), .S(n7472), .Q(n16042)
         );
  MUX21X1 U10003 ( .IN1(\mem1[191][13] ), .IN2(n980), .S(n7472), .Q(n16041) );
  MUX21X1 U10004 ( .IN1(\mem1[191][12] ), .IN2(n958), .S(n7472), .Q(n16040) );
  MUX21X1 U10005 ( .IN1(\mem1[191][11] ), .IN2(n936), .S(n7472), .Q(n16039) );
  MUX21X1 U10006 ( .IN1(\mem1[191][10] ), .IN2(n914), .S(n7472), .Q(n16038) );
  MUX21X1 U10007 ( .IN1(\mem1[191][9] ), .IN2(n892), .S(n7472), .Q(n16037) );
  MUX21X1 U10008 ( .IN1(\mem1[191][8] ), .IN2(n870), .S(n7472), .Q(n16036) );
  AND2X1 U10009 ( .IN1(n7473), .IN2(n7099), .Q(n7472) );
  MUX21X1 U10010 ( .IN1(\mem1[190][15] ), .IN2(n1024), .S(n7474), .Q(n16035)
         );
  MUX21X1 U10011 ( .IN1(\mem1[190][14] ), .IN2(n1002), .S(n7474), .Q(n16034)
         );
  MUX21X1 U10012 ( .IN1(\mem1[190][13] ), .IN2(n980), .S(n7474), .Q(n16033) );
  MUX21X1 U10013 ( .IN1(\mem1[190][12] ), .IN2(n958), .S(n7474), .Q(n16032) );
  MUX21X1 U10014 ( .IN1(\mem1[190][11] ), .IN2(n936), .S(n7474), .Q(n16031) );
  MUX21X1 U10015 ( .IN1(\mem1[190][10] ), .IN2(n914), .S(n7474), .Q(n16030) );
  MUX21X1 U10016 ( .IN1(\mem1[190][9] ), .IN2(n892), .S(n7474), .Q(n16029) );
  MUX21X1 U10017 ( .IN1(\mem1[190][8] ), .IN2(n870), .S(n7474), .Q(n16028) );
  AND2X1 U10018 ( .IN1(n7473), .IN2(n7102), .Q(n7474) );
  MUX21X1 U10019 ( .IN1(\mem1[189][15] ), .IN2(n1024), .S(n7475), .Q(n16027)
         );
  MUX21X1 U10020 ( .IN1(\mem1[189][14] ), .IN2(n1002), .S(n7475), .Q(n16026)
         );
  MUX21X1 U10021 ( .IN1(\mem1[189][13] ), .IN2(n980), .S(n7475), .Q(n16025) );
  MUX21X1 U10022 ( .IN1(\mem1[189][12] ), .IN2(n958), .S(n7475), .Q(n16024) );
  MUX21X1 U10023 ( .IN1(\mem1[189][11] ), .IN2(n936), .S(n7475), .Q(n16023) );
  MUX21X1 U10024 ( .IN1(\mem1[189][10] ), .IN2(n914), .S(n7475), .Q(n16022) );
  MUX21X1 U10025 ( .IN1(\mem1[189][9] ), .IN2(n892), .S(n7475), .Q(n16021) );
  MUX21X1 U10026 ( .IN1(\mem1[189][8] ), .IN2(n870), .S(n7475), .Q(n16020) );
  AND2X1 U10027 ( .IN1(n7473), .IN2(n7104), .Q(n7475) );
  MUX21X1 U10028 ( .IN1(\mem1[188][15] ), .IN2(n1024), .S(n7476), .Q(n16019)
         );
  MUX21X1 U10029 ( .IN1(\mem1[188][14] ), .IN2(n1002), .S(n7476), .Q(n16018)
         );
  MUX21X1 U10030 ( .IN1(\mem1[188][13] ), .IN2(n980), .S(n7476), .Q(n16017) );
  MUX21X1 U10031 ( .IN1(\mem1[188][12] ), .IN2(n958), .S(n7476), .Q(n16016) );
  MUX21X1 U10032 ( .IN1(\mem1[188][11] ), .IN2(n936), .S(n7476), .Q(n16015) );
  MUX21X1 U10033 ( .IN1(\mem1[188][10] ), .IN2(n914), .S(n7476), .Q(n16014) );
  MUX21X1 U10034 ( .IN1(\mem1[188][9] ), .IN2(n892), .S(n7476), .Q(n16013) );
  MUX21X1 U10035 ( .IN1(\mem1[188][8] ), .IN2(n870), .S(n7476), .Q(n16012) );
  AND2X1 U10036 ( .IN1(n7473), .IN2(n7106), .Q(n7476) );
  MUX21X1 U10037 ( .IN1(\mem1[187][15] ), .IN2(n1024), .S(n7477), .Q(n16011)
         );
  MUX21X1 U10038 ( .IN1(\mem1[187][14] ), .IN2(n1002), .S(n7477), .Q(n16010)
         );
  MUX21X1 U10039 ( .IN1(\mem1[187][13] ), .IN2(n980), .S(n7477), .Q(n16009) );
  MUX21X1 U10040 ( .IN1(\mem1[187][12] ), .IN2(n958), .S(n7477), .Q(n16008) );
  MUX21X1 U10041 ( .IN1(\mem1[187][11] ), .IN2(n936), .S(n7477), .Q(n16007) );
  MUX21X1 U10042 ( .IN1(\mem1[187][10] ), .IN2(n914), .S(n7477), .Q(n16006) );
  MUX21X1 U10043 ( .IN1(\mem1[187][9] ), .IN2(n892), .S(n7477), .Q(n16005) );
  MUX21X1 U10044 ( .IN1(\mem1[187][8] ), .IN2(n870), .S(n7477), .Q(n16004) );
  AND2X1 U10045 ( .IN1(n7473), .IN2(n7108), .Q(n7477) );
  MUX21X1 U10046 ( .IN1(\mem1[186][15] ), .IN2(n1024), .S(n7478), .Q(n16003)
         );
  MUX21X1 U10047 ( .IN1(\mem1[186][14] ), .IN2(n1002), .S(n7478), .Q(n16002)
         );
  MUX21X1 U10048 ( .IN1(\mem1[186][13] ), .IN2(n980), .S(n7478), .Q(n16001) );
  MUX21X1 U10049 ( .IN1(\mem1[186][12] ), .IN2(n958), .S(n7478), .Q(n16000) );
  MUX21X1 U10050 ( .IN1(\mem1[186][11] ), .IN2(n936), .S(n7478), .Q(n15999) );
  MUX21X1 U10051 ( .IN1(\mem1[186][10] ), .IN2(n914), .S(n7478), .Q(n15998) );
  MUX21X1 U10052 ( .IN1(\mem1[186][9] ), .IN2(n892), .S(n7478), .Q(n15997) );
  MUX21X1 U10053 ( .IN1(\mem1[186][8] ), .IN2(n870), .S(n7478), .Q(n15996) );
  AND2X1 U10054 ( .IN1(n7473), .IN2(n7110), .Q(n7478) );
  MUX21X1 U10055 ( .IN1(\mem1[185][15] ), .IN2(n1024), .S(n7479), .Q(n15995)
         );
  MUX21X1 U10056 ( .IN1(\mem1[185][14] ), .IN2(n1002), .S(n7479), .Q(n15994)
         );
  MUX21X1 U10057 ( .IN1(\mem1[185][13] ), .IN2(n980), .S(n7479), .Q(n15993) );
  MUX21X1 U10058 ( .IN1(\mem1[185][12] ), .IN2(n958), .S(n7479), .Q(n15992) );
  MUX21X1 U10059 ( .IN1(\mem1[185][11] ), .IN2(n936), .S(n7479), .Q(n15991) );
  MUX21X1 U10060 ( .IN1(\mem1[185][10] ), .IN2(n914), .S(n7479), .Q(n15990) );
  MUX21X1 U10061 ( .IN1(\mem1[185][9] ), .IN2(n892), .S(n7479), .Q(n15989) );
  MUX21X1 U10062 ( .IN1(\mem1[185][8] ), .IN2(n870), .S(n7479), .Q(n15988) );
  AND2X1 U10063 ( .IN1(n7473), .IN2(n7112), .Q(n7479) );
  MUX21X1 U10064 ( .IN1(\mem1[184][15] ), .IN2(n1024), .S(n7480), .Q(n15987)
         );
  MUX21X1 U10065 ( .IN1(\mem1[184][14] ), .IN2(n1002), .S(n7480), .Q(n15986)
         );
  MUX21X1 U10066 ( .IN1(\mem1[184][13] ), .IN2(n980), .S(n7480), .Q(n15985) );
  MUX21X1 U10067 ( .IN1(\mem1[184][12] ), .IN2(n958), .S(n7480), .Q(n15984) );
  MUX21X1 U10068 ( .IN1(\mem1[184][11] ), .IN2(n936), .S(n7480), .Q(n15983) );
  MUX21X1 U10069 ( .IN1(\mem1[184][10] ), .IN2(n914), .S(n7480), .Q(n15982) );
  MUX21X1 U10070 ( .IN1(\mem1[184][9] ), .IN2(n892), .S(n7480), .Q(n15981) );
  MUX21X1 U10071 ( .IN1(\mem1[184][8] ), .IN2(n870), .S(n7480), .Q(n15980) );
  AND2X1 U10072 ( .IN1(n7473), .IN2(n7114), .Q(n7480) );
  MUX21X1 U10073 ( .IN1(\mem1[183][15] ), .IN2(n1025), .S(n7481), .Q(n15979)
         );
  MUX21X1 U10074 ( .IN1(\mem1[183][14] ), .IN2(n1003), .S(n7481), .Q(n15978)
         );
  MUX21X1 U10075 ( .IN1(\mem1[183][13] ), .IN2(n981), .S(n7481), .Q(n15977) );
  MUX21X1 U10076 ( .IN1(\mem1[183][12] ), .IN2(n959), .S(n7481), .Q(n15976) );
  MUX21X1 U10077 ( .IN1(\mem1[183][11] ), .IN2(n937), .S(n7481), .Q(n15975) );
  MUX21X1 U10078 ( .IN1(\mem1[183][10] ), .IN2(n915), .S(n7481), .Q(n15974) );
  MUX21X1 U10079 ( .IN1(\mem1[183][9] ), .IN2(n893), .S(n7481), .Q(n15973) );
  MUX21X1 U10080 ( .IN1(\mem1[183][8] ), .IN2(n871), .S(n7481), .Q(n15972) );
  AND2X1 U10081 ( .IN1(n7473), .IN2(n7116), .Q(n7481) );
  MUX21X1 U10082 ( .IN1(\mem1[182][15] ), .IN2(n1025), .S(n7482), .Q(n15971)
         );
  MUX21X1 U10083 ( .IN1(\mem1[182][14] ), .IN2(n1003), .S(n7482), .Q(n15970)
         );
  MUX21X1 U10084 ( .IN1(\mem1[182][13] ), .IN2(n981), .S(n7482), .Q(n15969) );
  MUX21X1 U10085 ( .IN1(\mem1[182][12] ), .IN2(n959), .S(n7482), .Q(n15968) );
  MUX21X1 U10086 ( .IN1(\mem1[182][11] ), .IN2(n937), .S(n7482), .Q(n15967) );
  MUX21X1 U10087 ( .IN1(\mem1[182][10] ), .IN2(n915), .S(n7482), .Q(n15966) );
  MUX21X1 U10088 ( .IN1(\mem1[182][9] ), .IN2(n893), .S(n7482), .Q(n15965) );
  MUX21X1 U10089 ( .IN1(\mem1[182][8] ), .IN2(n871), .S(n7482), .Q(n15964) );
  AND2X1 U10090 ( .IN1(n7473), .IN2(n7118), .Q(n7482) );
  MUX21X1 U10091 ( .IN1(\mem1[181][15] ), .IN2(n1025), .S(n7483), .Q(n15963)
         );
  MUX21X1 U10092 ( .IN1(\mem1[181][14] ), .IN2(n1003), .S(n7483), .Q(n15962)
         );
  MUX21X1 U10093 ( .IN1(\mem1[181][13] ), .IN2(n981), .S(n7483), .Q(n15961) );
  MUX21X1 U10094 ( .IN1(\mem1[181][12] ), .IN2(n959), .S(n7483), .Q(n15960) );
  MUX21X1 U10095 ( .IN1(\mem1[181][11] ), .IN2(n937), .S(n7483), .Q(n15959) );
  MUX21X1 U10096 ( .IN1(\mem1[181][10] ), .IN2(n915), .S(n7483), .Q(n15958) );
  MUX21X1 U10097 ( .IN1(\mem1[181][9] ), .IN2(n893), .S(n7483), .Q(n15957) );
  MUX21X1 U10098 ( .IN1(\mem1[181][8] ), .IN2(n871), .S(n7483), .Q(n15956) );
  AND2X1 U10099 ( .IN1(n7473), .IN2(n7120), .Q(n7483) );
  MUX21X1 U10100 ( .IN1(\mem1[180][15] ), .IN2(n1025), .S(n7484), .Q(n15955)
         );
  MUX21X1 U10101 ( .IN1(\mem1[180][14] ), .IN2(n1003), .S(n7484), .Q(n15954)
         );
  MUX21X1 U10102 ( .IN1(\mem1[180][13] ), .IN2(n981), .S(n7484), .Q(n15953) );
  MUX21X1 U10103 ( .IN1(\mem1[180][12] ), .IN2(n959), .S(n7484), .Q(n15952) );
  MUX21X1 U10104 ( .IN1(\mem1[180][11] ), .IN2(n937), .S(n7484), .Q(n15951) );
  MUX21X1 U10105 ( .IN1(\mem1[180][10] ), .IN2(n915), .S(n7484), .Q(n15950) );
  MUX21X1 U10106 ( .IN1(\mem1[180][9] ), .IN2(n893), .S(n7484), .Q(n15949) );
  MUX21X1 U10107 ( .IN1(\mem1[180][8] ), .IN2(n871), .S(n7484), .Q(n15948) );
  AND2X1 U10108 ( .IN1(n7473), .IN2(n7122), .Q(n7484) );
  MUX21X1 U10109 ( .IN1(\mem1[179][15] ), .IN2(n1025), .S(n7485), .Q(n15947)
         );
  MUX21X1 U10110 ( .IN1(\mem1[179][14] ), .IN2(n1003), .S(n7485), .Q(n15946)
         );
  MUX21X1 U10111 ( .IN1(\mem1[179][13] ), .IN2(n981), .S(n7485), .Q(n15945) );
  MUX21X1 U10112 ( .IN1(\mem1[179][12] ), .IN2(n959), .S(n7485), .Q(n15944) );
  MUX21X1 U10113 ( .IN1(\mem1[179][11] ), .IN2(n937), .S(n7485), .Q(n15943) );
  MUX21X1 U10114 ( .IN1(\mem1[179][10] ), .IN2(n915), .S(n7485), .Q(n15942) );
  MUX21X1 U10115 ( .IN1(\mem1[179][9] ), .IN2(n893), .S(n7485), .Q(n15941) );
  MUX21X1 U10116 ( .IN1(\mem1[179][8] ), .IN2(n871), .S(n7485), .Q(n15940) );
  AND2X1 U10117 ( .IN1(n7473), .IN2(n7124), .Q(n7485) );
  MUX21X1 U10118 ( .IN1(\mem1[178][15] ), .IN2(n1025), .S(n7486), .Q(n15939)
         );
  MUX21X1 U10119 ( .IN1(\mem1[178][14] ), .IN2(n1003), .S(n7486), .Q(n15938)
         );
  MUX21X1 U10120 ( .IN1(\mem1[178][13] ), .IN2(n981), .S(n7486), .Q(n15937) );
  MUX21X1 U10121 ( .IN1(\mem1[178][12] ), .IN2(n959), .S(n7486), .Q(n15936) );
  MUX21X1 U10122 ( .IN1(\mem1[178][11] ), .IN2(n937), .S(n7486), .Q(n15935) );
  MUX21X1 U10123 ( .IN1(\mem1[178][10] ), .IN2(n915), .S(n7486), .Q(n15934) );
  MUX21X1 U10124 ( .IN1(\mem1[178][9] ), .IN2(n893), .S(n7486), .Q(n15933) );
  MUX21X1 U10125 ( .IN1(\mem1[178][8] ), .IN2(n871), .S(n7486), .Q(n15932) );
  AND2X1 U10126 ( .IN1(n7473), .IN2(n7126), .Q(n7486) );
  MUX21X1 U10127 ( .IN1(\mem1[177][15] ), .IN2(n1025), .S(n7487), .Q(n15931)
         );
  MUX21X1 U10128 ( .IN1(\mem1[177][14] ), .IN2(n1003), .S(n7487), .Q(n15930)
         );
  MUX21X1 U10129 ( .IN1(\mem1[177][13] ), .IN2(n981), .S(n7487), .Q(n15929) );
  MUX21X1 U10130 ( .IN1(\mem1[177][12] ), .IN2(n959), .S(n7487), .Q(n15928) );
  MUX21X1 U10131 ( .IN1(\mem1[177][11] ), .IN2(n937), .S(n7487), .Q(n15927) );
  MUX21X1 U10132 ( .IN1(\mem1[177][10] ), .IN2(n915), .S(n7487), .Q(n15926) );
  MUX21X1 U10133 ( .IN1(\mem1[177][9] ), .IN2(n893), .S(n7487), .Q(n15925) );
  MUX21X1 U10134 ( .IN1(\mem1[177][8] ), .IN2(n871), .S(n7487), .Q(n15924) );
  AND2X1 U10135 ( .IN1(n7473), .IN2(n7128), .Q(n7487) );
  MUX21X1 U10136 ( .IN1(\mem1[176][15] ), .IN2(n1025), .S(n7488), .Q(n15923)
         );
  MUX21X1 U10137 ( .IN1(\mem1[176][14] ), .IN2(n1003), .S(n7488), .Q(n15922)
         );
  MUX21X1 U10138 ( .IN1(\mem1[176][13] ), .IN2(n981), .S(n7488), .Q(n15921) );
  MUX21X1 U10139 ( .IN1(\mem1[176][12] ), .IN2(n959), .S(n7488), .Q(n15920) );
  MUX21X1 U10140 ( .IN1(\mem1[176][11] ), .IN2(n937), .S(n7488), .Q(n15919) );
  MUX21X1 U10141 ( .IN1(\mem1[176][10] ), .IN2(n915), .S(n7488), .Q(n15918) );
  MUX21X1 U10142 ( .IN1(\mem1[176][9] ), .IN2(n893), .S(n7488), .Q(n15917) );
  MUX21X1 U10143 ( .IN1(\mem1[176][8] ), .IN2(n871), .S(n7488), .Q(n15916) );
  AND2X1 U10144 ( .IN1(n7473), .IN2(n7130), .Q(n7488) );
  AND2X1 U10145 ( .IN1(n7420), .IN2(n7204), .Q(n7473) );
  MUX21X1 U10146 ( .IN1(\mem1[175][15] ), .IN2(n1025), .S(n7489), .Q(n15915)
         );
  MUX21X1 U10147 ( .IN1(\mem1[175][14] ), .IN2(n1003), .S(n7489), .Q(n15914)
         );
  MUX21X1 U10148 ( .IN1(\mem1[175][13] ), .IN2(n981), .S(n7489), .Q(n15913) );
  MUX21X1 U10149 ( .IN1(\mem1[175][12] ), .IN2(n959), .S(n7489), .Q(n15912) );
  MUX21X1 U10150 ( .IN1(\mem1[175][11] ), .IN2(n937), .S(n7489), .Q(n15911) );
  MUX21X1 U10151 ( .IN1(\mem1[175][10] ), .IN2(n915), .S(n7489), .Q(n15910) );
  MUX21X1 U10152 ( .IN1(\mem1[175][9] ), .IN2(n893), .S(n7489), .Q(n15909) );
  MUX21X1 U10153 ( .IN1(\mem1[175][8] ), .IN2(n871), .S(n7489), .Q(n15908) );
  AND2X1 U10154 ( .IN1(n7490), .IN2(n7099), .Q(n7489) );
  MUX21X1 U10155 ( .IN1(\mem1[174][15] ), .IN2(n1025), .S(n7491), .Q(n15907)
         );
  MUX21X1 U10156 ( .IN1(\mem1[174][14] ), .IN2(n1003), .S(n7491), .Q(n15906)
         );
  MUX21X1 U10157 ( .IN1(\mem1[174][13] ), .IN2(n981), .S(n7491), .Q(n15905) );
  MUX21X1 U10158 ( .IN1(\mem1[174][12] ), .IN2(n959), .S(n7491), .Q(n15904) );
  MUX21X1 U10159 ( .IN1(\mem1[174][11] ), .IN2(n937), .S(n7491), .Q(n15903) );
  MUX21X1 U10160 ( .IN1(\mem1[174][10] ), .IN2(n915), .S(n7491), .Q(n15902) );
  MUX21X1 U10161 ( .IN1(\mem1[174][9] ), .IN2(n893), .S(n7491), .Q(n15901) );
  MUX21X1 U10162 ( .IN1(\mem1[174][8] ), .IN2(n871), .S(n7491), .Q(n15900) );
  AND2X1 U10163 ( .IN1(n7490), .IN2(n7102), .Q(n7491) );
  MUX21X1 U10164 ( .IN1(\mem1[173][15] ), .IN2(n1025), .S(n7492), .Q(n15899)
         );
  MUX21X1 U10165 ( .IN1(\mem1[173][14] ), .IN2(n1003), .S(n7492), .Q(n15898)
         );
  MUX21X1 U10166 ( .IN1(\mem1[173][13] ), .IN2(n981), .S(n7492), .Q(n15897) );
  MUX21X1 U10167 ( .IN1(\mem1[173][12] ), .IN2(n959), .S(n7492), .Q(n15896) );
  MUX21X1 U10168 ( .IN1(\mem1[173][11] ), .IN2(n937), .S(n7492), .Q(n15895) );
  MUX21X1 U10169 ( .IN1(\mem1[173][10] ), .IN2(n915), .S(n7492), .Q(n15894) );
  MUX21X1 U10170 ( .IN1(\mem1[173][9] ), .IN2(n893), .S(n7492), .Q(n15893) );
  MUX21X1 U10171 ( .IN1(\mem1[173][8] ), .IN2(n871), .S(n7492), .Q(n15892) );
  AND2X1 U10172 ( .IN1(n7490), .IN2(n7104), .Q(n7492) );
  MUX21X1 U10173 ( .IN1(\mem1[172][15] ), .IN2(n1025), .S(n7493), .Q(n15891)
         );
  MUX21X1 U10174 ( .IN1(\mem1[172][14] ), .IN2(n1003), .S(n7493), .Q(n15890)
         );
  MUX21X1 U10175 ( .IN1(\mem1[172][13] ), .IN2(n981), .S(n7493), .Q(n15889) );
  MUX21X1 U10176 ( .IN1(\mem1[172][12] ), .IN2(n959), .S(n7493), .Q(n15888) );
  MUX21X1 U10177 ( .IN1(\mem1[172][11] ), .IN2(n937), .S(n7493), .Q(n15887) );
  MUX21X1 U10178 ( .IN1(\mem1[172][10] ), .IN2(n915), .S(n7493), .Q(n15886) );
  MUX21X1 U10179 ( .IN1(\mem1[172][9] ), .IN2(n893), .S(n7493), .Q(n15885) );
  MUX21X1 U10180 ( .IN1(\mem1[172][8] ), .IN2(n871), .S(n7493), .Q(n15884) );
  AND2X1 U10181 ( .IN1(n7490), .IN2(n7106), .Q(n7493) );
  MUX21X1 U10182 ( .IN1(\mem1[171][15] ), .IN2(n1026), .S(n7494), .Q(n15883)
         );
  MUX21X1 U10183 ( .IN1(\mem1[171][14] ), .IN2(n1004), .S(n7494), .Q(n15882)
         );
  MUX21X1 U10184 ( .IN1(\mem1[171][13] ), .IN2(n982), .S(n7494), .Q(n15881) );
  MUX21X1 U10185 ( .IN1(\mem1[171][12] ), .IN2(n960), .S(n7494), .Q(n15880) );
  MUX21X1 U10186 ( .IN1(\mem1[171][11] ), .IN2(n938), .S(n7494), .Q(n15879) );
  MUX21X1 U10187 ( .IN1(\mem1[171][10] ), .IN2(n916), .S(n7494), .Q(n15878) );
  MUX21X1 U10188 ( .IN1(\mem1[171][9] ), .IN2(n894), .S(n7494), .Q(n15877) );
  MUX21X1 U10189 ( .IN1(\mem1[171][8] ), .IN2(n872), .S(n7494), .Q(n15876) );
  AND2X1 U10190 ( .IN1(n7490), .IN2(n7108), .Q(n7494) );
  MUX21X1 U10191 ( .IN1(\mem1[170][15] ), .IN2(n1026), .S(n7495), .Q(n15875)
         );
  MUX21X1 U10192 ( .IN1(\mem1[170][14] ), .IN2(n1004), .S(n7495), .Q(n15874)
         );
  MUX21X1 U10193 ( .IN1(\mem1[170][13] ), .IN2(n982), .S(n7495), .Q(n15873) );
  MUX21X1 U10194 ( .IN1(\mem1[170][12] ), .IN2(n960), .S(n7495), .Q(n15872) );
  MUX21X1 U10195 ( .IN1(\mem1[170][11] ), .IN2(n938), .S(n7495), .Q(n15871) );
  MUX21X1 U10196 ( .IN1(\mem1[170][10] ), .IN2(n916), .S(n7495), .Q(n15870) );
  MUX21X1 U10197 ( .IN1(\mem1[170][9] ), .IN2(n894), .S(n7495), .Q(n15869) );
  MUX21X1 U10198 ( .IN1(\mem1[170][8] ), .IN2(n872), .S(n7495), .Q(n15868) );
  AND2X1 U10199 ( .IN1(n7490), .IN2(n7110), .Q(n7495) );
  MUX21X1 U10200 ( .IN1(\mem1[169][15] ), .IN2(n1026), .S(n7496), .Q(n15867)
         );
  MUX21X1 U10201 ( .IN1(\mem1[169][14] ), .IN2(n1004), .S(n7496), .Q(n15866)
         );
  MUX21X1 U10202 ( .IN1(\mem1[169][13] ), .IN2(n982), .S(n7496), .Q(n15865) );
  MUX21X1 U10203 ( .IN1(\mem1[169][12] ), .IN2(n960), .S(n7496), .Q(n15864) );
  MUX21X1 U10204 ( .IN1(\mem1[169][11] ), .IN2(n938), .S(n7496), .Q(n15863) );
  MUX21X1 U10205 ( .IN1(\mem1[169][10] ), .IN2(n916), .S(n7496), .Q(n15862) );
  MUX21X1 U10206 ( .IN1(\mem1[169][9] ), .IN2(n894), .S(n7496), .Q(n15861) );
  MUX21X1 U10207 ( .IN1(\mem1[169][8] ), .IN2(n872), .S(n7496), .Q(n15860) );
  AND2X1 U10208 ( .IN1(n7490), .IN2(n7112), .Q(n7496) );
  MUX21X1 U10209 ( .IN1(\mem1[168][15] ), .IN2(n1026), .S(n7497), .Q(n15859)
         );
  MUX21X1 U10210 ( .IN1(\mem1[168][14] ), .IN2(n1004), .S(n7497), .Q(n15858)
         );
  MUX21X1 U10211 ( .IN1(\mem1[168][13] ), .IN2(n982), .S(n7497), .Q(n15857) );
  MUX21X1 U10212 ( .IN1(\mem1[168][12] ), .IN2(n960), .S(n7497), .Q(n15856) );
  MUX21X1 U10213 ( .IN1(\mem1[168][11] ), .IN2(n938), .S(n7497), .Q(n15855) );
  MUX21X1 U10214 ( .IN1(\mem1[168][10] ), .IN2(n916), .S(n7497), .Q(n15854) );
  MUX21X1 U10215 ( .IN1(\mem1[168][9] ), .IN2(n894), .S(n7497), .Q(n15853) );
  MUX21X1 U10216 ( .IN1(\mem1[168][8] ), .IN2(n872), .S(n7497), .Q(n15852) );
  AND2X1 U10217 ( .IN1(n7490), .IN2(n7114), .Q(n7497) );
  MUX21X1 U10218 ( .IN1(\mem1[167][15] ), .IN2(n1026), .S(n7498), .Q(n15851)
         );
  MUX21X1 U10219 ( .IN1(\mem1[167][14] ), .IN2(n1004), .S(n7498), .Q(n15850)
         );
  MUX21X1 U10220 ( .IN1(\mem1[167][13] ), .IN2(n982), .S(n7498), .Q(n15849) );
  MUX21X1 U10221 ( .IN1(\mem1[167][12] ), .IN2(n960), .S(n7498), .Q(n15848) );
  MUX21X1 U10222 ( .IN1(\mem1[167][11] ), .IN2(n938), .S(n7498), .Q(n15847) );
  MUX21X1 U10223 ( .IN1(\mem1[167][10] ), .IN2(n916), .S(n7498), .Q(n15846) );
  MUX21X1 U10224 ( .IN1(\mem1[167][9] ), .IN2(n894), .S(n7498), .Q(n15845) );
  MUX21X1 U10225 ( .IN1(\mem1[167][8] ), .IN2(n872), .S(n7498), .Q(n15844) );
  AND2X1 U10226 ( .IN1(n7490), .IN2(n7116), .Q(n7498) );
  MUX21X1 U10227 ( .IN1(\mem1[166][15] ), .IN2(n1026), .S(n7499), .Q(n15843)
         );
  MUX21X1 U10228 ( .IN1(\mem1[166][14] ), .IN2(n1004), .S(n7499), .Q(n15842)
         );
  MUX21X1 U10229 ( .IN1(\mem1[166][13] ), .IN2(n982), .S(n7499), .Q(n15841) );
  MUX21X1 U10230 ( .IN1(\mem1[166][12] ), .IN2(n960), .S(n7499), .Q(n15840) );
  MUX21X1 U10231 ( .IN1(\mem1[166][11] ), .IN2(n938), .S(n7499), .Q(n15839) );
  MUX21X1 U10232 ( .IN1(\mem1[166][10] ), .IN2(n916), .S(n7499), .Q(n15838) );
  MUX21X1 U10233 ( .IN1(\mem1[166][9] ), .IN2(n894), .S(n7499), .Q(n15837) );
  MUX21X1 U10234 ( .IN1(\mem1[166][8] ), .IN2(n872), .S(n7499), .Q(n15836) );
  AND2X1 U10235 ( .IN1(n7490), .IN2(n7118), .Q(n7499) );
  MUX21X1 U10236 ( .IN1(\mem1[165][15] ), .IN2(n1026), .S(n7500), .Q(n15835)
         );
  MUX21X1 U10237 ( .IN1(\mem1[165][14] ), .IN2(n1004), .S(n7500), .Q(n15834)
         );
  MUX21X1 U10238 ( .IN1(\mem1[165][13] ), .IN2(n982), .S(n7500), .Q(n15833) );
  MUX21X1 U10239 ( .IN1(\mem1[165][12] ), .IN2(n960), .S(n7500), .Q(n15832) );
  MUX21X1 U10240 ( .IN1(\mem1[165][11] ), .IN2(n938), .S(n7500), .Q(n15831) );
  MUX21X1 U10241 ( .IN1(\mem1[165][10] ), .IN2(n916), .S(n7500), .Q(n15830) );
  MUX21X1 U10242 ( .IN1(\mem1[165][9] ), .IN2(n894), .S(n7500), .Q(n15829) );
  MUX21X1 U10243 ( .IN1(\mem1[165][8] ), .IN2(n872), .S(n7500), .Q(n15828) );
  AND2X1 U10244 ( .IN1(n7490), .IN2(n7120), .Q(n7500) );
  MUX21X1 U10245 ( .IN1(\mem1[164][15] ), .IN2(n1026), .S(n7501), .Q(n15827)
         );
  MUX21X1 U10246 ( .IN1(\mem1[164][14] ), .IN2(n1004), .S(n7501), .Q(n15826)
         );
  MUX21X1 U10247 ( .IN1(\mem1[164][13] ), .IN2(n982), .S(n7501), .Q(n15825) );
  MUX21X1 U10248 ( .IN1(\mem1[164][12] ), .IN2(n960), .S(n7501), .Q(n15824) );
  MUX21X1 U10249 ( .IN1(\mem1[164][11] ), .IN2(n938), .S(n7501), .Q(n15823) );
  MUX21X1 U10250 ( .IN1(\mem1[164][10] ), .IN2(n916), .S(n7501), .Q(n15822) );
  MUX21X1 U10251 ( .IN1(\mem1[164][9] ), .IN2(n894), .S(n7501), .Q(n15821) );
  MUX21X1 U10252 ( .IN1(\mem1[164][8] ), .IN2(n872), .S(n7501), .Q(n15820) );
  AND2X1 U10253 ( .IN1(n7490), .IN2(n7122), .Q(n7501) );
  MUX21X1 U10254 ( .IN1(\mem1[163][15] ), .IN2(n1026), .S(n7502), .Q(n15819)
         );
  MUX21X1 U10255 ( .IN1(\mem1[163][14] ), .IN2(n1004), .S(n7502), .Q(n15818)
         );
  MUX21X1 U10256 ( .IN1(\mem1[163][13] ), .IN2(n982), .S(n7502), .Q(n15817) );
  MUX21X1 U10257 ( .IN1(\mem1[163][12] ), .IN2(n960), .S(n7502), .Q(n15816) );
  MUX21X1 U10258 ( .IN1(\mem1[163][11] ), .IN2(n938), .S(n7502), .Q(n15815) );
  MUX21X1 U10259 ( .IN1(\mem1[163][10] ), .IN2(n916), .S(n7502), .Q(n15814) );
  MUX21X1 U10260 ( .IN1(\mem1[163][9] ), .IN2(n894), .S(n7502), .Q(n15813) );
  MUX21X1 U10261 ( .IN1(\mem1[163][8] ), .IN2(n872), .S(n7502), .Q(n15812) );
  AND2X1 U10262 ( .IN1(n7490), .IN2(n7124), .Q(n7502) );
  MUX21X1 U10263 ( .IN1(\mem1[162][15] ), .IN2(n1026), .S(n7503), .Q(n15811)
         );
  MUX21X1 U10264 ( .IN1(\mem1[162][14] ), .IN2(n1004), .S(n7503), .Q(n15810)
         );
  MUX21X1 U10265 ( .IN1(\mem1[162][13] ), .IN2(n982), .S(n7503), .Q(n15809) );
  MUX21X1 U10266 ( .IN1(\mem1[162][12] ), .IN2(n960), .S(n7503), .Q(n15808) );
  MUX21X1 U10267 ( .IN1(\mem1[162][11] ), .IN2(n938), .S(n7503), .Q(n15807) );
  MUX21X1 U10268 ( .IN1(\mem1[162][10] ), .IN2(n916), .S(n7503), .Q(n15806) );
  MUX21X1 U10269 ( .IN1(\mem1[162][9] ), .IN2(n894), .S(n7503), .Q(n15805) );
  MUX21X1 U10270 ( .IN1(\mem1[162][8] ), .IN2(n872), .S(n7503), .Q(n15804) );
  AND2X1 U10271 ( .IN1(n7490), .IN2(n7126), .Q(n7503) );
  MUX21X1 U10272 ( .IN1(\mem1[161][15] ), .IN2(n1026), .S(n7504), .Q(n15803)
         );
  MUX21X1 U10273 ( .IN1(\mem1[161][14] ), .IN2(n1004), .S(n7504), .Q(n15802)
         );
  MUX21X1 U10274 ( .IN1(\mem1[161][13] ), .IN2(n982), .S(n7504), .Q(n15801) );
  MUX21X1 U10275 ( .IN1(\mem1[161][12] ), .IN2(n960), .S(n7504), .Q(n15800) );
  MUX21X1 U10276 ( .IN1(\mem1[161][11] ), .IN2(n938), .S(n7504), .Q(n15799) );
  MUX21X1 U10277 ( .IN1(\mem1[161][10] ), .IN2(n916), .S(n7504), .Q(n15798) );
  MUX21X1 U10278 ( .IN1(\mem1[161][9] ), .IN2(n894), .S(n7504), .Q(n15797) );
  MUX21X1 U10279 ( .IN1(\mem1[161][8] ), .IN2(n872), .S(n7504), .Q(n15796) );
  AND2X1 U10280 ( .IN1(n7490), .IN2(n7128), .Q(n7504) );
  MUX21X1 U10281 ( .IN1(\mem1[160][15] ), .IN2(n1026), .S(n7505), .Q(n15795)
         );
  MUX21X1 U10282 ( .IN1(\mem1[160][14] ), .IN2(n1004), .S(n7505), .Q(n15794)
         );
  MUX21X1 U10283 ( .IN1(\mem1[160][13] ), .IN2(n982), .S(n7505), .Q(n15793) );
  MUX21X1 U10284 ( .IN1(\mem1[160][12] ), .IN2(n960), .S(n7505), .Q(n15792) );
  MUX21X1 U10285 ( .IN1(\mem1[160][11] ), .IN2(n938), .S(n7505), .Q(n15791) );
  MUX21X1 U10286 ( .IN1(\mem1[160][10] ), .IN2(n916), .S(n7505), .Q(n15790) );
  MUX21X1 U10287 ( .IN1(\mem1[160][9] ), .IN2(n894), .S(n7505), .Q(n15789) );
  MUX21X1 U10288 ( .IN1(\mem1[160][8] ), .IN2(n872), .S(n7505), .Q(n15788) );
  AND2X1 U10289 ( .IN1(n7490), .IN2(n7130), .Q(n7505) );
  AND2X1 U10290 ( .IN1(n7420), .IN2(n7222), .Q(n7490) );
  MUX21X1 U10291 ( .IN1(\mem1[159][15] ), .IN2(n1027), .S(n7506), .Q(n15787)
         );
  MUX21X1 U10292 ( .IN1(\mem1[159][14] ), .IN2(n1005), .S(n7506), .Q(n15786)
         );
  MUX21X1 U10293 ( .IN1(\mem1[159][13] ), .IN2(n983), .S(n7506), .Q(n15785) );
  MUX21X1 U10294 ( .IN1(\mem1[159][12] ), .IN2(n961), .S(n7506), .Q(n15784) );
  MUX21X1 U10295 ( .IN1(\mem1[159][11] ), .IN2(n939), .S(n7506), .Q(n15783) );
  MUX21X1 U10296 ( .IN1(\mem1[159][10] ), .IN2(n917), .S(n7506), .Q(n15782) );
  MUX21X1 U10297 ( .IN1(\mem1[159][9] ), .IN2(n895), .S(n7506), .Q(n15781) );
  MUX21X1 U10298 ( .IN1(\mem1[159][8] ), .IN2(n873), .S(n7506), .Q(n15780) );
  AND2X1 U10299 ( .IN1(n7507), .IN2(n7099), .Q(n7506) );
  MUX21X1 U10300 ( .IN1(\mem1[158][15] ), .IN2(n1027), .S(n7508), .Q(n15779)
         );
  MUX21X1 U10301 ( .IN1(\mem1[158][14] ), .IN2(n1005), .S(n7508), .Q(n15778)
         );
  MUX21X1 U10302 ( .IN1(\mem1[158][13] ), .IN2(n983), .S(n7508), .Q(n15777) );
  MUX21X1 U10303 ( .IN1(\mem1[158][12] ), .IN2(n961), .S(n7508), .Q(n15776) );
  MUX21X1 U10304 ( .IN1(\mem1[158][11] ), .IN2(n939), .S(n7508), .Q(n15775) );
  MUX21X1 U10305 ( .IN1(\mem1[158][10] ), .IN2(n917), .S(n7508), .Q(n15774) );
  MUX21X1 U10306 ( .IN1(\mem1[158][9] ), .IN2(n895), .S(n7508), .Q(n15773) );
  MUX21X1 U10307 ( .IN1(\mem1[158][8] ), .IN2(n873), .S(n7508), .Q(n15772) );
  AND2X1 U10308 ( .IN1(n7507), .IN2(n7102), .Q(n7508) );
  MUX21X1 U10309 ( .IN1(\mem1[157][15] ), .IN2(n1027), .S(n7509), .Q(n15771)
         );
  MUX21X1 U10310 ( .IN1(\mem1[157][14] ), .IN2(n1005), .S(n7509), .Q(n15770)
         );
  MUX21X1 U10311 ( .IN1(\mem1[157][13] ), .IN2(n983), .S(n7509), .Q(n15769) );
  MUX21X1 U10312 ( .IN1(\mem1[157][12] ), .IN2(n961), .S(n7509), .Q(n15768) );
  MUX21X1 U10313 ( .IN1(\mem1[157][11] ), .IN2(n939), .S(n7509), .Q(n15767) );
  MUX21X1 U10314 ( .IN1(\mem1[157][10] ), .IN2(n917), .S(n7509), .Q(n15766) );
  MUX21X1 U10315 ( .IN1(\mem1[157][9] ), .IN2(n895), .S(n7509), .Q(n15765) );
  MUX21X1 U10316 ( .IN1(\mem1[157][8] ), .IN2(n873), .S(n7509), .Q(n15764) );
  AND2X1 U10317 ( .IN1(n7507), .IN2(n7104), .Q(n7509) );
  MUX21X1 U10318 ( .IN1(\mem1[156][15] ), .IN2(n1027), .S(n7510), .Q(n15763)
         );
  MUX21X1 U10319 ( .IN1(\mem1[156][14] ), .IN2(n1005), .S(n7510), .Q(n15762)
         );
  MUX21X1 U10320 ( .IN1(\mem1[156][13] ), .IN2(n983), .S(n7510), .Q(n15761) );
  MUX21X1 U10321 ( .IN1(\mem1[156][12] ), .IN2(n961), .S(n7510), .Q(n15760) );
  MUX21X1 U10322 ( .IN1(\mem1[156][11] ), .IN2(n939), .S(n7510), .Q(n15759) );
  MUX21X1 U10323 ( .IN1(\mem1[156][10] ), .IN2(n917), .S(n7510), .Q(n15758) );
  MUX21X1 U10324 ( .IN1(\mem1[156][9] ), .IN2(n895), .S(n7510), .Q(n15757) );
  MUX21X1 U10325 ( .IN1(\mem1[156][8] ), .IN2(n873), .S(n7510), .Q(n15756) );
  AND2X1 U10326 ( .IN1(n7507), .IN2(n7106), .Q(n7510) );
  MUX21X1 U10327 ( .IN1(\mem1[155][15] ), .IN2(n1027), .S(n7511), .Q(n15755)
         );
  MUX21X1 U10328 ( .IN1(\mem1[155][14] ), .IN2(n1005), .S(n7511), .Q(n15754)
         );
  MUX21X1 U10329 ( .IN1(\mem1[155][13] ), .IN2(n983), .S(n7511), .Q(n15753) );
  MUX21X1 U10330 ( .IN1(\mem1[155][12] ), .IN2(n961), .S(n7511), .Q(n15752) );
  MUX21X1 U10331 ( .IN1(\mem1[155][11] ), .IN2(n939), .S(n7511), .Q(n15751) );
  MUX21X1 U10332 ( .IN1(\mem1[155][10] ), .IN2(n917), .S(n7511), .Q(n15750) );
  MUX21X1 U10333 ( .IN1(\mem1[155][9] ), .IN2(n895), .S(n7511), .Q(n15749) );
  MUX21X1 U10334 ( .IN1(\mem1[155][8] ), .IN2(n873), .S(n7511), .Q(n15748) );
  AND2X1 U10335 ( .IN1(n7507), .IN2(n7108), .Q(n7511) );
  MUX21X1 U10336 ( .IN1(\mem1[154][15] ), .IN2(n1027), .S(n7512), .Q(n15747)
         );
  MUX21X1 U10337 ( .IN1(\mem1[154][14] ), .IN2(n1005), .S(n7512), .Q(n15746)
         );
  MUX21X1 U10338 ( .IN1(\mem1[154][13] ), .IN2(n983), .S(n7512), .Q(n15745) );
  MUX21X1 U10339 ( .IN1(\mem1[154][12] ), .IN2(n961), .S(n7512), .Q(n15744) );
  MUX21X1 U10340 ( .IN1(\mem1[154][11] ), .IN2(n939), .S(n7512), .Q(n15743) );
  MUX21X1 U10341 ( .IN1(\mem1[154][10] ), .IN2(n917), .S(n7512), .Q(n15742) );
  MUX21X1 U10342 ( .IN1(\mem1[154][9] ), .IN2(n895), .S(n7512), .Q(n15741) );
  MUX21X1 U10343 ( .IN1(\mem1[154][8] ), .IN2(n873), .S(n7512), .Q(n15740) );
  AND2X1 U10344 ( .IN1(n7507), .IN2(n7110), .Q(n7512) );
  MUX21X1 U10345 ( .IN1(\mem1[153][15] ), .IN2(n1027), .S(n7513), .Q(n15739)
         );
  MUX21X1 U10346 ( .IN1(\mem1[153][14] ), .IN2(n1005), .S(n7513), .Q(n15738)
         );
  MUX21X1 U10347 ( .IN1(\mem1[153][13] ), .IN2(n983), .S(n7513), .Q(n15737) );
  MUX21X1 U10348 ( .IN1(\mem1[153][12] ), .IN2(n961), .S(n7513), .Q(n15736) );
  MUX21X1 U10349 ( .IN1(\mem1[153][11] ), .IN2(n939), .S(n7513), .Q(n15735) );
  MUX21X1 U10350 ( .IN1(\mem1[153][10] ), .IN2(n917), .S(n7513), .Q(n15734) );
  MUX21X1 U10351 ( .IN1(\mem1[153][9] ), .IN2(n895), .S(n7513), .Q(n15733) );
  MUX21X1 U10352 ( .IN1(\mem1[153][8] ), .IN2(n873), .S(n7513), .Q(n15732) );
  AND2X1 U10353 ( .IN1(n7507), .IN2(n7112), .Q(n7513) );
  MUX21X1 U10354 ( .IN1(\mem1[152][15] ), .IN2(n1027), .S(n7514), .Q(n15731)
         );
  MUX21X1 U10355 ( .IN1(\mem1[152][14] ), .IN2(n1005), .S(n7514), .Q(n15730)
         );
  MUX21X1 U10356 ( .IN1(\mem1[152][13] ), .IN2(n983), .S(n7514), .Q(n15729) );
  MUX21X1 U10357 ( .IN1(\mem1[152][12] ), .IN2(n961), .S(n7514), .Q(n15728) );
  MUX21X1 U10358 ( .IN1(\mem1[152][11] ), .IN2(n939), .S(n7514), .Q(n15727) );
  MUX21X1 U10359 ( .IN1(\mem1[152][10] ), .IN2(n917), .S(n7514), .Q(n15726) );
  MUX21X1 U10360 ( .IN1(\mem1[152][9] ), .IN2(n895), .S(n7514), .Q(n15725) );
  MUX21X1 U10361 ( .IN1(\mem1[152][8] ), .IN2(n873), .S(n7514), .Q(n15724) );
  AND2X1 U10362 ( .IN1(n7507), .IN2(n7114), .Q(n7514) );
  MUX21X1 U10363 ( .IN1(\mem1[151][15] ), .IN2(n1027), .S(n7515), .Q(n15723)
         );
  MUX21X1 U10364 ( .IN1(\mem1[151][14] ), .IN2(n1005), .S(n7515), .Q(n15722)
         );
  MUX21X1 U10365 ( .IN1(\mem1[151][13] ), .IN2(n983), .S(n7515), .Q(n15721) );
  MUX21X1 U10366 ( .IN1(\mem1[151][12] ), .IN2(n961), .S(n7515), .Q(n15720) );
  MUX21X1 U10367 ( .IN1(\mem1[151][11] ), .IN2(n939), .S(n7515), .Q(n15719) );
  MUX21X1 U10368 ( .IN1(\mem1[151][10] ), .IN2(n917), .S(n7515), .Q(n15718) );
  MUX21X1 U10369 ( .IN1(\mem1[151][9] ), .IN2(n895), .S(n7515), .Q(n15717) );
  MUX21X1 U10370 ( .IN1(\mem1[151][8] ), .IN2(n873), .S(n7515), .Q(n15716) );
  AND2X1 U10371 ( .IN1(n7507), .IN2(n7116), .Q(n7515) );
  MUX21X1 U10372 ( .IN1(\mem1[150][15] ), .IN2(n1027), .S(n7516), .Q(n15715)
         );
  MUX21X1 U10373 ( .IN1(\mem1[150][14] ), .IN2(n1005), .S(n7516), .Q(n15714)
         );
  MUX21X1 U10374 ( .IN1(\mem1[150][13] ), .IN2(n983), .S(n7516), .Q(n15713) );
  MUX21X1 U10375 ( .IN1(\mem1[150][12] ), .IN2(n961), .S(n7516), .Q(n15712) );
  MUX21X1 U10376 ( .IN1(\mem1[150][11] ), .IN2(n939), .S(n7516), .Q(n15711) );
  MUX21X1 U10377 ( .IN1(\mem1[150][10] ), .IN2(n917), .S(n7516), .Q(n15710) );
  MUX21X1 U10378 ( .IN1(\mem1[150][9] ), .IN2(n895), .S(n7516), .Q(n15709) );
  MUX21X1 U10379 ( .IN1(\mem1[150][8] ), .IN2(n873), .S(n7516), .Q(n15708) );
  AND2X1 U10380 ( .IN1(n7507), .IN2(n7118), .Q(n7516) );
  MUX21X1 U10381 ( .IN1(\mem1[149][15] ), .IN2(n1027), .S(n7517), .Q(n15707)
         );
  MUX21X1 U10382 ( .IN1(\mem1[149][14] ), .IN2(n1005), .S(n7517), .Q(n15706)
         );
  MUX21X1 U10383 ( .IN1(\mem1[149][13] ), .IN2(n983), .S(n7517), .Q(n15705) );
  MUX21X1 U10384 ( .IN1(\mem1[149][12] ), .IN2(n961), .S(n7517), .Q(n15704) );
  MUX21X1 U10385 ( .IN1(\mem1[149][11] ), .IN2(n939), .S(n7517), .Q(n15703) );
  MUX21X1 U10386 ( .IN1(\mem1[149][10] ), .IN2(n917), .S(n7517), .Q(n15702) );
  MUX21X1 U10387 ( .IN1(\mem1[149][9] ), .IN2(n895), .S(n7517), .Q(n15701) );
  MUX21X1 U10388 ( .IN1(\mem1[149][8] ), .IN2(n873), .S(n7517), .Q(n15700) );
  AND2X1 U10389 ( .IN1(n7507), .IN2(n7120), .Q(n7517) );
  MUX21X1 U10390 ( .IN1(\mem1[148][15] ), .IN2(n1027), .S(n7518), .Q(n15699)
         );
  MUX21X1 U10391 ( .IN1(\mem1[148][14] ), .IN2(n1005), .S(n7518), .Q(n15698)
         );
  MUX21X1 U10392 ( .IN1(\mem1[148][13] ), .IN2(n983), .S(n7518), .Q(n15697) );
  MUX21X1 U10393 ( .IN1(\mem1[148][12] ), .IN2(n961), .S(n7518), .Q(n15696) );
  MUX21X1 U10394 ( .IN1(\mem1[148][11] ), .IN2(n939), .S(n7518), .Q(n15695) );
  MUX21X1 U10395 ( .IN1(\mem1[148][10] ), .IN2(n917), .S(n7518), .Q(n15694) );
  MUX21X1 U10396 ( .IN1(\mem1[148][9] ), .IN2(n895), .S(n7518), .Q(n15693) );
  MUX21X1 U10397 ( .IN1(\mem1[148][8] ), .IN2(n873), .S(n7518), .Q(n15692) );
  AND2X1 U10398 ( .IN1(n7507), .IN2(n7122), .Q(n7518) );
  MUX21X1 U10399 ( .IN1(\mem1[147][15] ), .IN2(n1028), .S(n7519), .Q(n15691)
         );
  MUX21X1 U10400 ( .IN1(\mem1[147][14] ), .IN2(n1006), .S(n7519), .Q(n15690)
         );
  MUX21X1 U10401 ( .IN1(\mem1[147][13] ), .IN2(n984), .S(n7519), .Q(n15689) );
  MUX21X1 U10402 ( .IN1(\mem1[147][12] ), .IN2(n962), .S(n7519), .Q(n15688) );
  MUX21X1 U10403 ( .IN1(\mem1[147][11] ), .IN2(n940), .S(n7519), .Q(n15687) );
  MUX21X1 U10404 ( .IN1(\mem1[147][10] ), .IN2(n918), .S(n7519), .Q(n15686) );
  MUX21X1 U10405 ( .IN1(\mem1[147][9] ), .IN2(n896), .S(n7519), .Q(n15685) );
  MUX21X1 U10406 ( .IN1(\mem1[147][8] ), .IN2(n874), .S(n7519), .Q(n15684) );
  AND2X1 U10407 ( .IN1(n7507), .IN2(n7124), .Q(n7519) );
  MUX21X1 U10408 ( .IN1(\mem1[146][15] ), .IN2(n1028), .S(n7520), .Q(n15683)
         );
  MUX21X1 U10409 ( .IN1(\mem1[146][14] ), .IN2(n1006), .S(n7520), .Q(n15682)
         );
  MUX21X1 U10410 ( .IN1(\mem1[146][13] ), .IN2(n984), .S(n7520), .Q(n15681) );
  MUX21X1 U10411 ( .IN1(\mem1[146][12] ), .IN2(n962), .S(n7520), .Q(n15680) );
  MUX21X1 U10412 ( .IN1(\mem1[146][11] ), .IN2(n940), .S(n7520), .Q(n15679) );
  MUX21X1 U10413 ( .IN1(\mem1[146][10] ), .IN2(n918), .S(n7520), .Q(n15678) );
  MUX21X1 U10414 ( .IN1(\mem1[146][9] ), .IN2(n896), .S(n7520), .Q(n15677) );
  MUX21X1 U10415 ( .IN1(\mem1[146][8] ), .IN2(n874), .S(n7520), .Q(n15676) );
  AND2X1 U10416 ( .IN1(n7507), .IN2(n7126), .Q(n7520) );
  MUX21X1 U10417 ( .IN1(\mem1[145][15] ), .IN2(n1028), .S(n7521), .Q(n15675)
         );
  MUX21X1 U10418 ( .IN1(\mem1[145][14] ), .IN2(n1006), .S(n7521), .Q(n15674)
         );
  MUX21X1 U10419 ( .IN1(\mem1[145][13] ), .IN2(n984), .S(n7521), .Q(n15673) );
  MUX21X1 U10420 ( .IN1(\mem1[145][12] ), .IN2(n962), .S(n7521), .Q(n15672) );
  MUX21X1 U10421 ( .IN1(\mem1[145][11] ), .IN2(n940), .S(n7521), .Q(n15671) );
  MUX21X1 U10422 ( .IN1(\mem1[145][10] ), .IN2(n918), .S(n7521), .Q(n15670) );
  MUX21X1 U10423 ( .IN1(\mem1[145][9] ), .IN2(n896), .S(n7521), .Q(n15669) );
  MUX21X1 U10424 ( .IN1(\mem1[145][8] ), .IN2(n874), .S(n7521), .Q(n15668) );
  AND2X1 U10425 ( .IN1(n7507), .IN2(n7128), .Q(n7521) );
  MUX21X1 U10426 ( .IN1(\mem1[144][15] ), .IN2(n1028), .S(n7522), .Q(n15667)
         );
  MUX21X1 U10427 ( .IN1(\mem1[144][14] ), .IN2(n1006), .S(n7522), .Q(n15666)
         );
  MUX21X1 U10428 ( .IN1(\mem1[144][13] ), .IN2(n984), .S(n7522), .Q(n15665) );
  MUX21X1 U10429 ( .IN1(\mem1[144][12] ), .IN2(n962), .S(n7522), .Q(n15664) );
  MUX21X1 U10430 ( .IN1(\mem1[144][11] ), .IN2(n940), .S(n7522), .Q(n15663) );
  MUX21X1 U10431 ( .IN1(\mem1[144][10] ), .IN2(n918), .S(n7522), .Q(n15662) );
  MUX21X1 U10432 ( .IN1(\mem1[144][9] ), .IN2(n896), .S(n7522), .Q(n15661) );
  MUX21X1 U10433 ( .IN1(\mem1[144][8] ), .IN2(n874), .S(n7522), .Q(n15660) );
  AND2X1 U10434 ( .IN1(n7507), .IN2(n7130), .Q(n7522) );
  AND2X1 U10435 ( .IN1(n7420), .IN2(n7240), .Q(n7507) );
  MUX21X1 U10436 ( .IN1(\mem1[143][15] ), .IN2(n1028), .S(n7523), .Q(n15659)
         );
  MUX21X1 U10437 ( .IN1(\mem1[143][14] ), .IN2(n1006), .S(n7523), .Q(n15658)
         );
  MUX21X1 U10438 ( .IN1(\mem1[143][13] ), .IN2(n984), .S(n7523), .Q(n15657) );
  MUX21X1 U10439 ( .IN1(\mem1[143][12] ), .IN2(n962), .S(n7523), .Q(n15656) );
  MUX21X1 U10440 ( .IN1(\mem1[143][11] ), .IN2(n940), .S(n7523), .Q(n15655) );
  MUX21X1 U10441 ( .IN1(\mem1[143][10] ), .IN2(n918), .S(n7523), .Q(n15654) );
  MUX21X1 U10442 ( .IN1(\mem1[143][9] ), .IN2(n896), .S(n7523), .Q(n15653) );
  MUX21X1 U10443 ( .IN1(\mem1[143][8] ), .IN2(n874), .S(n7523), .Q(n15652) );
  AND2X1 U10444 ( .IN1(n7524), .IN2(n7099), .Q(n7523) );
  MUX21X1 U10445 ( .IN1(\mem1[142][15] ), .IN2(n1028), .S(n7525), .Q(n15651)
         );
  MUX21X1 U10446 ( .IN1(\mem1[142][14] ), .IN2(n1006), .S(n7525), .Q(n15650)
         );
  MUX21X1 U10447 ( .IN1(\mem1[142][13] ), .IN2(n984), .S(n7525), .Q(n15649) );
  MUX21X1 U10448 ( .IN1(\mem1[142][12] ), .IN2(n962), .S(n7525), .Q(n15648) );
  MUX21X1 U10449 ( .IN1(\mem1[142][11] ), .IN2(n940), .S(n7525), .Q(n15647) );
  MUX21X1 U10450 ( .IN1(\mem1[142][10] ), .IN2(n918), .S(n7525), .Q(n15646) );
  MUX21X1 U10451 ( .IN1(\mem1[142][9] ), .IN2(n896), .S(n7525), .Q(n15645) );
  MUX21X1 U10452 ( .IN1(\mem1[142][8] ), .IN2(n874), .S(n7525), .Q(n15644) );
  AND2X1 U10453 ( .IN1(n7524), .IN2(n7102), .Q(n7525) );
  MUX21X1 U10454 ( .IN1(\mem1[141][15] ), .IN2(n1028), .S(n7526), .Q(n15643)
         );
  MUX21X1 U10455 ( .IN1(\mem1[141][14] ), .IN2(n1006), .S(n7526), .Q(n15642)
         );
  MUX21X1 U10456 ( .IN1(\mem1[141][13] ), .IN2(n984), .S(n7526), .Q(n15641) );
  MUX21X1 U10457 ( .IN1(\mem1[141][12] ), .IN2(n962), .S(n7526), .Q(n15640) );
  MUX21X1 U10458 ( .IN1(\mem1[141][11] ), .IN2(n940), .S(n7526), .Q(n15639) );
  MUX21X1 U10459 ( .IN1(\mem1[141][10] ), .IN2(n918), .S(n7526), .Q(n15638) );
  MUX21X1 U10460 ( .IN1(\mem1[141][9] ), .IN2(n896), .S(n7526), .Q(n15637) );
  MUX21X1 U10461 ( .IN1(\mem1[141][8] ), .IN2(n874), .S(n7526), .Q(n15636) );
  AND2X1 U10462 ( .IN1(n7524), .IN2(n7104), .Q(n7526) );
  MUX21X1 U10463 ( .IN1(\mem1[140][15] ), .IN2(n1028), .S(n7527), .Q(n15635)
         );
  MUX21X1 U10464 ( .IN1(\mem1[140][14] ), .IN2(n1006), .S(n7527), .Q(n15634)
         );
  MUX21X1 U10465 ( .IN1(\mem1[140][13] ), .IN2(n984), .S(n7527), .Q(n15633) );
  MUX21X1 U10466 ( .IN1(\mem1[140][12] ), .IN2(n962), .S(n7527), .Q(n15632) );
  MUX21X1 U10467 ( .IN1(\mem1[140][11] ), .IN2(n940), .S(n7527), .Q(n15631) );
  MUX21X1 U10468 ( .IN1(\mem1[140][10] ), .IN2(n918), .S(n7527), .Q(n15630) );
  MUX21X1 U10469 ( .IN1(\mem1[140][9] ), .IN2(n896), .S(n7527), .Q(n15629) );
  MUX21X1 U10470 ( .IN1(\mem1[140][8] ), .IN2(n874), .S(n7527), .Q(n15628) );
  AND2X1 U10471 ( .IN1(n7524), .IN2(n7106), .Q(n7527) );
  MUX21X1 U10472 ( .IN1(\mem1[139][15] ), .IN2(n1028), .S(n7528), .Q(n15627)
         );
  MUX21X1 U10473 ( .IN1(\mem1[139][14] ), .IN2(n1006), .S(n7528), .Q(n15626)
         );
  MUX21X1 U10474 ( .IN1(\mem1[139][13] ), .IN2(n984), .S(n7528), .Q(n15625) );
  MUX21X1 U10475 ( .IN1(\mem1[139][12] ), .IN2(n962), .S(n7528), .Q(n15624) );
  MUX21X1 U10476 ( .IN1(\mem1[139][11] ), .IN2(n940), .S(n7528), .Q(n15623) );
  MUX21X1 U10477 ( .IN1(\mem1[139][10] ), .IN2(n918), .S(n7528), .Q(n15622) );
  MUX21X1 U10478 ( .IN1(\mem1[139][9] ), .IN2(n896), .S(n7528), .Q(n15621) );
  MUX21X1 U10479 ( .IN1(\mem1[139][8] ), .IN2(n874), .S(n7528), .Q(n15620) );
  AND2X1 U10480 ( .IN1(n7524), .IN2(n7108), .Q(n7528) );
  MUX21X1 U10481 ( .IN1(\mem1[138][15] ), .IN2(n1028), .S(n7529), .Q(n15619)
         );
  MUX21X1 U10482 ( .IN1(\mem1[138][14] ), .IN2(n1006), .S(n7529), .Q(n15618)
         );
  MUX21X1 U10483 ( .IN1(\mem1[138][13] ), .IN2(n984), .S(n7529), .Q(n15617) );
  MUX21X1 U10484 ( .IN1(\mem1[138][12] ), .IN2(n962), .S(n7529), .Q(n15616) );
  MUX21X1 U10485 ( .IN1(\mem1[138][11] ), .IN2(n940), .S(n7529), .Q(n15615) );
  MUX21X1 U10486 ( .IN1(\mem1[138][10] ), .IN2(n918), .S(n7529), .Q(n15614) );
  MUX21X1 U10487 ( .IN1(\mem1[138][9] ), .IN2(n896), .S(n7529), .Q(n15613) );
  MUX21X1 U10488 ( .IN1(\mem1[138][8] ), .IN2(n874), .S(n7529), .Q(n15612) );
  AND2X1 U10489 ( .IN1(n7524), .IN2(n7110), .Q(n7529) );
  MUX21X1 U10490 ( .IN1(\mem1[137][15] ), .IN2(n1028), .S(n7530), .Q(n15611)
         );
  MUX21X1 U10491 ( .IN1(\mem1[137][14] ), .IN2(n1006), .S(n7530), .Q(n15610)
         );
  MUX21X1 U10492 ( .IN1(\mem1[137][13] ), .IN2(n984), .S(n7530), .Q(n15609) );
  MUX21X1 U10493 ( .IN1(\mem1[137][12] ), .IN2(n962), .S(n7530), .Q(n15608) );
  MUX21X1 U10494 ( .IN1(\mem1[137][11] ), .IN2(n940), .S(n7530), .Q(n15607) );
  MUX21X1 U10495 ( .IN1(\mem1[137][10] ), .IN2(n918), .S(n7530), .Q(n15606) );
  MUX21X1 U10496 ( .IN1(\mem1[137][9] ), .IN2(n896), .S(n7530), .Q(n15605) );
  MUX21X1 U10497 ( .IN1(\mem1[137][8] ), .IN2(n874), .S(n7530), .Q(n15604) );
  AND2X1 U10498 ( .IN1(n7524), .IN2(n7112), .Q(n7530) );
  MUX21X1 U10499 ( .IN1(\mem1[136][15] ), .IN2(n1028), .S(n7531), .Q(n15603)
         );
  MUX21X1 U10500 ( .IN1(\mem1[136][14] ), .IN2(n1006), .S(n7531), .Q(n15602)
         );
  MUX21X1 U10501 ( .IN1(\mem1[136][13] ), .IN2(n984), .S(n7531), .Q(n15601) );
  MUX21X1 U10502 ( .IN1(\mem1[136][12] ), .IN2(n962), .S(n7531), .Q(n15600) );
  MUX21X1 U10503 ( .IN1(\mem1[136][11] ), .IN2(n940), .S(n7531), .Q(n15599) );
  MUX21X1 U10504 ( .IN1(\mem1[136][10] ), .IN2(n918), .S(n7531), .Q(n15598) );
  MUX21X1 U10505 ( .IN1(\mem1[136][9] ), .IN2(n896), .S(n7531), .Q(n15597) );
  MUX21X1 U10506 ( .IN1(\mem1[136][8] ), .IN2(n874), .S(n7531), .Q(n15596) );
  AND2X1 U10507 ( .IN1(n7524), .IN2(n7114), .Q(n7531) );
  MUX21X1 U10508 ( .IN1(\mem1[135][15] ), .IN2(n1029), .S(n7532), .Q(n15595)
         );
  MUX21X1 U10509 ( .IN1(\mem1[135][14] ), .IN2(n1007), .S(n7532), .Q(n15594)
         );
  MUX21X1 U10510 ( .IN1(\mem1[135][13] ), .IN2(n985), .S(n7532), .Q(n15593) );
  MUX21X1 U10511 ( .IN1(\mem1[135][12] ), .IN2(n963), .S(n7532), .Q(n15592) );
  MUX21X1 U10512 ( .IN1(\mem1[135][11] ), .IN2(n941), .S(n7532), .Q(n15591) );
  MUX21X1 U10513 ( .IN1(\mem1[135][10] ), .IN2(n919), .S(n7532), .Q(n15590) );
  MUX21X1 U10514 ( .IN1(\mem1[135][9] ), .IN2(n897), .S(n7532), .Q(n15589) );
  MUX21X1 U10515 ( .IN1(\mem1[135][8] ), .IN2(n875), .S(n7532), .Q(n15588) );
  AND2X1 U10516 ( .IN1(n7524), .IN2(n7116), .Q(n7532) );
  MUX21X1 U10517 ( .IN1(\mem1[134][15] ), .IN2(n1029), .S(n7533), .Q(n15587)
         );
  MUX21X1 U10518 ( .IN1(\mem1[134][14] ), .IN2(n1007), .S(n7533), .Q(n15586)
         );
  MUX21X1 U10519 ( .IN1(\mem1[134][13] ), .IN2(n985), .S(n7533), .Q(n15585) );
  MUX21X1 U10520 ( .IN1(\mem1[134][12] ), .IN2(n963), .S(n7533), .Q(n15584) );
  MUX21X1 U10521 ( .IN1(\mem1[134][11] ), .IN2(n941), .S(n7533), .Q(n15583) );
  MUX21X1 U10522 ( .IN1(\mem1[134][10] ), .IN2(n919), .S(n7533), .Q(n15582) );
  MUX21X1 U10523 ( .IN1(\mem1[134][9] ), .IN2(n897), .S(n7533), .Q(n15581) );
  MUX21X1 U10524 ( .IN1(\mem1[134][8] ), .IN2(n875), .S(n7533), .Q(n15580) );
  AND2X1 U10525 ( .IN1(n7524), .IN2(n7118), .Q(n7533) );
  MUX21X1 U10526 ( .IN1(\mem1[133][15] ), .IN2(n1029), .S(n7534), .Q(n15579)
         );
  MUX21X1 U10527 ( .IN1(\mem1[133][14] ), .IN2(n1007), .S(n7534), .Q(n15578)
         );
  MUX21X1 U10528 ( .IN1(\mem1[133][13] ), .IN2(n985), .S(n7534), .Q(n15577) );
  MUX21X1 U10529 ( .IN1(\mem1[133][12] ), .IN2(n963), .S(n7534), .Q(n15576) );
  MUX21X1 U10530 ( .IN1(\mem1[133][11] ), .IN2(n941), .S(n7534), .Q(n15575) );
  MUX21X1 U10531 ( .IN1(\mem1[133][10] ), .IN2(n919), .S(n7534), .Q(n15574) );
  MUX21X1 U10532 ( .IN1(\mem1[133][9] ), .IN2(n897), .S(n7534), .Q(n15573) );
  MUX21X1 U10533 ( .IN1(\mem1[133][8] ), .IN2(n875), .S(n7534), .Q(n15572) );
  AND2X1 U10534 ( .IN1(n7524), .IN2(n7120), .Q(n7534) );
  MUX21X1 U10535 ( .IN1(\mem1[132][15] ), .IN2(n1029), .S(n7535), .Q(n15571)
         );
  MUX21X1 U10536 ( .IN1(\mem1[132][14] ), .IN2(n1007), .S(n7535), .Q(n15570)
         );
  MUX21X1 U10537 ( .IN1(\mem1[132][13] ), .IN2(n985), .S(n7535), .Q(n15569) );
  MUX21X1 U10538 ( .IN1(\mem1[132][12] ), .IN2(n963), .S(n7535), .Q(n15568) );
  MUX21X1 U10539 ( .IN1(\mem1[132][11] ), .IN2(n941), .S(n7535), .Q(n15567) );
  MUX21X1 U10540 ( .IN1(\mem1[132][10] ), .IN2(n919), .S(n7535), .Q(n15566) );
  MUX21X1 U10541 ( .IN1(\mem1[132][9] ), .IN2(n897), .S(n7535), .Q(n15565) );
  MUX21X1 U10542 ( .IN1(\mem1[132][8] ), .IN2(n875), .S(n7535), .Q(n15564) );
  AND2X1 U10543 ( .IN1(n7524), .IN2(n7122), .Q(n7535) );
  MUX21X1 U10544 ( .IN1(\mem1[131][15] ), .IN2(n1029), .S(n7536), .Q(n15563)
         );
  MUX21X1 U10545 ( .IN1(\mem1[131][14] ), .IN2(n1007), .S(n7536), .Q(n15562)
         );
  MUX21X1 U10546 ( .IN1(\mem1[131][13] ), .IN2(n985), .S(n7536), .Q(n15561) );
  MUX21X1 U10547 ( .IN1(\mem1[131][12] ), .IN2(n963), .S(n7536), .Q(n15560) );
  MUX21X1 U10548 ( .IN1(\mem1[131][11] ), .IN2(n941), .S(n7536), .Q(n15559) );
  MUX21X1 U10549 ( .IN1(\mem1[131][10] ), .IN2(n919), .S(n7536), .Q(n15558) );
  MUX21X1 U10550 ( .IN1(\mem1[131][9] ), .IN2(n897), .S(n7536), .Q(n15557) );
  MUX21X1 U10551 ( .IN1(\mem1[131][8] ), .IN2(n875), .S(n7536), .Q(n15556) );
  AND2X1 U10552 ( .IN1(n7524), .IN2(n7124), .Q(n7536) );
  MUX21X1 U10553 ( .IN1(\mem1[130][15] ), .IN2(n1029), .S(n7537), .Q(n15555)
         );
  MUX21X1 U10554 ( .IN1(\mem1[130][14] ), .IN2(n1007), .S(n7537), .Q(n15554)
         );
  MUX21X1 U10555 ( .IN1(\mem1[130][13] ), .IN2(n985), .S(n7537), .Q(n15553) );
  MUX21X1 U10556 ( .IN1(\mem1[130][12] ), .IN2(n963), .S(n7537), .Q(n15552) );
  MUX21X1 U10557 ( .IN1(\mem1[130][11] ), .IN2(n941), .S(n7537), .Q(n15551) );
  MUX21X1 U10558 ( .IN1(\mem1[130][10] ), .IN2(n919), .S(n7537), .Q(n15550) );
  MUX21X1 U10559 ( .IN1(\mem1[130][9] ), .IN2(n897), .S(n7537), .Q(n15549) );
  MUX21X1 U10560 ( .IN1(\mem1[130][8] ), .IN2(n875), .S(n7537), .Q(n15548) );
  AND2X1 U10561 ( .IN1(n7524), .IN2(n7126), .Q(n7537) );
  MUX21X1 U10562 ( .IN1(\mem1[129][15] ), .IN2(n1029), .S(n7538), .Q(n15547)
         );
  MUX21X1 U10563 ( .IN1(\mem1[129][14] ), .IN2(n1007), .S(n7538), .Q(n15546)
         );
  MUX21X1 U10564 ( .IN1(\mem1[129][13] ), .IN2(n985), .S(n7538), .Q(n15545) );
  MUX21X1 U10565 ( .IN1(\mem1[129][12] ), .IN2(n963), .S(n7538), .Q(n15544) );
  MUX21X1 U10566 ( .IN1(\mem1[129][11] ), .IN2(n941), .S(n7538), .Q(n15543) );
  MUX21X1 U10567 ( .IN1(\mem1[129][10] ), .IN2(n919), .S(n7538), .Q(n15542) );
  MUX21X1 U10568 ( .IN1(\mem1[129][9] ), .IN2(n897), .S(n7538), .Q(n15541) );
  MUX21X1 U10569 ( .IN1(\mem1[129][8] ), .IN2(n875), .S(n7538), .Q(n15540) );
  AND2X1 U10570 ( .IN1(n7524), .IN2(n7128), .Q(n7538) );
  MUX21X1 U10571 ( .IN1(\mem1[128][15] ), .IN2(n1029), .S(n7539), .Q(n15539)
         );
  MUX21X1 U10572 ( .IN1(\mem1[128][14] ), .IN2(n1007), .S(n7539), .Q(n15538)
         );
  MUX21X1 U10573 ( .IN1(\mem1[128][13] ), .IN2(n985), .S(n7539), .Q(n15537) );
  MUX21X1 U10574 ( .IN1(\mem1[128][12] ), .IN2(n963), .S(n7539), .Q(n15536) );
  MUX21X1 U10575 ( .IN1(\mem1[128][11] ), .IN2(n941), .S(n7539), .Q(n15535) );
  MUX21X1 U10576 ( .IN1(\mem1[128][10] ), .IN2(n919), .S(n7539), .Q(n15534) );
  MUX21X1 U10577 ( .IN1(\mem1[128][9] ), .IN2(n897), .S(n7539), .Q(n15533) );
  MUX21X1 U10578 ( .IN1(\mem1[128][8] ), .IN2(n875), .S(n7539), .Q(n15532) );
  AND2X1 U10579 ( .IN1(n7524), .IN2(n7130), .Q(n7539) );
  AND2X1 U10580 ( .IN1(n7420), .IN2(n7258), .Q(n7524) );
  MUX21X1 U10581 ( .IN1(\mem1[127][15] ), .IN2(n1029), .S(n7540), .Q(n15531)
         );
  MUX21X1 U10582 ( .IN1(\mem1[127][14] ), .IN2(n1007), .S(n7540), .Q(n15530)
         );
  MUX21X1 U10583 ( .IN1(\mem1[127][13] ), .IN2(n985), .S(n7540), .Q(n15529) );
  MUX21X1 U10584 ( .IN1(\mem1[127][12] ), .IN2(n963), .S(n7540), .Q(n15528) );
  MUX21X1 U10585 ( .IN1(\mem1[127][11] ), .IN2(n941), .S(n7540), .Q(n15527) );
  MUX21X1 U10586 ( .IN1(\mem1[127][10] ), .IN2(n919), .S(n7540), .Q(n15526) );
  MUX21X1 U10587 ( .IN1(\mem1[127][9] ), .IN2(n897), .S(n7540), .Q(n15525) );
  MUX21X1 U10588 ( .IN1(\mem1[127][8] ), .IN2(n875), .S(n7540), .Q(n15524) );
  AND2X1 U10589 ( .IN1(n7541), .IN2(n7099), .Q(n7540) );
  MUX21X1 U10590 ( .IN1(\mem1[126][15] ), .IN2(n1029), .S(n7542), .Q(n15523)
         );
  MUX21X1 U10591 ( .IN1(\mem1[126][14] ), .IN2(n1007), .S(n7542), .Q(n15522)
         );
  MUX21X1 U10592 ( .IN1(\mem1[126][13] ), .IN2(n985), .S(n7542), .Q(n15521) );
  MUX21X1 U10593 ( .IN1(\mem1[126][12] ), .IN2(n963), .S(n7542), .Q(n15520) );
  MUX21X1 U10594 ( .IN1(\mem1[126][11] ), .IN2(n941), .S(n7542), .Q(n15519) );
  MUX21X1 U10595 ( .IN1(\mem1[126][10] ), .IN2(n919), .S(n7542), .Q(n15518) );
  MUX21X1 U10596 ( .IN1(\mem1[126][9] ), .IN2(n897), .S(n7542), .Q(n15517) );
  MUX21X1 U10597 ( .IN1(\mem1[126][8] ), .IN2(n875), .S(n7542), .Q(n15516) );
  AND2X1 U10598 ( .IN1(n7541), .IN2(n7102), .Q(n7542) );
  MUX21X1 U10599 ( .IN1(\mem1[125][15] ), .IN2(n1029), .S(n7543), .Q(n15515)
         );
  MUX21X1 U10600 ( .IN1(\mem1[125][14] ), .IN2(n1007), .S(n7543), .Q(n15514)
         );
  MUX21X1 U10601 ( .IN1(\mem1[125][13] ), .IN2(n985), .S(n7543), .Q(n15513) );
  MUX21X1 U10602 ( .IN1(\mem1[125][12] ), .IN2(n963), .S(n7543), .Q(n15512) );
  MUX21X1 U10603 ( .IN1(\mem1[125][11] ), .IN2(n941), .S(n7543), .Q(n15511) );
  MUX21X1 U10604 ( .IN1(\mem1[125][10] ), .IN2(n919), .S(n7543), .Q(n15510) );
  MUX21X1 U10605 ( .IN1(\mem1[125][9] ), .IN2(n897), .S(n7543), .Q(n15509) );
  MUX21X1 U10606 ( .IN1(\mem1[125][8] ), .IN2(n875), .S(n7543), .Q(n15508) );
  AND2X1 U10607 ( .IN1(n7541), .IN2(n7104), .Q(n7543) );
  MUX21X1 U10608 ( .IN1(\mem1[124][15] ), .IN2(n1029), .S(n7544), .Q(n15507)
         );
  MUX21X1 U10609 ( .IN1(\mem1[124][14] ), .IN2(n1007), .S(n7544), .Q(n15506)
         );
  MUX21X1 U10610 ( .IN1(\mem1[124][13] ), .IN2(n985), .S(n7544), .Q(n15505) );
  MUX21X1 U10611 ( .IN1(\mem1[124][12] ), .IN2(n963), .S(n7544), .Q(n15504) );
  MUX21X1 U10612 ( .IN1(\mem1[124][11] ), .IN2(n941), .S(n7544), .Q(n15503) );
  MUX21X1 U10613 ( .IN1(\mem1[124][10] ), .IN2(n919), .S(n7544), .Q(n15502) );
  MUX21X1 U10614 ( .IN1(\mem1[124][9] ), .IN2(n897), .S(n7544), .Q(n15501) );
  MUX21X1 U10615 ( .IN1(\mem1[124][8] ), .IN2(n875), .S(n7544), .Q(n15500) );
  AND2X1 U10616 ( .IN1(n7541), .IN2(n7106), .Q(n7544) );
  MUX21X1 U10617 ( .IN1(\mem1[123][15] ), .IN2(n1030), .S(n7545), .Q(n15499)
         );
  MUX21X1 U10618 ( .IN1(\mem1[123][14] ), .IN2(n1008), .S(n7545), .Q(n15498)
         );
  MUX21X1 U10619 ( .IN1(\mem1[123][13] ), .IN2(n986), .S(n7545), .Q(n15497) );
  MUX21X1 U10620 ( .IN1(\mem1[123][12] ), .IN2(n964), .S(n7545), .Q(n15496) );
  MUX21X1 U10621 ( .IN1(\mem1[123][11] ), .IN2(n942), .S(n7545), .Q(n15495) );
  MUX21X1 U10622 ( .IN1(\mem1[123][10] ), .IN2(n920), .S(n7545), .Q(n15494) );
  MUX21X1 U10623 ( .IN1(\mem1[123][9] ), .IN2(n898), .S(n7545), .Q(n15493) );
  MUX21X1 U10624 ( .IN1(\mem1[123][8] ), .IN2(n876), .S(n7545), .Q(n15492) );
  AND2X1 U10625 ( .IN1(n7541), .IN2(n7108), .Q(n7545) );
  MUX21X1 U10626 ( .IN1(\mem1[122][15] ), .IN2(n1030), .S(n7546), .Q(n15491)
         );
  MUX21X1 U10627 ( .IN1(\mem1[122][14] ), .IN2(n1008), .S(n7546), .Q(n15490)
         );
  MUX21X1 U10628 ( .IN1(\mem1[122][13] ), .IN2(n986), .S(n7546), .Q(n15489) );
  MUX21X1 U10629 ( .IN1(\mem1[122][12] ), .IN2(n964), .S(n7546), .Q(n15488) );
  MUX21X1 U10630 ( .IN1(\mem1[122][11] ), .IN2(n942), .S(n7546), .Q(n15487) );
  MUX21X1 U10631 ( .IN1(\mem1[122][10] ), .IN2(n920), .S(n7546), .Q(n15486) );
  MUX21X1 U10632 ( .IN1(\mem1[122][9] ), .IN2(n898), .S(n7546), .Q(n15485) );
  MUX21X1 U10633 ( .IN1(\mem1[122][8] ), .IN2(n876), .S(n7546), .Q(n15484) );
  AND2X1 U10634 ( .IN1(n7541), .IN2(n7110), .Q(n7546) );
  MUX21X1 U10635 ( .IN1(\mem1[121][15] ), .IN2(n1030), .S(n7547), .Q(n15483)
         );
  MUX21X1 U10636 ( .IN1(\mem1[121][14] ), .IN2(n1008), .S(n7547), .Q(n15482)
         );
  MUX21X1 U10637 ( .IN1(\mem1[121][13] ), .IN2(n986), .S(n7547), .Q(n15481) );
  MUX21X1 U10638 ( .IN1(\mem1[121][12] ), .IN2(n964), .S(n7547), .Q(n15480) );
  MUX21X1 U10639 ( .IN1(\mem1[121][11] ), .IN2(n942), .S(n7547), .Q(n15479) );
  MUX21X1 U10640 ( .IN1(\mem1[121][10] ), .IN2(n920), .S(n7547), .Q(n15478) );
  MUX21X1 U10641 ( .IN1(\mem1[121][9] ), .IN2(n898), .S(n7547), .Q(n15477) );
  MUX21X1 U10642 ( .IN1(\mem1[121][8] ), .IN2(n876), .S(n7547), .Q(n15476) );
  AND2X1 U10643 ( .IN1(n7541), .IN2(n7112), .Q(n7547) );
  MUX21X1 U10644 ( .IN1(\mem1[120][15] ), .IN2(n1030), .S(n7548), .Q(n15475)
         );
  MUX21X1 U10645 ( .IN1(\mem1[120][14] ), .IN2(n1008), .S(n7548), .Q(n15474)
         );
  MUX21X1 U10646 ( .IN1(\mem1[120][13] ), .IN2(n986), .S(n7548), .Q(n15473) );
  MUX21X1 U10647 ( .IN1(\mem1[120][12] ), .IN2(n964), .S(n7548), .Q(n15472) );
  MUX21X1 U10648 ( .IN1(\mem1[120][11] ), .IN2(n942), .S(n7548), .Q(n15471) );
  MUX21X1 U10649 ( .IN1(\mem1[120][10] ), .IN2(n920), .S(n7548), .Q(n15470) );
  MUX21X1 U10650 ( .IN1(\mem1[120][9] ), .IN2(n898), .S(n7548), .Q(n15469) );
  MUX21X1 U10651 ( .IN1(\mem1[120][8] ), .IN2(n876), .S(n7548), .Q(n15468) );
  AND2X1 U10652 ( .IN1(n7541), .IN2(n7114), .Q(n7548) );
  MUX21X1 U10653 ( .IN1(\mem1[119][15] ), .IN2(n1030), .S(n7549), .Q(n15467)
         );
  MUX21X1 U10654 ( .IN1(\mem1[119][14] ), .IN2(n1008), .S(n7549), .Q(n15466)
         );
  MUX21X1 U10655 ( .IN1(\mem1[119][13] ), .IN2(n986), .S(n7549), .Q(n15465) );
  MUX21X1 U10656 ( .IN1(\mem1[119][12] ), .IN2(n964), .S(n7549), .Q(n15464) );
  MUX21X1 U10657 ( .IN1(\mem1[119][11] ), .IN2(n942), .S(n7549), .Q(n15463) );
  MUX21X1 U10658 ( .IN1(\mem1[119][10] ), .IN2(n920), .S(n7549), .Q(n15462) );
  MUX21X1 U10659 ( .IN1(\mem1[119][9] ), .IN2(n898), .S(n7549), .Q(n15461) );
  MUX21X1 U10660 ( .IN1(\mem1[119][8] ), .IN2(n876), .S(n7549), .Q(n15460) );
  AND2X1 U10661 ( .IN1(n7541), .IN2(n7116), .Q(n7549) );
  MUX21X1 U10662 ( .IN1(\mem1[118][15] ), .IN2(n1030), .S(n7550), .Q(n15459)
         );
  MUX21X1 U10663 ( .IN1(\mem1[118][14] ), .IN2(n1008), .S(n7550), .Q(n15458)
         );
  MUX21X1 U10664 ( .IN1(\mem1[118][13] ), .IN2(n986), .S(n7550), .Q(n15457) );
  MUX21X1 U10665 ( .IN1(\mem1[118][12] ), .IN2(n964), .S(n7550), .Q(n15456) );
  MUX21X1 U10666 ( .IN1(\mem1[118][11] ), .IN2(n942), .S(n7550), .Q(n15455) );
  MUX21X1 U10667 ( .IN1(\mem1[118][10] ), .IN2(n920), .S(n7550), .Q(n15454) );
  MUX21X1 U10668 ( .IN1(\mem1[118][9] ), .IN2(n898), .S(n7550), .Q(n15453) );
  MUX21X1 U10669 ( .IN1(\mem1[118][8] ), .IN2(n876), .S(n7550), .Q(n15452) );
  AND2X1 U10670 ( .IN1(n7541), .IN2(n7118), .Q(n7550) );
  MUX21X1 U10671 ( .IN1(\mem1[117][15] ), .IN2(n1030), .S(n7551), .Q(n15451)
         );
  MUX21X1 U10672 ( .IN1(\mem1[117][14] ), .IN2(n1008), .S(n7551), .Q(n15450)
         );
  MUX21X1 U10673 ( .IN1(\mem1[117][13] ), .IN2(n986), .S(n7551), .Q(n15449) );
  MUX21X1 U10674 ( .IN1(\mem1[117][12] ), .IN2(n964), .S(n7551), .Q(n15448) );
  MUX21X1 U10675 ( .IN1(\mem1[117][11] ), .IN2(n942), .S(n7551), .Q(n15447) );
  MUX21X1 U10676 ( .IN1(\mem1[117][10] ), .IN2(n920), .S(n7551), .Q(n15446) );
  MUX21X1 U10677 ( .IN1(\mem1[117][9] ), .IN2(n898), .S(n7551), .Q(n15445) );
  MUX21X1 U10678 ( .IN1(\mem1[117][8] ), .IN2(n876), .S(n7551), .Q(n15444) );
  AND2X1 U10679 ( .IN1(n7541), .IN2(n7120), .Q(n7551) );
  MUX21X1 U10680 ( .IN1(\mem1[116][15] ), .IN2(n1030), .S(n7552), .Q(n15443)
         );
  MUX21X1 U10681 ( .IN1(\mem1[116][14] ), .IN2(n1008), .S(n7552), .Q(n15442)
         );
  MUX21X1 U10682 ( .IN1(\mem1[116][13] ), .IN2(n986), .S(n7552), .Q(n15441) );
  MUX21X1 U10683 ( .IN1(\mem1[116][12] ), .IN2(n964), .S(n7552), .Q(n15440) );
  MUX21X1 U10684 ( .IN1(\mem1[116][11] ), .IN2(n942), .S(n7552), .Q(n15439) );
  MUX21X1 U10685 ( .IN1(\mem1[116][10] ), .IN2(n920), .S(n7552), .Q(n15438) );
  MUX21X1 U10686 ( .IN1(\mem1[116][9] ), .IN2(n898), .S(n7552), .Q(n15437) );
  MUX21X1 U10687 ( .IN1(\mem1[116][8] ), .IN2(n876), .S(n7552), .Q(n15436) );
  AND2X1 U10688 ( .IN1(n7541), .IN2(n7122), .Q(n7552) );
  MUX21X1 U10689 ( .IN1(\mem1[115][15] ), .IN2(n1030), .S(n7553), .Q(n15435)
         );
  MUX21X1 U10690 ( .IN1(\mem1[115][14] ), .IN2(n1008), .S(n7553), .Q(n15434)
         );
  MUX21X1 U10691 ( .IN1(\mem1[115][13] ), .IN2(n986), .S(n7553), .Q(n15433) );
  MUX21X1 U10692 ( .IN1(\mem1[115][12] ), .IN2(n964), .S(n7553), .Q(n15432) );
  MUX21X1 U10693 ( .IN1(\mem1[115][11] ), .IN2(n942), .S(n7553), .Q(n15431) );
  MUX21X1 U10694 ( .IN1(\mem1[115][10] ), .IN2(n920), .S(n7553), .Q(n15430) );
  MUX21X1 U10695 ( .IN1(\mem1[115][9] ), .IN2(n898), .S(n7553), .Q(n15429) );
  MUX21X1 U10696 ( .IN1(\mem1[115][8] ), .IN2(n876), .S(n7553), .Q(n15428) );
  AND2X1 U10697 ( .IN1(n7541), .IN2(n7124), .Q(n7553) );
  MUX21X1 U10698 ( .IN1(\mem1[114][15] ), .IN2(n1030), .S(n7554), .Q(n15427)
         );
  MUX21X1 U10699 ( .IN1(\mem1[114][14] ), .IN2(n1008), .S(n7554), .Q(n15426)
         );
  MUX21X1 U10700 ( .IN1(\mem1[114][13] ), .IN2(n986), .S(n7554), .Q(n15425) );
  MUX21X1 U10701 ( .IN1(\mem1[114][12] ), .IN2(n964), .S(n7554), .Q(n15424) );
  MUX21X1 U10702 ( .IN1(\mem1[114][11] ), .IN2(n942), .S(n7554), .Q(n15423) );
  MUX21X1 U10703 ( .IN1(\mem1[114][10] ), .IN2(n920), .S(n7554), .Q(n15422) );
  MUX21X1 U10704 ( .IN1(\mem1[114][9] ), .IN2(n898), .S(n7554), .Q(n15421) );
  MUX21X1 U10705 ( .IN1(\mem1[114][8] ), .IN2(n876), .S(n7554), .Q(n15420) );
  AND2X1 U10706 ( .IN1(n7541), .IN2(n7126), .Q(n7554) );
  MUX21X1 U10707 ( .IN1(\mem1[113][15] ), .IN2(n1030), .S(n7555), .Q(n15419)
         );
  MUX21X1 U10708 ( .IN1(\mem1[113][14] ), .IN2(n1008), .S(n7555), .Q(n15418)
         );
  MUX21X1 U10709 ( .IN1(\mem1[113][13] ), .IN2(n986), .S(n7555), .Q(n15417) );
  MUX21X1 U10710 ( .IN1(\mem1[113][12] ), .IN2(n964), .S(n7555), .Q(n15416) );
  MUX21X1 U10711 ( .IN1(\mem1[113][11] ), .IN2(n942), .S(n7555), .Q(n15415) );
  MUX21X1 U10712 ( .IN1(\mem1[113][10] ), .IN2(n920), .S(n7555), .Q(n15414) );
  MUX21X1 U10713 ( .IN1(\mem1[113][9] ), .IN2(n898), .S(n7555), .Q(n15413) );
  MUX21X1 U10714 ( .IN1(\mem1[113][8] ), .IN2(n876), .S(n7555), .Q(n15412) );
  AND2X1 U10715 ( .IN1(n7541), .IN2(n7128), .Q(n7555) );
  MUX21X1 U10716 ( .IN1(\mem1[112][15] ), .IN2(n1030), .S(n7556), .Q(n15411)
         );
  MUX21X1 U10717 ( .IN1(\mem1[112][14] ), .IN2(n1008), .S(n7556), .Q(n15410)
         );
  MUX21X1 U10718 ( .IN1(\mem1[112][13] ), .IN2(n986), .S(n7556), .Q(n15409) );
  MUX21X1 U10719 ( .IN1(\mem1[112][12] ), .IN2(n964), .S(n7556), .Q(n15408) );
  MUX21X1 U10720 ( .IN1(\mem1[112][11] ), .IN2(n942), .S(n7556), .Q(n15407) );
  MUX21X1 U10721 ( .IN1(\mem1[112][10] ), .IN2(n920), .S(n7556), .Q(n15406) );
  MUX21X1 U10722 ( .IN1(\mem1[112][9] ), .IN2(n898), .S(n7556), .Q(n15405) );
  MUX21X1 U10723 ( .IN1(\mem1[112][8] ), .IN2(n876), .S(n7556), .Q(n15404) );
  AND2X1 U10724 ( .IN1(n7541), .IN2(n7130), .Q(n7556) );
  AND2X1 U10725 ( .IN1(n7420), .IN2(n7276), .Q(n7541) );
  MUX21X1 U10726 ( .IN1(\mem1[111][15] ), .IN2(n1031), .S(n7557), .Q(n15403)
         );
  MUX21X1 U10727 ( .IN1(\mem1[111][14] ), .IN2(n1009), .S(n7557), .Q(n15402)
         );
  MUX21X1 U10728 ( .IN1(\mem1[111][13] ), .IN2(n987), .S(n7557), .Q(n15401) );
  MUX21X1 U10729 ( .IN1(\mem1[111][12] ), .IN2(n965), .S(n7557), .Q(n15400) );
  MUX21X1 U10730 ( .IN1(\mem1[111][11] ), .IN2(n943), .S(n7557), .Q(n15399) );
  MUX21X1 U10731 ( .IN1(\mem1[111][10] ), .IN2(n921), .S(n7557), .Q(n15398) );
  MUX21X1 U10732 ( .IN1(\mem1[111][9] ), .IN2(n899), .S(n7557), .Q(n15397) );
  MUX21X1 U10733 ( .IN1(\mem1[111][8] ), .IN2(n877), .S(n7557), .Q(n15396) );
  AND2X1 U10734 ( .IN1(n7558), .IN2(n7099), .Q(n7557) );
  MUX21X1 U10735 ( .IN1(\mem1[110][15] ), .IN2(n1031), .S(n7559), .Q(n15395)
         );
  MUX21X1 U10736 ( .IN1(\mem1[110][14] ), .IN2(n1009), .S(n7559), .Q(n15394)
         );
  MUX21X1 U10737 ( .IN1(\mem1[110][13] ), .IN2(n987), .S(n7559), .Q(n15393) );
  MUX21X1 U10738 ( .IN1(\mem1[110][12] ), .IN2(n965), .S(n7559), .Q(n15392) );
  MUX21X1 U10739 ( .IN1(\mem1[110][11] ), .IN2(n943), .S(n7559), .Q(n15391) );
  MUX21X1 U10740 ( .IN1(\mem1[110][10] ), .IN2(n921), .S(n7559), .Q(n15390) );
  MUX21X1 U10741 ( .IN1(\mem1[110][9] ), .IN2(n899), .S(n7559), .Q(n15389) );
  MUX21X1 U10742 ( .IN1(\mem1[110][8] ), .IN2(n877), .S(n7559), .Q(n15388) );
  AND2X1 U10743 ( .IN1(n7558), .IN2(n7102), .Q(n7559) );
  MUX21X1 U10744 ( .IN1(\mem1[109][15] ), .IN2(n1031), .S(n7560), .Q(n15387)
         );
  MUX21X1 U10745 ( .IN1(\mem1[109][14] ), .IN2(n1009), .S(n7560), .Q(n15386)
         );
  MUX21X1 U10746 ( .IN1(\mem1[109][13] ), .IN2(n987), .S(n7560), .Q(n15385) );
  MUX21X1 U10747 ( .IN1(\mem1[109][12] ), .IN2(n965), .S(n7560), .Q(n15384) );
  MUX21X1 U10748 ( .IN1(\mem1[109][11] ), .IN2(n943), .S(n7560), .Q(n15383) );
  MUX21X1 U10749 ( .IN1(\mem1[109][10] ), .IN2(n921), .S(n7560), .Q(n15382) );
  MUX21X1 U10750 ( .IN1(\mem1[109][9] ), .IN2(n899), .S(n7560), .Q(n15381) );
  MUX21X1 U10751 ( .IN1(\mem1[109][8] ), .IN2(n877), .S(n7560), .Q(n15380) );
  AND2X1 U10752 ( .IN1(n7558), .IN2(n7104), .Q(n7560) );
  MUX21X1 U10753 ( .IN1(\mem1[108][15] ), .IN2(n1031), .S(n7561), .Q(n15379)
         );
  MUX21X1 U10754 ( .IN1(\mem1[108][14] ), .IN2(n1009), .S(n7561), .Q(n15378)
         );
  MUX21X1 U10755 ( .IN1(\mem1[108][13] ), .IN2(n987), .S(n7561), .Q(n15377) );
  MUX21X1 U10756 ( .IN1(\mem1[108][12] ), .IN2(n965), .S(n7561), .Q(n15376) );
  MUX21X1 U10757 ( .IN1(\mem1[108][11] ), .IN2(n943), .S(n7561), .Q(n15375) );
  MUX21X1 U10758 ( .IN1(\mem1[108][10] ), .IN2(n921), .S(n7561), .Q(n15374) );
  MUX21X1 U10759 ( .IN1(\mem1[108][9] ), .IN2(n899), .S(n7561), .Q(n15373) );
  MUX21X1 U10760 ( .IN1(\mem1[108][8] ), .IN2(n877), .S(n7561), .Q(n15372) );
  AND2X1 U10761 ( .IN1(n7558), .IN2(n7106), .Q(n7561) );
  MUX21X1 U10762 ( .IN1(\mem1[107][15] ), .IN2(n1031), .S(n7562), .Q(n15371)
         );
  MUX21X1 U10763 ( .IN1(\mem1[107][14] ), .IN2(n1009), .S(n7562), .Q(n15370)
         );
  MUX21X1 U10764 ( .IN1(\mem1[107][13] ), .IN2(n987), .S(n7562), .Q(n15369) );
  MUX21X1 U10765 ( .IN1(\mem1[107][12] ), .IN2(n965), .S(n7562), .Q(n15368) );
  MUX21X1 U10766 ( .IN1(\mem1[107][11] ), .IN2(n943), .S(n7562), .Q(n15367) );
  MUX21X1 U10767 ( .IN1(\mem1[107][10] ), .IN2(n921), .S(n7562), .Q(n15366) );
  MUX21X1 U10768 ( .IN1(\mem1[107][9] ), .IN2(n899), .S(n7562), .Q(n15365) );
  MUX21X1 U10769 ( .IN1(\mem1[107][8] ), .IN2(n877), .S(n7562), .Q(n15364) );
  AND2X1 U10770 ( .IN1(n7558), .IN2(n7108), .Q(n7562) );
  MUX21X1 U10771 ( .IN1(\mem1[106][15] ), .IN2(n1031), .S(n7563), .Q(n15363)
         );
  MUX21X1 U10772 ( .IN1(\mem1[106][14] ), .IN2(n1009), .S(n7563), .Q(n15362)
         );
  MUX21X1 U10773 ( .IN1(\mem1[106][13] ), .IN2(n987), .S(n7563), .Q(n15361) );
  MUX21X1 U10774 ( .IN1(\mem1[106][12] ), .IN2(n965), .S(n7563), .Q(n15360) );
  MUX21X1 U10775 ( .IN1(\mem1[106][11] ), .IN2(n943), .S(n7563), .Q(n15359) );
  MUX21X1 U10776 ( .IN1(\mem1[106][10] ), .IN2(n921), .S(n7563), .Q(n15358) );
  MUX21X1 U10777 ( .IN1(\mem1[106][9] ), .IN2(n899), .S(n7563), .Q(n15357) );
  MUX21X1 U10778 ( .IN1(\mem1[106][8] ), .IN2(n877), .S(n7563), .Q(n15356) );
  AND2X1 U10779 ( .IN1(n7558), .IN2(n7110), .Q(n7563) );
  MUX21X1 U10780 ( .IN1(\mem1[105][15] ), .IN2(n1031), .S(n7564), .Q(n15355)
         );
  MUX21X1 U10781 ( .IN1(\mem1[105][14] ), .IN2(n1009), .S(n7564), .Q(n15354)
         );
  MUX21X1 U10782 ( .IN1(\mem1[105][13] ), .IN2(n987), .S(n7564), .Q(n15353) );
  MUX21X1 U10783 ( .IN1(\mem1[105][12] ), .IN2(n965), .S(n7564), .Q(n15352) );
  MUX21X1 U10784 ( .IN1(\mem1[105][11] ), .IN2(n943), .S(n7564), .Q(n15351) );
  MUX21X1 U10785 ( .IN1(\mem1[105][10] ), .IN2(n921), .S(n7564), .Q(n15350) );
  MUX21X1 U10786 ( .IN1(\mem1[105][9] ), .IN2(n899), .S(n7564), .Q(n15349) );
  MUX21X1 U10787 ( .IN1(\mem1[105][8] ), .IN2(n877), .S(n7564), .Q(n15348) );
  AND2X1 U10788 ( .IN1(n7558), .IN2(n7112), .Q(n7564) );
  MUX21X1 U10789 ( .IN1(\mem1[104][15] ), .IN2(n1031), .S(n7565), .Q(n15347)
         );
  MUX21X1 U10790 ( .IN1(\mem1[104][14] ), .IN2(n1009), .S(n7565), .Q(n15346)
         );
  MUX21X1 U10791 ( .IN1(\mem1[104][13] ), .IN2(n987), .S(n7565), .Q(n15345) );
  MUX21X1 U10792 ( .IN1(\mem1[104][12] ), .IN2(n965), .S(n7565), .Q(n15344) );
  MUX21X1 U10793 ( .IN1(\mem1[104][11] ), .IN2(n943), .S(n7565), .Q(n15343) );
  MUX21X1 U10794 ( .IN1(\mem1[104][10] ), .IN2(n921), .S(n7565), .Q(n15342) );
  MUX21X1 U10795 ( .IN1(\mem1[104][9] ), .IN2(n899), .S(n7565), .Q(n15341) );
  MUX21X1 U10796 ( .IN1(\mem1[104][8] ), .IN2(n877), .S(n7565), .Q(n15340) );
  AND2X1 U10797 ( .IN1(n7558), .IN2(n7114), .Q(n7565) );
  MUX21X1 U10798 ( .IN1(\mem1[103][15] ), .IN2(n1031), .S(n7566), .Q(n15339)
         );
  MUX21X1 U10799 ( .IN1(\mem1[103][14] ), .IN2(n1009), .S(n7566), .Q(n15338)
         );
  MUX21X1 U10800 ( .IN1(\mem1[103][13] ), .IN2(n987), .S(n7566), .Q(n15337) );
  MUX21X1 U10801 ( .IN1(\mem1[103][12] ), .IN2(n965), .S(n7566), .Q(n15336) );
  MUX21X1 U10802 ( .IN1(\mem1[103][11] ), .IN2(n943), .S(n7566), .Q(n15335) );
  MUX21X1 U10803 ( .IN1(\mem1[103][10] ), .IN2(n921), .S(n7566), .Q(n15334) );
  MUX21X1 U10804 ( .IN1(\mem1[103][9] ), .IN2(n899), .S(n7566), .Q(n15333) );
  MUX21X1 U10805 ( .IN1(\mem1[103][8] ), .IN2(n877), .S(n7566), .Q(n15332) );
  AND2X1 U10806 ( .IN1(n7558), .IN2(n7116), .Q(n7566) );
  MUX21X1 U10807 ( .IN1(\mem1[102][15] ), .IN2(n1031), .S(n7567), .Q(n15331)
         );
  MUX21X1 U10808 ( .IN1(\mem1[102][14] ), .IN2(n1009), .S(n7567), .Q(n15330)
         );
  MUX21X1 U10809 ( .IN1(\mem1[102][13] ), .IN2(n987), .S(n7567), .Q(n15329) );
  MUX21X1 U10810 ( .IN1(\mem1[102][12] ), .IN2(n965), .S(n7567), .Q(n15328) );
  MUX21X1 U10811 ( .IN1(\mem1[102][11] ), .IN2(n943), .S(n7567), .Q(n15327) );
  MUX21X1 U10812 ( .IN1(\mem1[102][10] ), .IN2(n921), .S(n7567), .Q(n15326) );
  MUX21X1 U10813 ( .IN1(\mem1[102][9] ), .IN2(n899), .S(n7567), .Q(n15325) );
  MUX21X1 U10814 ( .IN1(\mem1[102][8] ), .IN2(n877), .S(n7567), .Q(n15324) );
  AND2X1 U10815 ( .IN1(n7558), .IN2(n7118), .Q(n7567) );
  MUX21X1 U10816 ( .IN1(\mem1[101][15] ), .IN2(n1031), .S(n7568), .Q(n15323)
         );
  MUX21X1 U10817 ( .IN1(\mem1[101][14] ), .IN2(n1009), .S(n7568), .Q(n15322)
         );
  MUX21X1 U10818 ( .IN1(\mem1[101][13] ), .IN2(n987), .S(n7568), .Q(n15321) );
  MUX21X1 U10819 ( .IN1(\mem1[101][12] ), .IN2(n965), .S(n7568), .Q(n15320) );
  MUX21X1 U10820 ( .IN1(\mem1[101][11] ), .IN2(n943), .S(n7568), .Q(n15319) );
  MUX21X1 U10821 ( .IN1(\mem1[101][10] ), .IN2(n921), .S(n7568), .Q(n15318) );
  MUX21X1 U10822 ( .IN1(\mem1[101][9] ), .IN2(n899), .S(n7568), .Q(n15317) );
  MUX21X1 U10823 ( .IN1(\mem1[101][8] ), .IN2(n877), .S(n7568), .Q(n15316) );
  AND2X1 U10824 ( .IN1(n7558), .IN2(n7120), .Q(n7568) );
  MUX21X1 U10825 ( .IN1(\mem1[100][15] ), .IN2(n1031), .S(n7569), .Q(n15315)
         );
  MUX21X1 U10826 ( .IN1(\mem1[100][14] ), .IN2(n1009), .S(n7569), .Q(n15314)
         );
  MUX21X1 U10827 ( .IN1(\mem1[100][13] ), .IN2(n987), .S(n7569), .Q(n15313) );
  MUX21X1 U10828 ( .IN1(\mem1[100][12] ), .IN2(n965), .S(n7569), .Q(n15312) );
  MUX21X1 U10829 ( .IN1(\mem1[100][11] ), .IN2(n943), .S(n7569), .Q(n15311) );
  MUX21X1 U10830 ( .IN1(\mem1[100][10] ), .IN2(n921), .S(n7569), .Q(n15310) );
  MUX21X1 U10831 ( .IN1(\mem1[100][9] ), .IN2(n899), .S(n7569), .Q(n15309) );
  MUX21X1 U10832 ( .IN1(\mem1[100][8] ), .IN2(n877), .S(n7569), .Q(n15308) );
  AND2X1 U10833 ( .IN1(n7558), .IN2(n7122), .Q(n7569) );
  MUX21X1 U10834 ( .IN1(\mem1[99][15] ), .IN2(n1032), .S(n7570), .Q(n15307) );
  MUX21X1 U10835 ( .IN1(\mem1[99][14] ), .IN2(n1010), .S(n7570), .Q(n15306) );
  MUX21X1 U10836 ( .IN1(\mem1[99][13] ), .IN2(n988), .S(n7570), .Q(n15305) );
  MUX21X1 U10837 ( .IN1(\mem1[99][12] ), .IN2(n966), .S(n7570), .Q(n15304) );
  MUX21X1 U10838 ( .IN1(\mem1[99][11] ), .IN2(n944), .S(n7570), .Q(n15303) );
  MUX21X1 U10839 ( .IN1(\mem1[99][10] ), .IN2(n922), .S(n7570), .Q(n15302) );
  MUX21X1 U10840 ( .IN1(\mem1[99][9] ), .IN2(n900), .S(n7570), .Q(n15301) );
  MUX21X1 U10841 ( .IN1(\mem1[99][8] ), .IN2(n878), .S(n7570), .Q(n15300) );
  AND2X1 U10842 ( .IN1(n7558), .IN2(n7124), .Q(n7570) );
  MUX21X1 U10843 ( .IN1(\mem1[98][15] ), .IN2(n1032), .S(n7571), .Q(n15299) );
  MUX21X1 U10844 ( .IN1(\mem1[98][14] ), .IN2(n1010), .S(n7571), .Q(n15298) );
  MUX21X1 U10845 ( .IN1(\mem1[98][13] ), .IN2(n988), .S(n7571), .Q(n15297) );
  MUX21X1 U10846 ( .IN1(\mem1[98][12] ), .IN2(n966), .S(n7571), .Q(n15296) );
  MUX21X1 U10847 ( .IN1(\mem1[98][11] ), .IN2(n944), .S(n7571), .Q(n15295) );
  MUX21X1 U10848 ( .IN1(\mem1[98][10] ), .IN2(n922), .S(n7571), .Q(n15294) );
  MUX21X1 U10849 ( .IN1(\mem1[98][9] ), .IN2(n900), .S(n7571), .Q(n15293) );
  MUX21X1 U10850 ( .IN1(\mem1[98][8] ), .IN2(n878), .S(n7571), .Q(n15292) );
  AND2X1 U10851 ( .IN1(n7558), .IN2(n7126), .Q(n7571) );
  MUX21X1 U10852 ( .IN1(\mem1[97][15] ), .IN2(n1032), .S(n7572), .Q(n15291) );
  MUX21X1 U10853 ( .IN1(\mem1[97][14] ), .IN2(n1010), .S(n7572), .Q(n15290) );
  MUX21X1 U10854 ( .IN1(\mem1[97][13] ), .IN2(n988), .S(n7572), .Q(n15289) );
  MUX21X1 U10855 ( .IN1(\mem1[97][12] ), .IN2(n966), .S(n7572), .Q(n15288) );
  MUX21X1 U10856 ( .IN1(\mem1[97][11] ), .IN2(n944), .S(n7572), .Q(n15287) );
  MUX21X1 U10857 ( .IN1(\mem1[97][10] ), .IN2(n922), .S(n7572), .Q(n15286) );
  MUX21X1 U10858 ( .IN1(\mem1[97][9] ), .IN2(n900), .S(n7572), .Q(n15285) );
  MUX21X1 U10859 ( .IN1(\mem1[97][8] ), .IN2(n878), .S(n7572), .Q(n15284) );
  AND2X1 U10860 ( .IN1(n7558), .IN2(n7128), .Q(n7572) );
  MUX21X1 U10861 ( .IN1(\mem1[96][15] ), .IN2(n1032), .S(n7573), .Q(n15283) );
  MUX21X1 U10862 ( .IN1(\mem1[96][14] ), .IN2(n1010), .S(n7573), .Q(n15282) );
  MUX21X1 U10863 ( .IN1(\mem1[96][13] ), .IN2(n988), .S(n7573), .Q(n15281) );
  MUX21X1 U10864 ( .IN1(\mem1[96][12] ), .IN2(n966), .S(n7573), .Q(n15280) );
  MUX21X1 U10865 ( .IN1(\mem1[96][11] ), .IN2(n944), .S(n7573), .Q(n15279) );
  MUX21X1 U10866 ( .IN1(\mem1[96][10] ), .IN2(n922), .S(n7573), .Q(n15278) );
  MUX21X1 U10867 ( .IN1(\mem1[96][9] ), .IN2(n900), .S(n7573), .Q(n15277) );
  MUX21X1 U10868 ( .IN1(\mem1[96][8] ), .IN2(n878), .S(n7573), .Q(n15276) );
  AND2X1 U10869 ( .IN1(n7558), .IN2(n7130), .Q(n7573) );
  AND2X1 U10870 ( .IN1(n7420), .IN2(n7294), .Q(n7558) );
  MUX21X1 U10871 ( .IN1(\mem1[95][15] ), .IN2(n1032), .S(n7574), .Q(n15275) );
  MUX21X1 U10872 ( .IN1(\mem1[95][14] ), .IN2(n1010), .S(n7574), .Q(n15274) );
  MUX21X1 U10873 ( .IN1(\mem1[95][13] ), .IN2(n988), .S(n7574), .Q(n15273) );
  MUX21X1 U10874 ( .IN1(\mem1[95][12] ), .IN2(n966), .S(n7574), .Q(n15272) );
  MUX21X1 U10875 ( .IN1(\mem1[95][11] ), .IN2(n944), .S(n7574), .Q(n15271) );
  MUX21X1 U10876 ( .IN1(\mem1[95][10] ), .IN2(n922), .S(n7574), .Q(n15270) );
  MUX21X1 U10877 ( .IN1(\mem1[95][9] ), .IN2(n900), .S(n7574), .Q(n15269) );
  MUX21X1 U10878 ( .IN1(\mem1[95][8] ), .IN2(n878), .S(n7574), .Q(n15268) );
  AND2X1 U10879 ( .IN1(n7575), .IN2(n7099), .Q(n7574) );
  MUX21X1 U10880 ( .IN1(\mem1[94][15] ), .IN2(n1032), .S(n7576), .Q(n15267) );
  MUX21X1 U10881 ( .IN1(\mem1[94][14] ), .IN2(n1010), .S(n7576), .Q(n15266) );
  MUX21X1 U10882 ( .IN1(\mem1[94][13] ), .IN2(n988), .S(n7576), .Q(n15265) );
  MUX21X1 U10883 ( .IN1(\mem1[94][12] ), .IN2(n966), .S(n7576), .Q(n15264) );
  MUX21X1 U10884 ( .IN1(\mem1[94][11] ), .IN2(n944), .S(n7576), .Q(n15263) );
  MUX21X1 U10885 ( .IN1(\mem1[94][10] ), .IN2(n922), .S(n7576), .Q(n15262) );
  MUX21X1 U10886 ( .IN1(\mem1[94][9] ), .IN2(n900), .S(n7576), .Q(n15261) );
  MUX21X1 U10887 ( .IN1(\mem1[94][8] ), .IN2(n878), .S(n7576), .Q(n15260) );
  AND2X1 U10888 ( .IN1(n7575), .IN2(n7102), .Q(n7576) );
  MUX21X1 U10889 ( .IN1(\mem1[93][15] ), .IN2(n1032), .S(n7577), .Q(n15259) );
  MUX21X1 U10890 ( .IN1(\mem1[93][14] ), .IN2(n1010), .S(n7577), .Q(n15258) );
  MUX21X1 U10891 ( .IN1(\mem1[93][13] ), .IN2(n988), .S(n7577), .Q(n15257) );
  MUX21X1 U10892 ( .IN1(\mem1[93][12] ), .IN2(n966), .S(n7577), .Q(n15256) );
  MUX21X1 U10893 ( .IN1(\mem1[93][11] ), .IN2(n944), .S(n7577), .Q(n15255) );
  MUX21X1 U10894 ( .IN1(\mem1[93][10] ), .IN2(n922), .S(n7577), .Q(n15254) );
  MUX21X1 U10895 ( .IN1(\mem1[93][9] ), .IN2(n900), .S(n7577), .Q(n15253) );
  MUX21X1 U10896 ( .IN1(\mem1[93][8] ), .IN2(n878), .S(n7577), .Q(n15252) );
  AND2X1 U10897 ( .IN1(n7575), .IN2(n7104), .Q(n7577) );
  MUX21X1 U10898 ( .IN1(\mem1[92][15] ), .IN2(n1032), .S(n7578), .Q(n15251) );
  MUX21X1 U10899 ( .IN1(\mem1[92][14] ), .IN2(n1010), .S(n7578), .Q(n15250) );
  MUX21X1 U10900 ( .IN1(\mem1[92][13] ), .IN2(n988), .S(n7578), .Q(n15249) );
  MUX21X1 U10901 ( .IN1(\mem1[92][12] ), .IN2(n966), .S(n7578), .Q(n15248) );
  MUX21X1 U10902 ( .IN1(\mem1[92][11] ), .IN2(n944), .S(n7578), .Q(n15247) );
  MUX21X1 U10903 ( .IN1(\mem1[92][10] ), .IN2(n922), .S(n7578), .Q(n15246) );
  MUX21X1 U10904 ( .IN1(\mem1[92][9] ), .IN2(n900), .S(n7578), .Q(n15245) );
  MUX21X1 U10905 ( .IN1(\mem1[92][8] ), .IN2(n878), .S(n7578), .Q(n15244) );
  AND2X1 U10906 ( .IN1(n7575), .IN2(n7106), .Q(n7578) );
  MUX21X1 U10907 ( .IN1(\mem1[91][15] ), .IN2(n1032), .S(n7579), .Q(n15243) );
  MUX21X1 U10908 ( .IN1(\mem1[91][14] ), .IN2(n1010), .S(n7579), .Q(n15242) );
  MUX21X1 U10909 ( .IN1(\mem1[91][13] ), .IN2(n988), .S(n7579), .Q(n15241) );
  MUX21X1 U10910 ( .IN1(\mem1[91][12] ), .IN2(n966), .S(n7579), .Q(n15240) );
  MUX21X1 U10911 ( .IN1(\mem1[91][11] ), .IN2(n944), .S(n7579), .Q(n15239) );
  MUX21X1 U10912 ( .IN1(\mem1[91][10] ), .IN2(n922), .S(n7579), .Q(n15238) );
  MUX21X1 U10913 ( .IN1(\mem1[91][9] ), .IN2(n900), .S(n7579), .Q(n15237) );
  MUX21X1 U10914 ( .IN1(\mem1[91][8] ), .IN2(n878), .S(n7579), .Q(n15236) );
  AND2X1 U10915 ( .IN1(n7575), .IN2(n7108), .Q(n7579) );
  MUX21X1 U10916 ( .IN1(\mem1[90][15] ), .IN2(n1032), .S(n7580), .Q(n15235) );
  MUX21X1 U10917 ( .IN1(\mem1[90][14] ), .IN2(n1010), .S(n7580), .Q(n15234) );
  MUX21X1 U10918 ( .IN1(\mem1[90][13] ), .IN2(n988), .S(n7580), .Q(n15233) );
  MUX21X1 U10919 ( .IN1(\mem1[90][12] ), .IN2(n966), .S(n7580), .Q(n15232) );
  MUX21X1 U10920 ( .IN1(\mem1[90][11] ), .IN2(n944), .S(n7580), .Q(n15231) );
  MUX21X1 U10921 ( .IN1(\mem1[90][10] ), .IN2(n922), .S(n7580), .Q(n15230) );
  MUX21X1 U10922 ( .IN1(\mem1[90][9] ), .IN2(n900), .S(n7580), .Q(n15229) );
  MUX21X1 U10923 ( .IN1(\mem1[90][8] ), .IN2(n878), .S(n7580), .Q(n15228) );
  AND2X1 U10924 ( .IN1(n7575), .IN2(n7110), .Q(n7580) );
  MUX21X1 U10925 ( .IN1(\mem1[89][15] ), .IN2(n1032), .S(n7581), .Q(n15227) );
  MUX21X1 U10926 ( .IN1(\mem1[89][14] ), .IN2(n1010), .S(n7581), .Q(n15226) );
  MUX21X1 U10927 ( .IN1(\mem1[89][13] ), .IN2(n988), .S(n7581), .Q(n15225) );
  MUX21X1 U10928 ( .IN1(\mem1[89][12] ), .IN2(n966), .S(n7581), .Q(n15224) );
  MUX21X1 U10929 ( .IN1(\mem1[89][11] ), .IN2(n944), .S(n7581), .Q(n15223) );
  MUX21X1 U10930 ( .IN1(\mem1[89][10] ), .IN2(n922), .S(n7581), .Q(n15222) );
  MUX21X1 U10931 ( .IN1(\mem1[89][9] ), .IN2(n900), .S(n7581), .Q(n15221) );
  MUX21X1 U10932 ( .IN1(\mem1[89][8] ), .IN2(n878), .S(n7581), .Q(n15220) );
  AND2X1 U10933 ( .IN1(n7575), .IN2(n7112), .Q(n7581) );
  MUX21X1 U10934 ( .IN1(\mem1[88][15] ), .IN2(n1032), .S(n7582), .Q(n15219) );
  MUX21X1 U10935 ( .IN1(\mem1[88][14] ), .IN2(n1010), .S(n7582), .Q(n15218) );
  MUX21X1 U10936 ( .IN1(\mem1[88][13] ), .IN2(n988), .S(n7582), .Q(n15217) );
  MUX21X1 U10937 ( .IN1(\mem1[88][12] ), .IN2(n966), .S(n7582), .Q(n15216) );
  MUX21X1 U10938 ( .IN1(\mem1[88][11] ), .IN2(n944), .S(n7582), .Q(n15215) );
  MUX21X1 U10939 ( .IN1(\mem1[88][10] ), .IN2(n922), .S(n7582), .Q(n15214) );
  MUX21X1 U10940 ( .IN1(\mem1[88][9] ), .IN2(n900), .S(n7582), .Q(n15213) );
  MUX21X1 U10941 ( .IN1(\mem1[88][8] ), .IN2(n878), .S(n7582), .Q(n15212) );
  AND2X1 U10942 ( .IN1(n7575), .IN2(n7114), .Q(n7582) );
  MUX21X1 U10943 ( .IN1(\mem1[87][15] ), .IN2(n1033), .S(n7583), .Q(n15211) );
  MUX21X1 U10944 ( .IN1(\mem1[87][14] ), .IN2(n1011), .S(n7583), .Q(n15210) );
  MUX21X1 U10945 ( .IN1(\mem1[87][13] ), .IN2(n989), .S(n7583), .Q(n15209) );
  MUX21X1 U10946 ( .IN1(\mem1[87][12] ), .IN2(n967), .S(n7583), .Q(n15208) );
  MUX21X1 U10947 ( .IN1(\mem1[87][11] ), .IN2(n945), .S(n7583), .Q(n15207) );
  MUX21X1 U10948 ( .IN1(\mem1[87][10] ), .IN2(n923), .S(n7583), .Q(n15206) );
  MUX21X1 U10949 ( .IN1(\mem1[87][9] ), .IN2(n901), .S(n7583), .Q(n15205) );
  MUX21X1 U10950 ( .IN1(\mem1[87][8] ), .IN2(n879), .S(n7583), .Q(n15204) );
  AND2X1 U10951 ( .IN1(n7575), .IN2(n7116), .Q(n7583) );
  MUX21X1 U10952 ( .IN1(\mem1[86][15] ), .IN2(n1033), .S(n7584), .Q(n15203) );
  MUX21X1 U10953 ( .IN1(\mem1[86][14] ), .IN2(n1011), .S(n7584), .Q(n15202) );
  MUX21X1 U10954 ( .IN1(\mem1[86][13] ), .IN2(n989), .S(n7584), .Q(n15201) );
  MUX21X1 U10955 ( .IN1(\mem1[86][12] ), .IN2(n967), .S(n7584), .Q(n15200) );
  MUX21X1 U10956 ( .IN1(\mem1[86][11] ), .IN2(n945), .S(n7584), .Q(n15199) );
  MUX21X1 U10957 ( .IN1(\mem1[86][10] ), .IN2(n923), .S(n7584), .Q(n15198) );
  MUX21X1 U10958 ( .IN1(\mem1[86][9] ), .IN2(n901), .S(n7584), .Q(n15197) );
  MUX21X1 U10959 ( .IN1(\mem1[86][8] ), .IN2(n879), .S(n7584), .Q(n15196) );
  AND2X1 U10960 ( .IN1(n7575), .IN2(n7118), .Q(n7584) );
  MUX21X1 U10961 ( .IN1(\mem1[85][15] ), .IN2(n1033), .S(n7585), .Q(n15195) );
  MUX21X1 U10962 ( .IN1(\mem1[85][14] ), .IN2(n1011), .S(n7585), .Q(n15194) );
  MUX21X1 U10963 ( .IN1(\mem1[85][13] ), .IN2(n989), .S(n7585), .Q(n15193) );
  MUX21X1 U10964 ( .IN1(\mem1[85][12] ), .IN2(n967), .S(n7585), .Q(n15192) );
  MUX21X1 U10965 ( .IN1(\mem1[85][11] ), .IN2(n945), .S(n7585), .Q(n15191) );
  MUX21X1 U10966 ( .IN1(\mem1[85][10] ), .IN2(n923), .S(n7585), .Q(n15190) );
  MUX21X1 U10967 ( .IN1(\mem1[85][9] ), .IN2(n901), .S(n7585), .Q(n15189) );
  MUX21X1 U10968 ( .IN1(\mem1[85][8] ), .IN2(n879), .S(n7585), .Q(n15188) );
  AND2X1 U10969 ( .IN1(n7575), .IN2(n7120), .Q(n7585) );
  MUX21X1 U10970 ( .IN1(\mem1[84][15] ), .IN2(n1033), .S(n7586), .Q(n15187) );
  MUX21X1 U10971 ( .IN1(\mem1[84][14] ), .IN2(n1011), .S(n7586), .Q(n15186) );
  MUX21X1 U10972 ( .IN1(\mem1[84][13] ), .IN2(n989), .S(n7586), .Q(n15185) );
  MUX21X1 U10973 ( .IN1(\mem1[84][12] ), .IN2(n967), .S(n7586), .Q(n15184) );
  MUX21X1 U10974 ( .IN1(\mem1[84][11] ), .IN2(n945), .S(n7586), .Q(n15183) );
  MUX21X1 U10975 ( .IN1(\mem1[84][10] ), .IN2(n923), .S(n7586), .Q(n15182) );
  MUX21X1 U10976 ( .IN1(\mem1[84][9] ), .IN2(n901), .S(n7586), .Q(n15181) );
  MUX21X1 U10977 ( .IN1(\mem1[84][8] ), .IN2(n879), .S(n7586), .Q(n15180) );
  AND2X1 U10978 ( .IN1(n7575), .IN2(n7122), .Q(n7586) );
  MUX21X1 U10979 ( .IN1(\mem1[83][15] ), .IN2(n1033), .S(n7587), .Q(n15179) );
  MUX21X1 U10980 ( .IN1(\mem1[83][14] ), .IN2(n1011), .S(n7587), .Q(n15178) );
  MUX21X1 U10981 ( .IN1(\mem1[83][13] ), .IN2(n989), .S(n7587), .Q(n15177) );
  MUX21X1 U10982 ( .IN1(\mem1[83][12] ), .IN2(n967), .S(n7587), .Q(n15176) );
  MUX21X1 U10983 ( .IN1(\mem1[83][11] ), .IN2(n945), .S(n7587), .Q(n15175) );
  MUX21X1 U10984 ( .IN1(\mem1[83][10] ), .IN2(n923), .S(n7587), .Q(n15174) );
  MUX21X1 U10985 ( .IN1(\mem1[83][9] ), .IN2(n901), .S(n7587), .Q(n15173) );
  MUX21X1 U10986 ( .IN1(\mem1[83][8] ), .IN2(n879), .S(n7587), .Q(n15172) );
  AND2X1 U10987 ( .IN1(n7575), .IN2(n7124), .Q(n7587) );
  MUX21X1 U10988 ( .IN1(\mem1[82][15] ), .IN2(n1033), .S(n7588), .Q(n15171) );
  MUX21X1 U10989 ( .IN1(\mem1[82][14] ), .IN2(n1011), .S(n7588), .Q(n15170) );
  MUX21X1 U10990 ( .IN1(\mem1[82][13] ), .IN2(n989), .S(n7588), .Q(n15169) );
  MUX21X1 U10991 ( .IN1(\mem1[82][12] ), .IN2(n967), .S(n7588), .Q(n15168) );
  MUX21X1 U10992 ( .IN1(\mem1[82][11] ), .IN2(n945), .S(n7588), .Q(n15167) );
  MUX21X1 U10993 ( .IN1(\mem1[82][10] ), .IN2(n923), .S(n7588), .Q(n15166) );
  MUX21X1 U10994 ( .IN1(\mem1[82][9] ), .IN2(n901), .S(n7588), .Q(n15165) );
  MUX21X1 U10995 ( .IN1(\mem1[82][8] ), .IN2(n879), .S(n7588), .Q(n15164) );
  AND2X1 U10996 ( .IN1(n7575), .IN2(n7126), .Q(n7588) );
  MUX21X1 U10997 ( .IN1(\mem1[81][15] ), .IN2(n1033), .S(n7589), .Q(n15163) );
  MUX21X1 U10998 ( .IN1(\mem1[81][14] ), .IN2(n1011), .S(n7589), .Q(n15162) );
  MUX21X1 U10999 ( .IN1(\mem1[81][13] ), .IN2(n989), .S(n7589), .Q(n15161) );
  MUX21X1 U11000 ( .IN1(\mem1[81][12] ), .IN2(n967), .S(n7589), .Q(n15160) );
  MUX21X1 U11001 ( .IN1(\mem1[81][11] ), .IN2(n945), .S(n7589), .Q(n15159) );
  MUX21X1 U11002 ( .IN1(\mem1[81][10] ), .IN2(n923), .S(n7589), .Q(n15158) );
  MUX21X1 U11003 ( .IN1(\mem1[81][9] ), .IN2(n901), .S(n7589), .Q(n15157) );
  MUX21X1 U11004 ( .IN1(\mem1[81][8] ), .IN2(n879), .S(n7589), .Q(n15156) );
  AND2X1 U11005 ( .IN1(n7575), .IN2(n7128), .Q(n7589) );
  MUX21X1 U11006 ( .IN1(\mem1[80][15] ), .IN2(n1033), .S(n7590), .Q(n15155) );
  MUX21X1 U11007 ( .IN1(\mem1[80][14] ), .IN2(n1011), .S(n7590), .Q(n15154) );
  MUX21X1 U11008 ( .IN1(\mem1[80][13] ), .IN2(n989), .S(n7590), .Q(n15153) );
  MUX21X1 U11009 ( .IN1(\mem1[80][12] ), .IN2(n967), .S(n7590), .Q(n15152) );
  MUX21X1 U11010 ( .IN1(\mem1[80][11] ), .IN2(n945), .S(n7590), .Q(n15151) );
  MUX21X1 U11011 ( .IN1(\mem1[80][10] ), .IN2(n923), .S(n7590), .Q(n15150) );
  MUX21X1 U11012 ( .IN1(\mem1[80][9] ), .IN2(n901), .S(n7590), .Q(n15149) );
  MUX21X1 U11013 ( .IN1(\mem1[80][8] ), .IN2(n879), .S(n7590), .Q(n15148) );
  AND2X1 U11014 ( .IN1(n7575), .IN2(n7130), .Q(n7590) );
  AND2X1 U11015 ( .IN1(n7420), .IN2(n7312), .Q(n7575) );
  MUX21X1 U11016 ( .IN1(\mem1[79][15] ), .IN2(n1033), .S(n7591), .Q(n15147) );
  MUX21X1 U11017 ( .IN1(\mem1[79][14] ), .IN2(n1011), .S(n7591), .Q(n15146) );
  MUX21X1 U11018 ( .IN1(\mem1[79][13] ), .IN2(n989), .S(n7591), .Q(n15145) );
  MUX21X1 U11019 ( .IN1(\mem1[79][12] ), .IN2(n967), .S(n7591), .Q(n15144) );
  MUX21X1 U11020 ( .IN1(\mem1[79][11] ), .IN2(n945), .S(n7591), .Q(n15143) );
  MUX21X1 U11021 ( .IN1(\mem1[79][10] ), .IN2(n923), .S(n7591), .Q(n15142) );
  MUX21X1 U11022 ( .IN1(\mem1[79][9] ), .IN2(n901), .S(n7591), .Q(n15141) );
  MUX21X1 U11023 ( .IN1(\mem1[79][8] ), .IN2(n879), .S(n7591), .Q(n15140) );
  AND2X1 U11024 ( .IN1(n7592), .IN2(n7099), .Q(n7591) );
  MUX21X1 U11025 ( .IN1(\mem1[78][15] ), .IN2(n1033), .S(n7593), .Q(n15139) );
  MUX21X1 U11026 ( .IN1(\mem1[78][14] ), .IN2(n1011), .S(n7593), .Q(n15138) );
  MUX21X1 U11027 ( .IN1(\mem1[78][13] ), .IN2(n989), .S(n7593), .Q(n15137) );
  MUX21X1 U11028 ( .IN1(\mem1[78][12] ), .IN2(n967), .S(n7593), .Q(n15136) );
  MUX21X1 U11029 ( .IN1(\mem1[78][11] ), .IN2(n945), .S(n7593), .Q(n15135) );
  MUX21X1 U11030 ( .IN1(\mem1[78][10] ), .IN2(n923), .S(n7593), .Q(n15134) );
  MUX21X1 U11031 ( .IN1(\mem1[78][9] ), .IN2(n901), .S(n7593), .Q(n15133) );
  MUX21X1 U11032 ( .IN1(\mem1[78][8] ), .IN2(n879), .S(n7593), .Q(n15132) );
  AND2X1 U11033 ( .IN1(n7592), .IN2(n7102), .Q(n7593) );
  MUX21X1 U11034 ( .IN1(\mem1[77][15] ), .IN2(n1033), .S(n7594), .Q(n15131) );
  MUX21X1 U11035 ( .IN1(\mem1[77][14] ), .IN2(n1011), .S(n7594), .Q(n15130) );
  MUX21X1 U11036 ( .IN1(\mem1[77][13] ), .IN2(n989), .S(n7594), .Q(n15129) );
  MUX21X1 U11037 ( .IN1(\mem1[77][12] ), .IN2(n967), .S(n7594), .Q(n15128) );
  MUX21X1 U11038 ( .IN1(\mem1[77][11] ), .IN2(n945), .S(n7594), .Q(n15127) );
  MUX21X1 U11039 ( .IN1(\mem1[77][10] ), .IN2(n923), .S(n7594), .Q(n15126) );
  MUX21X1 U11040 ( .IN1(\mem1[77][9] ), .IN2(n901), .S(n7594), .Q(n15125) );
  MUX21X1 U11041 ( .IN1(\mem1[77][8] ), .IN2(n879), .S(n7594), .Q(n15124) );
  AND2X1 U11042 ( .IN1(n7592), .IN2(n7104), .Q(n7594) );
  MUX21X1 U11043 ( .IN1(\mem1[76][15] ), .IN2(n1033), .S(n7595), .Q(n15123) );
  MUX21X1 U11044 ( .IN1(\mem1[76][14] ), .IN2(n1011), .S(n7595), .Q(n15122) );
  MUX21X1 U11045 ( .IN1(\mem1[76][13] ), .IN2(n989), .S(n7595), .Q(n15121) );
  MUX21X1 U11046 ( .IN1(\mem1[76][12] ), .IN2(n967), .S(n7595), .Q(n15120) );
  MUX21X1 U11047 ( .IN1(\mem1[76][11] ), .IN2(n945), .S(n7595), .Q(n15119) );
  MUX21X1 U11048 ( .IN1(\mem1[76][10] ), .IN2(n923), .S(n7595), .Q(n15118) );
  MUX21X1 U11049 ( .IN1(\mem1[76][9] ), .IN2(n901), .S(n7595), .Q(n15117) );
  MUX21X1 U11050 ( .IN1(\mem1[76][8] ), .IN2(n879), .S(n7595), .Q(n15116) );
  AND2X1 U11051 ( .IN1(n7592), .IN2(n7106), .Q(n7595) );
  MUX21X1 U11052 ( .IN1(\mem1[75][15] ), .IN2(n1034), .S(n7596), .Q(n15115) );
  MUX21X1 U11053 ( .IN1(\mem1[75][14] ), .IN2(n1012), .S(n7596), .Q(n15114) );
  MUX21X1 U11054 ( .IN1(\mem1[75][13] ), .IN2(n990), .S(n7596), .Q(n15113) );
  MUX21X1 U11055 ( .IN1(\mem1[75][12] ), .IN2(n968), .S(n7596), .Q(n15112) );
  MUX21X1 U11056 ( .IN1(\mem1[75][11] ), .IN2(n946), .S(n7596), .Q(n15111) );
  MUX21X1 U11057 ( .IN1(\mem1[75][10] ), .IN2(n924), .S(n7596), .Q(n15110) );
  MUX21X1 U11058 ( .IN1(\mem1[75][9] ), .IN2(n902), .S(n7596), .Q(n15109) );
  MUX21X1 U11059 ( .IN1(\mem1[75][8] ), .IN2(n880), .S(n7596), .Q(n15108) );
  AND2X1 U11060 ( .IN1(n7592), .IN2(n7108), .Q(n7596) );
  MUX21X1 U11061 ( .IN1(\mem1[74][15] ), .IN2(n1034), .S(n7597), .Q(n15107) );
  MUX21X1 U11062 ( .IN1(\mem1[74][14] ), .IN2(n1012), .S(n7597), .Q(n15106) );
  MUX21X1 U11063 ( .IN1(\mem1[74][13] ), .IN2(n990), .S(n7597), .Q(n15105) );
  MUX21X1 U11064 ( .IN1(\mem1[74][12] ), .IN2(n968), .S(n7597), .Q(n15104) );
  MUX21X1 U11065 ( .IN1(\mem1[74][11] ), .IN2(n946), .S(n7597), .Q(n15103) );
  MUX21X1 U11066 ( .IN1(\mem1[74][10] ), .IN2(n924), .S(n7597), .Q(n15102) );
  MUX21X1 U11067 ( .IN1(\mem1[74][9] ), .IN2(n902), .S(n7597), .Q(n15101) );
  MUX21X1 U11068 ( .IN1(\mem1[74][8] ), .IN2(n880), .S(n7597), .Q(n15100) );
  AND2X1 U11069 ( .IN1(n7592), .IN2(n7110), .Q(n7597) );
  MUX21X1 U11070 ( .IN1(\mem1[73][15] ), .IN2(n1034), .S(n7598), .Q(n15099) );
  MUX21X1 U11071 ( .IN1(\mem1[73][14] ), .IN2(n1012), .S(n7598), .Q(n15098) );
  MUX21X1 U11072 ( .IN1(\mem1[73][13] ), .IN2(n990), .S(n7598), .Q(n15097) );
  MUX21X1 U11073 ( .IN1(\mem1[73][12] ), .IN2(n968), .S(n7598), .Q(n15096) );
  MUX21X1 U11074 ( .IN1(\mem1[73][11] ), .IN2(n946), .S(n7598), .Q(n15095) );
  MUX21X1 U11075 ( .IN1(\mem1[73][10] ), .IN2(n924), .S(n7598), .Q(n15094) );
  MUX21X1 U11076 ( .IN1(\mem1[73][9] ), .IN2(n902), .S(n7598), .Q(n15093) );
  MUX21X1 U11077 ( .IN1(\mem1[73][8] ), .IN2(n880), .S(n7598), .Q(n15092) );
  AND2X1 U11078 ( .IN1(n7592), .IN2(n7112), .Q(n7598) );
  MUX21X1 U11079 ( .IN1(\mem1[72][15] ), .IN2(n1034), .S(n7599), .Q(n15091) );
  MUX21X1 U11080 ( .IN1(\mem1[72][14] ), .IN2(n1012), .S(n7599), .Q(n15090) );
  MUX21X1 U11081 ( .IN1(\mem1[72][13] ), .IN2(n990), .S(n7599), .Q(n15089) );
  MUX21X1 U11082 ( .IN1(\mem1[72][12] ), .IN2(n968), .S(n7599), .Q(n15088) );
  MUX21X1 U11083 ( .IN1(\mem1[72][11] ), .IN2(n946), .S(n7599), .Q(n15087) );
  MUX21X1 U11084 ( .IN1(\mem1[72][10] ), .IN2(n924), .S(n7599), .Q(n15086) );
  MUX21X1 U11085 ( .IN1(\mem1[72][9] ), .IN2(n902), .S(n7599), .Q(n15085) );
  MUX21X1 U11086 ( .IN1(\mem1[72][8] ), .IN2(n880), .S(n7599), .Q(n15084) );
  AND2X1 U11087 ( .IN1(n7592), .IN2(n7114), .Q(n7599) );
  MUX21X1 U11088 ( .IN1(\mem1[71][15] ), .IN2(n1034), .S(n7600), .Q(n15083) );
  MUX21X1 U11089 ( .IN1(\mem1[71][14] ), .IN2(n1012), .S(n7600), .Q(n15082) );
  MUX21X1 U11090 ( .IN1(\mem1[71][13] ), .IN2(n990), .S(n7600), .Q(n15081) );
  MUX21X1 U11091 ( .IN1(\mem1[71][12] ), .IN2(n968), .S(n7600), .Q(n15080) );
  MUX21X1 U11092 ( .IN1(\mem1[71][11] ), .IN2(n946), .S(n7600), .Q(n15079) );
  MUX21X1 U11093 ( .IN1(\mem1[71][10] ), .IN2(n924), .S(n7600), .Q(n15078) );
  MUX21X1 U11094 ( .IN1(\mem1[71][9] ), .IN2(n902), .S(n7600), .Q(n15077) );
  MUX21X1 U11095 ( .IN1(\mem1[71][8] ), .IN2(n880), .S(n7600), .Q(n15076) );
  AND2X1 U11096 ( .IN1(n7592), .IN2(n7116), .Q(n7600) );
  MUX21X1 U11097 ( .IN1(\mem1[70][15] ), .IN2(n1034), .S(n7601), .Q(n15075) );
  MUX21X1 U11098 ( .IN1(\mem1[70][14] ), .IN2(n1012), .S(n7601), .Q(n15074) );
  MUX21X1 U11099 ( .IN1(\mem1[70][13] ), .IN2(n990), .S(n7601), .Q(n15073) );
  MUX21X1 U11100 ( .IN1(\mem1[70][12] ), .IN2(n968), .S(n7601), .Q(n15072) );
  MUX21X1 U11101 ( .IN1(\mem1[70][11] ), .IN2(n946), .S(n7601), .Q(n15071) );
  MUX21X1 U11102 ( .IN1(\mem1[70][10] ), .IN2(n924), .S(n7601), .Q(n15070) );
  MUX21X1 U11103 ( .IN1(\mem1[70][9] ), .IN2(n902), .S(n7601), .Q(n15069) );
  MUX21X1 U11104 ( .IN1(\mem1[70][8] ), .IN2(n880), .S(n7601), .Q(n15068) );
  AND2X1 U11105 ( .IN1(n7592), .IN2(n7118), .Q(n7601) );
  MUX21X1 U11106 ( .IN1(\mem1[69][15] ), .IN2(n1034), .S(n7602), .Q(n15067) );
  MUX21X1 U11107 ( .IN1(\mem1[69][14] ), .IN2(n1012), .S(n7602), .Q(n15066) );
  MUX21X1 U11108 ( .IN1(\mem1[69][13] ), .IN2(n990), .S(n7602), .Q(n15065) );
  MUX21X1 U11109 ( .IN1(\mem1[69][12] ), .IN2(n968), .S(n7602), .Q(n15064) );
  MUX21X1 U11110 ( .IN1(\mem1[69][11] ), .IN2(n946), .S(n7602), .Q(n15063) );
  MUX21X1 U11111 ( .IN1(\mem1[69][10] ), .IN2(n924), .S(n7602), .Q(n15062) );
  MUX21X1 U11112 ( .IN1(\mem1[69][9] ), .IN2(n902), .S(n7602), .Q(n15061) );
  MUX21X1 U11113 ( .IN1(\mem1[69][8] ), .IN2(n880), .S(n7602), .Q(n15060) );
  AND2X1 U11114 ( .IN1(n7592), .IN2(n7120), .Q(n7602) );
  MUX21X1 U11115 ( .IN1(\mem1[68][15] ), .IN2(n1034), .S(n7603), .Q(n15059) );
  MUX21X1 U11116 ( .IN1(\mem1[68][14] ), .IN2(n1012), .S(n7603), .Q(n15058) );
  MUX21X1 U11117 ( .IN1(\mem1[68][13] ), .IN2(n990), .S(n7603), .Q(n15057) );
  MUX21X1 U11118 ( .IN1(\mem1[68][12] ), .IN2(n968), .S(n7603), .Q(n15056) );
  MUX21X1 U11119 ( .IN1(\mem1[68][11] ), .IN2(n946), .S(n7603), .Q(n15055) );
  MUX21X1 U11120 ( .IN1(\mem1[68][10] ), .IN2(n924), .S(n7603), .Q(n15054) );
  MUX21X1 U11121 ( .IN1(\mem1[68][9] ), .IN2(n902), .S(n7603), .Q(n15053) );
  MUX21X1 U11122 ( .IN1(\mem1[68][8] ), .IN2(n880), .S(n7603), .Q(n15052) );
  AND2X1 U11123 ( .IN1(n7592), .IN2(n7122), .Q(n7603) );
  MUX21X1 U11124 ( .IN1(\mem1[67][15] ), .IN2(n1034), .S(n7604), .Q(n15051) );
  MUX21X1 U11125 ( .IN1(\mem1[67][14] ), .IN2(n1012), .S(n7604), .Q(n15050) );
  MUX21X1 U11126 ( .IN1(\mem1[67][13] ), .IN2(n990), .S(n7604), .Q(n15049) );
  MUX21X1 U11127 ( .IN1(\mem1[67][12] ), .IN2(n968), .S(n7604), .Q(n15048) );
  MUX21X1 U11128 ( .IN1(\mem1[67][11] ), .IN2(n946), .S(n7604), .Q(n15047) );
  MUX21X1 U11129 ( .IN1(\mem1[67][10] ), .IN2(n924), .S(n7604), .Q(n15046) );
  MUX21X1 U11130 ( .IN1(\mem1[67][9] ), .IN2(n902), .S(n7604), .Q(n15045) );
  MUX21X1 U11131 ( .IN1(\mem1[67][8] ), .IN2(n880), .S(n7604), .Q(n15044) );
  AND2X1 U11132 ( .IN1(n7592), .IN2(n7124), .Q(n7604) );
  MUX21X1 U11133 ( .IN1(\mem1[66][15] ), .IN2(n1034), .S(n7605), .Q(n15043) );
  MUX21X1 U11134 ( .IN1(\mem1[66][14] ), .IN2(n1012), .S(n7605), .Q(n15042) );
  MUX21X1 U11135 ( .IN1(\mem1[66][13] ), .IN2(n990), .S(n7605), .Q(n15041) );
  MUX21X1 U11136 ( .IN1(\mem1[66][12] ), .IN2(n968), .S(n7605), .Q(n15040) );
  MUX21X1 U11137 ( .IN1(\mem1[66][11] ), .IN2(n946), .S(n7605), .Q(n15039) );
  MUX21X1 U11138 ( .IN1(\mem1[66][10] ), .IN2(n924), .S(n7605), .Q(n15038) );
  MUX21X1 U11139 ( .IN1(\mem1[66][9] ), .IN2(n902), .S(n7605), .Q(n15037) );
  MUX21X1 U11140 ( .IN1(\mem1[66][8] ), .IN2(n880), .S(n7605), .Q(n15036) );
  AND2X1 U11141 ( .IN1(n7592), .IN2(n7126), .Q(n7605) );
  MUX21X1 U11142 ( .IN1(\mem1[65][15] ), .IN2(n1034), .S(n7606), .Q(n15035) );
  MUX21X1 U11143 ( .IN1(\mem1[65][14] ), .IN2(n1012), .S(n7606), .Q(n15034) );
  MUX21X1 U11144 ( .IN1(\mem1[65][13] ), .IN2(n990), .S(n7606), .Q(n15033) );
  MUX21X1 U11145 ( .IN1(\mem1[65][12] ), .IN2(n968), .S(n7606), .Q(n15032) );
  MUX21X1 U11146 ( .IN1(\mem1[65][11] ), .IN2(n946), .S(n7606), .Q(n15031) );
  MUX21X1 U11147 ( .IN1(\mem1[65][10] ), .IN2(n924), .S(n7606), .Q(n15030) );
  MUX21X1 U11148 ( .IN1(\mem1[65][9] ), .IN2(n902), .S(n7606), .Q(n15029) );
  MUX21X1 U11149 ( .IN1(\mem1[65][8] ), .IN2(n880), .S(n7606), .Q(n15028) );
  AND2X1 U11150 ( .IN1(n7592), .IN2(n7128), .Q(n7606) );
  MUX21X1 U11151 ( .IN1(\mem1[64][15] ), .IN2(n1034), .S(n7607), .Q(n15027) );
  MUX21X1 U11152 ( .IN1(\mem1[64][14] ), .IN2(n1012), .S(n7607), .Q(n15026) );
  MUX21X1 U11153 ( .IN1(\mem1[64][13] ), .IN2(n990), .S(n7607), .Q(n15025) );
  MUX21X1 U11154 ( .IN1(\mem1[64][12] ), .IN2(n968), .S(n7607), .Q(n15024) );
  MUX21X1 U11155 ( .IN1(\mem1[64][11] ), .IN2(n946), .S(n7607), .Q(n15023) );
  MUX21X1 U11156 ( .IN1(\mem1[64][10] ), .IN2(n924), .S(n7607), .Q(n15022) );
  MUX21X1 U11157 ( .IN1(\mem1[64][9] ), .IN2(n902), .S(n7607), .Q(n15021) );
  MUX21X1 U11158 ( .IN1(\mem1[64][8] ), .IN2(n880), .S(n7607), .Q(n15020) );
  AND2X1 U11159 ( .IN1(n7592), .IN2(n7130), .Q(n7607) );
  AND2X1 U11160 ( .IN1(n7420), .IN2(n7330), .Q(n7592) );
  MUX21X1 U11161 ( .IN1(\mem1[63][15] ), .IN2(n1035), .S(n7608), .Q(n15019) );
  MUX21X1 U11162 ( .IN1(\mem1[63][14] ), .IN2(n1013), .S(n7608), .Q(n15018) );
  MUX21X1 U11163 ( .IN1(\mem1[63][13] ), .IN2(n991), .S(n7608), .Q(n15017) );
  MUX21X1 U11164 ( .IN1(\mem1[63][12] ), .IN2(n969), .S(n7608), .Q(n15016) );
  MUX21X1 U11165 ( .IN1(\mem1[63][11] ), .IN2(n947), .S(n7608), .Q(n15015) );
  MUX21X1 U11166 ( .IN1(\mem1[63][10] ), .IN2(n925), .S(n7608), .Q(n15014) );
  MUX21X1 U11167 ( .IN1(\mem1[63][9] ), .IN2(n903), .S(n7608), .Q(n15013) );
  MUX21X1 U11168 ( .IN1(\mem1[63][8] ), .IN2(n881), .S(n7608), .Q(n15012) );
  AND2X1 U11169 ( .IN1(n7609), .IN2(n7099), .Q(n7608) );
  MUX21X1 U11170 ( .IN1(\mem1[62][15] ), .IN2(n1035), .S(n7610), .Q(n15011) );
  MUX21X1 U11171 ( .IN1(\mem1[62][14] ), .IN2(n1013), .S(n7610), .Q(n15010) );
  MUX21X1 U11172 ( .IN1(\mem1[62][13] ), .IN2(n991), .S(n7610), .Q(n15009) );
  MUX21X1 U11173 ( .IN1(\mem1[62][12] ), .IN2(n969), .S(n7610), .Q(n15008) );
  MUX21X1 U11174 ( .IN1(\mem1[62][11] ), .IN2(n947), .S(n7610), .Q(n15007) );
  MUX21X1 U11175 ( .IN1(\mem1[62][10] ), .IN2(n925), .S(n7610), .Q(n15006) );
  MUX21X1 U11176 ( .IN1(\mem1[62][9] ), .IN2(n903), .S(n7610), .Q(n15005) );
  MUX21X1 U11177 ( .IN1(\mem1[62][8] ), .IN2(n881), .S(n7610), .Q(n15004) );
  AND2X1 U11178 ( .IN1(n7609), .IN2(n7102), .Q(n7610) );
  MUX21X1 U11179 ( .IN1(\mem1[61][15] ), .IN2(n1035), .S(n7611), .Q(n15003) );
  MUX21X1 U11180 ( .IN1(\mem1[61][14] ), .IN2(n1013), .S(n7611), .Q(n15002) );
  MUX21X1 U11181 ( .IN1(\mem1[61][13] ), .IN2(n991), .S(n7611), .Q(n15001) );
  MUX21X1 U11182 ( .IN1(\mem1[61][12] ), .IN2(n969), .S(n7611), .Q(n15000) );
  MUX21X1 U11183 ( .IN1(\mem1[61][11] ), .IN2(n947), .S(n7611), .Q(n14999) );
  MUX21X1 U11184 ( .IN1(\mem1[61][10] ), .IN2(n925), .S(n7611), .Q(n14998) );
  MUX21X1 U11185 ( .IN1(\mem1[61][9] ), .IN2(n903), .S(n7611), .Q(n14997) );
  MUX21X1 U11186 ( .IN1(\mem1[61][8] ), .IN2(n881), .S(n7611), .Q(n14996) );
  AND2X1 U11187 ( .IN1(n7609), .IN2(n7104), .Q(n7611) );
  MUX21X1 U11188 ( .IN1(\mem1[60][15] ), .IN2(n1035), .S(n7612), .Q(n14995) );
  MUX21X1 U11189 ( .IN1(\mem1[60][14] ), .IN2(n1013), .S(n7612), .Q(n14994) );
  MUX21X1 U11190 ( .IN1(\mem1[60][13] ), .IN2(n991), .S(n7612), .Q(n14993) );
  MUX21X1 U11191 ( .IN1(\mem1[60][12] ), .IN2(n969), .S(n7612), .Q(n14992) );
  MUX21X1 U11192 ( .IN1(\mem1[60][11] ), .IN2(n947), .S(n7612), .Q(n14991) );
  MUX21X1 U11193 ( .IN1(\mem1[60][10] ), .IN2(n925), .S(n7612), .Q(n14990) );
  MUX21X1 U11194 ( .IN1(\mem1[60][9] ), .IN2(n903), .S(n7612), .Q(n14989) );
  MUX21X1 U11195 ( .IN1(\mem1[60][8] ), .IN2(n881), .S(n7612), .Q(n14988) );
  AND2X1 U11196 ( .IN1(n7609), .IN2(n7106), .Q(n7612) );
  MUX21X1 U11197 ( .IN1(\mem1[59][15] ), .IN2(n1035), .S(n7613), .Q(n14987) );
  MUX21X1 U11198 ( .IN1(\mem1[59][14] ), .IN2(n1013), .S(n7613), .Q(n14986) );
  MUX21X1 U11199 ( .IN1(\mem1[59][13] ), .IN2(n991), .S(n7613), .Q(n14985) );
  MUX21X1 U11200 ( .IN1(\mem1[59][12] ), .IN2(n969), .S(n7613), .Q(n14984) );
  MUX21X1 U11201 ( .IN1(\mem1[59][11] ), .IN2(n947), .S(n7613), .Q(n14983) );
  MUX21X1 U11202 ( .IN1(\mem1[59][10] ), .IN2(n925), .S(n7613), .Q(n14982) );
  MUX21X1 U11203 ( .IN1(\mem1[59][9] ), .IN2(n903), .S(n7613), .Q(n14981) );
  MUX21X1 U11204 ( .IN1(\mem1[59][8] ), .IN2(n881), .S(n7613), .Q(n14980) );
  AND2X1 U11205 ( .IN1(n7609), .IN2(n7108), .Q(n7613) );
  MUX21X1 U11206 ( .IN1(\mem1[58][15] ), .IN2(n1035), .S(n7614), .Q(n14979) );
  MUX21X1 U11207 ( .IN1(\mem1[58][14] ), .IN2(n1013), .S(n7614), .Q(n14978) );
  MUX21X1 U11208 ( .IN1(\mem1[58][13] ), .IN2(n991), .S(n7614), .Q(n14977) );
  MUX21X1 U11209 ( .IN1(\mem1[58][12] ), .IN2(n969), .S(n7614), .Q(n14976) );
  MUX21X1 U11210 ( .IN1(\mem1[58][11] ), .IN2(n947), .S(n7614), .Q(n14975) );
  MUX21X1 U11211 ( .IN1(\mem1[58][10] ), .IN2(n925), .S(n7614), .Q(n14974) );
  MUX21X1 U11212 ( .IN1(\mem1[58][9] ), .IN2(n903), .S(n7614), .Q(n14973) );
  MUX21X1 U11213 ( .IN1(\mem1[58][8] ), .IN2(n881), .S(n7614), .Q(n14972) );
  AND2X1 U11214 ( .IN1(n7609), .IN2(n7110), .Q(n7614) );
  MUX21X1 U11215 ( .IN1(\mem1[57][15] ), .IN2(n1035), .S(n7615), .Q(n14971) );
  MUX21X1 U11216 ( .IN1(\mem1[57][14] ), .IN2(n1013), .S(n7615), .Q(n14970) );
  MUX21X1 U11217 ( .IN1(\mem1[57][13] ), .IN2(n991), .S(n7615), .Q(n14969) );
  MUX21X1 U11218 ( .IN1(\mem1[57][12] ), .IN2(n969), .S(n7615), .Q(n14968) );
  MUX21X1 U11219 ( .IN1(\mem1[57][11] ), .IN2(n947), .S(n7615), .Q(n14967) );
  MUX21X1 U11220 ( .IN1(\mem1[57][10] ), .IN2(n925), .S(n7615), .Q(n14966) );
  MUX21X1 U11221 ( .IN1(\mem1[57][9] ), .IN2(n903), .S(n7615), .Q(n14965) );
  MUX21X1 U11222 ( .IN1(\mem1[57][8] ), .IN2(n881), .S(n7615), .Q(n14964) );
  AND2X1 U11223 ( .IN1(n7609), .IN2(n7112), .Q(n7615) );
  MUX21X1 U11224 ( .IN1(\mem1[56][15] ), .IN2(n1035), .S(n7616), .Q(n14963) );
  MUX21X1 U11225 ( .IN1(\mem1[56][14] ), .IN2(n1013), .S(n7616), .Q(n14962) );
  MUX21X1 U11226 ( .IN1(\mem1[56][13] ), .IN2(n991), .S(n7616), .Q(n14961) );
  MUX21X1 U11227 ( .IN1(\mem1[56][12] ), .IN2(n969), .S(n7616), .Q(n14960) );
  MUX21X1 U11228 ( .IN1(\mem1[56][11] ), .IN2(n947), .S(n7616), .Q(n14959) );
  MUX21X1 U11229 ( .IN1(\mem1[56][10] ), .IN2(n925), .S(n7616), .Q(n14958) );
  MUX21X1 U11230 ( .IN1(\mem1[56][9] ), .IN2(n903), .S(n7616), .Q(n14957) );
  MUX21X1 U11231 ( .IN1(\mem1[56][8] ), .IN2(n881), .S(n7616), .Q(n14956) );
  AND2X1 U11232 ( .IN1(n7609), .IN2(n7114), .Q(n7616) );
  MUX21X1 U11233 ( .IN1(\mem1[55][15] ), .IN2(n1035), .S(n7617), .Q(n14955) );
  MUX21X1 U11234 ( .IN1(\mem1[55][14] ), .IN2(n1013), .S(n7617), .Q(n14954) );
  MUX21X1 U11235 ( .IN1(\mem1[55][13] ), .IN2(n991), .S(n7617), .Q(n14953) );
  MUX21X1 U11236 ( .IN1(\mem1[55][12] ), .IN2(n969), .S(n7617), .Q(n14952) );
  MUX21X1 U11237 ( .IN1(\mem1[55][11] ), .IN2(n947), .S(n7617), .Q(n14951) );
  MUX21X1 U11238 ( .IN1(\mem1[55][10] ), .IN2(n925), .S(n7617), .Q(n14950) );
  MUX21X1 U11239 ( .IN1(\mem1[55][9] ), .IN2(n903), .S(n7617), .Q(n14949) );
  MUX21X1 U11240 ( .IN1(\mem1[55][8] ), .IN2(n881), .S(n7617), .Q(n14948) );
  AND2X1 U11241 ( .IN1(n7609), .IN2(n7116), .Q(n7617) );
  MUX21X1 U11242 ( .IN1(\mem1[54][15] ), .IN2(n1035), .S(n7618), .Q(n14947) );
  MUX21X1 U11243 ( .IN1(\mem1[54][14] ), .IN2(n1013), .S(n7618), .Q(n14946) );
  MUX21X1 U11244 ( .IN1(\mem1[54][13] ), .IN2(n991), .S(n7618), .Q(n14945) );
  MUX21X1 U11245 ( .IN1(\mem1[54][12] ), .IN2(n969), .S(n7618), .Q(n14944) );
  MUX21X1 U11246 ( .IN1(\mem1[54][11] ), .IN2(n947), .S(n7618), .Q(n14943) );
  MUX21X1 U11247 ( .IN1(\mem1[54][10] ), .IN2(n925), .S(n7618), .Q(n14942) );
  MUX21X1 U11248 ( .IN1(\mem1[54][9] ), .IN2(n903), .S(n7618), .Q(n14941) );
  MUX21X1 U11249 ( .IN1(\mem1[54][8] ), .IN2(n881), .S(n7618), .Q(n14940) );
  AND2X1 U11250 ( .IN1(n7609), .IN2(n7118), .Q(n7618) );
  MUX21X1 U11251 ( .IN1(\mem1[53][15] ), .IN2(n1035), .S(n7619), .Q(n14939) );
  MUX21X1 U11252 ( .IN1(\mem1[53][14] ), .IN2(n1013), .S(n7619), .Q(n14938) );
  MUX21X1 U11253 ( .IN1(\mem1[53][13] ), .IN2(n991), .S(n7619), .Q(n14937) );
  MUX21X1 U11254 ( .IN1(\mem1[53][12] ), .IN2(n969), .S(n7619), .Q(n14936) );
  MUX21X1 U11255 ( .IN1(\mem1[53][11] ), .IN2(n947), .S(n7619), .Q(n14935) );
  MUX21X1 U11256 ( .IN1(\mem1[53][10] ), .IN2(n925), .S(n7619), .Q(n14934) );
  MUX21X1 U11257 ( .IN1(\mem1[53][9] ), .IN2(n903), .S(n7619), .Q(n14933) );
  MUX21X1 U11258 ( .IN1(\mem1[53][8] ), .IN2(n881), .S(n7619), .Q(n14932) );
  AND2X1 U11259 ( .IN1(n7609), .IN2(n7120), .Q(n7619) );
  MUX21X1 U11260 ( .IN1(\mem1[52][15] ), .IN2(n1035), .S(n7620), .Q(n14931) );
  MUX21X1 U11261 ( .IN1(\mem1[52][14] ), .IN2(n1013), .S(n7620), .Q(n14930) );
  MUX21X1 U11262 ( .IN1(\mem1[52][13] ), .IN2(n991), .S(n7620), .Q(n14929) );
  MUX21X1 U11263 ( .IN1(\mem1[52][12] ), .IN2(n969), .S(n7620), .Q(n14928) );
  MUX21X1 U11264 ( .IN1(\mem1[52][11] ), .IN2(n947), .S(n7620), .Q(n14927) );
  MUX21X1 U11265 ( .IN1(\mem1[52][10] ), .IN2(n925), .S(n7620), .Q(n14926) );
  MUX21X1 U11266 ( .IN1(\mem1[52][9] ), .IN2(n903), .S(n7620), .Q(n14925) );
  MUX21X1 U11267 ( .IN1(\mem1[52][8] ), .IN2(n881), .S(n7620), .Q(n14924) );
  AND2X1 U11268 ( .IN1(n7609), .IN2(n7122), .Q(n7620) );
  MUX21X1 U11269 ( .IN1(\mem1[51][15] ), .IN2(n1036), .S(n7621), .Q(n14923) );
  MUX21X1 U11270 ( .IN1(\mem1[51][14] ), .IN2(n1014), .S(n7621), .Q(n14922) );
  MUX21X1 U11271 ( .IN1(\mem1[51][13] ), .IN2(n992), .S(n7621), .Q(n14921) );
  MUX21X1 U11272 ( .IN1(\mem1[51][12] ), .IN2(n970), .S(n7621), .Q(n14920) );
  MUX21X1 U11273 ( .IN1(\mem1[51][11] ), .IN2(n948), .S(n7621), .Q(n14919) );
  MUX21X1 U11274 ( .IN1(\mem1[51][10] ), .IN2(n926), .S(n7621), .Q(n14918) );
  MUX21X1 U11275 ( .IN1(\mem1[51][9] ), .IN2(n904), .S(n7621), .Q(n14917) );
  MUX21X1 U11276 ( .IN1(\mem1[51][8] ), .IN2(n882), .S(n7621), .Q(n14916) );
  AND2X1 U11277 ( .IN1(n7609), .IN2(n7124), .Q(n7621) );
  MUX21X1 U11278 ( .IN1(\mem1[50][15] ), .IN2(n1036), .S(n7622), .Q(n14915) );
  MUX21X1 U11279 ( .IN1(\mem1[50][14] ), .IN2(n1014), .S(n7622), .Q(n14914) );
  MUX21X1 U11280 ( .IN1(\mem1[50][13] ), .IN2(n992), .S(n7622), .Q(n14913) );
  MUX21X1 U11281 ( .IN1(\mem1[50][12] ), .IN2(n970), .S(n7622), .Q(n14912) );
  MUX21X1 U11282 ( .IN1(\mem1[50][11] ), .IN2(n948), .S(n7622), .Q(n14911) );
  MUX21X1 U11283 ( .IN1(\mem1[50][10] ), .IN2(n926), .S(n7622), .Q(n14910) );
  MUX21X1 U11284 ( .IN1(\mem1[50][9] ), .IN2(n904), .S(n7622), .Q(n14909) );
  MUX21X1 U11285 ( .IN1(\mem1[50][8] ), .IN2(n882), .S(n7622), .Q(n14908) );
  AND2X1 U11286 ( .IN1(n7609), .IN2(n7126), .Q(n7622) );
  MUX21X1 U11287 ( .IN1(\mem1[49][15] ), .IN2(n1036), .S(n7623), .Q(n14907) );
  MUX21X1 U11288 ( .IN1(\mem1[49][14] ), .IN2(n1014), .S(n7623), .Q(n14906) );
  MUX21X1 U11289 ( .IN1(\mem1[49][13] ), .IN2(n992), .S(n7623), .Q(n14905) );
  MUX21X1 U11290 ( .IN1(\mem1[49][12] ), .IN2(n970), .S(n7623), .Q(n14904) );
  MUX21X1 U11291 ( .IN1(\mem1[49][11] ), .IN2(n948), .S(n7623), .Q(n14903) );
  MUX21X1 U11292 ( .IN1(\mem1[49][10] ), .IN2(n926), .S(n7623), .Q(n14902) );
  MUX21X1 U11293 ( .IN1(\mem1[49][9] ), .IN2(n904), .S(n7623), .Q(n14901) );
  MUX21X1 U11294 ( .IN1(\mem1[49][8] ), .IN2(n882), .S(n7623), .Q(n14900) );
  AND2X1 U11295 ( .IN1(n7609), .IN2(n7128), .Q(n7623) );
  MUX21X1 U11296 ( .IN1(\mem1[48][15] ), .IN2(n1036), .S(n7624), .Q(n14899) );
  MUX21X1 U11297 ( .IN1(\mem1[48][14] ), .IN2(n1014), .S(n7624), .Q(n14898) );
  MUX21X1 U11298 ( .IN1(\mem1[48][13] ), .IN2(n992), .S(n7624), .Q(n14897) );
  MUX21X1 U11299 ( .IN1(\mem1[48][12] ), .IN2(n970), .S(n7624), .Q(n14896) );
  MUX21X1 U11300 ( .IN1(\mem1[48][11] ), .IN2(n948), .S(n7624), .Q(n14895) );
  MUX21X1 U11301 ( .IN1(\mem1[48][10] ), .IN2(n926), .S(n7624), .Q(n14894) );
  MUX21X1 U11302 ( .IN1(\mem1[48][9] ), .IN2(n904), .S(n7624), .Q(n14893) );
  MUX21X1 U11303 ( .IN1(\mem1[48][8] ), .IN2(n882), .S(n7624), .Q(n14892) );
  AND2X1 U11304 ( .IN1(n7609), .IN2(n7130), .Q(n7624) );
  AND2X1 U11305 ( .IN1(n7420), .IN2(n7348), .Q(n7609) );
  MUX21X1 U11306 ( .IN1(\mem1[47][15] ), .IN2(n1036), .S(n7625), .Q(n14891) );
  MUX21X1 U11307 ( .IN1(\mem1[47][14] ), .IN2(n1014), .S(n7625), .Q(n14890) );
  MUX21X1 U11308 ( .IN1(\mem1[47][13] ), .IN2(n992), .S(n7625), .Q(n14889) );
  MUX21X1 U11309 ( .IN1(\mem1[47][12] ), .IN2(n970), .S(n7625), .Q(n14888) );
  MUX21X1 U11310 ( .IN1(\mem1[47][11] ), .IN2(n948), .S(n7625), .Q(n14887) );
  MUX21X1 U11311 ( .IN1(\mem1[47][10] ), .IN2(n926), .S(n7625), .Q(n14886) );
  MUX21X1 U11312 ( .IN1(\mem1[47][9] ), .IN2(n904), .S(n7625), .Q(n14885) );
  MUX21X1 U11313 ( .IN1(\mem1[47][8] ), .IN2(n882), .S(n7625), .Q(n14884) );
  AND2X1 U11314 ( .IN1(n7626), .IN2(n7099), .Q(n7625) );
  MUX21X1 U11315 ( .IN1(\mem1[46][15] ), .IN2(n1036), .S(n7627), .Q(n14883) );
  MUX21X1 U11316 ( .IN1(\mem1[46][14] ), .IN2(n1014), .S(n7627), .Q(n14882) );
  MUX21X1 U11317 ( .IN1(\mem1[46][13] ), .IN2(n992), .S(n7627), .Q(n14881) );
  MUX21X1 U11318 ( .IN1(\mem1[46][12] ), .IN2(n970), .S(n7627), .Q(n14880) );
  MUX21X1 U11319 ( .IN1(\mem1[46][11] ), .IN2(n948), .S(n7627), .Q(n14879) );
  MUX21X1 U11320 ( .IN1(\mem1[46][10] ), .IN2(n926), .S(n7627), .Q(n14878) );
  MUX21X1 U11321 ( .IN1(\mem1[46][9] ), .IN2(n904), .S(n7627), .Q(n14877) );
  MUX21X1 U11322 ( .IN1(\mem1[46][8] ), .IN2(n882), .S(n7627), .Q(n14876) );
  AND2X1 U11323 ( .IN1(n7626), .IN2(n7102), .Q(n7627) );
  MUX21X1 U11324 ( .IN1(\mem1[45][15] ), .IN2(n1036), .S(n7628), .Q(n14875) );
  MUX21X1 U11325 ( .IN1(\mem1[45][14] ), .IN2(n1014), .S(n7628), .Q(n14874) );
  MUX21X1 U11326 ( .IN1(\mem1[45][13] ), .IN2(n992), .S(n7628), .Q(n14873) );
  MUX21X1 U11327 ( .IN1(\mem1[45][12] ), .IN2(n970), .S(n7628), .Q(n14872) );
  MUX21X1 U11328 ( .IN1(\mem1[45][11] ), .IN2(n948), .S(n7628), .Q(n14871) );
  MUX21X1 U11329 ( .IN1(\mem1[45][10] ), .IN2(n926), .S(n7628), .Q(n14870) );
  MUX21X1 U11330 ( .IN1(\mem1[45][9] ), .IN2(n904), .S(n7628), .Q(n14869) );
  MUX21X1 U11331 ( .IN1(\mem1[45][8] ), .IN2(n882), .S(n7628), .Q(n14868) );
  AND2X1 U11332 ( .IN1(n7626), .IN2(n7104), .Q(n7628) );
  MUX21X1 U11333 ( .IN1(\mem1[44][15] ), .IN2(n1036), .S(n7629), .Q(n14867) );
  MUX21X1 U11334 ( .IN1(\mem1[44][14] ), .IN2(n1014), .S(n7629), .Q(n14866) );
  MUX21X1 U11335 ( .IN1(\mem1[44][13] ), .IN2(n992), .S(n7629), .Q(n14865) );
  MUX21X1 U11336 ( .IN1(\mem1[44][12] ), .IN2(n970), .S(n7629), .Q(n14864) );
  MUX21X1 U11337 ( .IN1(\mem1[44][11] ), .IN2(n948), .S(n7629), .Q(n14863) );
  MUX21X1 U11338 ( .IN1(\mem1[44][10] ), .IN2(n926), .S(n7629), .Q(n14862) );
  MUX21X1 U11339 ( .IN1(\mem1[44][9] ), .IN2(n904), .S(n7629), .Q(n14861) );
  MUX21X1 U11340 ( .IN1(\mem1[44][8] ), .IN2(n882), .S(n7629), .Q(n14860) );
  AND2X1 U11341 ( .IN1(n7626), .IN2(n7106), .Q(n7629) );
  MUX21X1 U11342 ( .IN1(\mem1[43][15] ), .IN2(n1036), .S(n7630), .Q(n14859) );
  MUX21X1 U11343 ( .IN1(\mem1[43][14] ), .IN2(n1014), .S(n7630), .Q(n14858) );
  MUX21X1 U11344 ( .IN1(\mem1[43][13] ), .IN2(n992), .S(n7630), .Q(n14857) );
  MUX21X1 U11345 ( .IN1(\mem1[43][12] ), .IN2(n970), .S(n7630), .Q(n14856) );
  MUX21X1 U11346 ( .IN1(\mem1[43][11] ), .IN2(n948), .S(n7630), .Q(n14855) );
  MUX21X1 U11347 ( .IN1(\mem1[43][10] ), .IN2(n926), .S(n7630), .Q(n14854) );
  MUX21X1 U11348 ( .IN1(\mem1[43][9] ), .IN2(n904), .S(n7630), .Q(n14853) );
  MUX21X1 U11349 ( .IN1(\mem1[43][8] ), .IN2(n882), .S(n7630), .Q(n14852) );
  AND2X1 U11350 ( .IN1(n7626), .IN2(n7108), .Q(n7630) );
  MUX21X1 U11351 ( .IN1(\mem1[42][15] ), .IN2(n1036), .S(n7631), .Q(n14851) );
  MUX21X1 U11352 ( .IN1(\mem1[42][14] ), .IN2(n1014), .S(n7631), .Q(n14850) );
  MUX21X1 U11353 ( .IN1(\mem1[42][13] ), .IN2(n992), .S(n7631), .Q(n14849) );
  MUX21X1 U11354 ( .IN1(\mem1[42][12] ), .IN2(n970), .S(n7631), .Q(n14848) );
  MUX21X1 U11355 ( .IN1(\mem1[42][11] ), .IN2(n948), .S(n7631), .Q(n14847) );
  MUX21X1 U11356 ( .IN1(\mem1[42][10] ), .IN2(n926), .S(n7631), .Q(n14846) );
  MUX21X1 U11357 ( .IN1(\mem1[42][9] ), .IN2(n904), .S(n7631), .Q(n14845) );
  MUX21X1 U11358 ( .IN1(\mem1[42][8] ), .IN2(n882), .S(n7631), .Q(n14844) );
  AND2X1 U11359 ( .IN1(n7626), .IN2(n7110), .Q(n7631) );
  MUX21X1 U11360 ( .IN1(\mem1[41][15] ), .IN2(n1036), .S(n7632), .Q(n14843) );
  MUX21X1 U11361 ( .IN1(\mem1[41][14] ), .IN2(n1014), .S(n7632), .Q(n14842) );
  MUX21X1 U11362 ( .IN1(\mem1[41][13] ), .IN2(n992), .S(n7632), .Q(n14841) );
  MUX21X1 U11363 ( .IN1(\mem1[41][12] ), .IN2(n970), .S(n7632), .Q(n14840) );
  MUX21X1 U11364 ( .IN1(\mem1[41][11] ), .IN2(n948), .S(n7632), .Q(n14839) );
  MUX21X1 U11365 ( .IN1(\mem1[41][10] ), .IN2(n926), .S(n7632), .Q(n14838) );
  MUX21X1 U11366 ( .IN1(\mem1[41][9] ), .IN2(n904), .S(n7632), .Q(n14837) );
  MUX21X1 U11367 ( .IN1(\mem1[41][8] ), .IN2(n882), .S(n7632), .Q(n14836) );
  AND2X1 U11368 ( .IN1(n7626), .IN2(n7112), .Q(n7632) );
  MUX21X1 U11369 ( .IN1(\mem1[40][15] ), .IN2(n1036), .S(n7633), .Q(n14835) );
  MUX21X1 U11370 ( .IN1(\mem1[40][14] ), .IN2(n1014), .S(n7633), .Q(n14834) );
  MUX21X1 U11371 ( .IN1(\mem1[40][13] ), .IN2(n992), .S(n7633), .Q(n14833) );
  MUX21X1 U11372 ( .IN1(\mem1[40][12] ), .IN2(n970), .S(n7633), .Q(n14832) );
  MUX21X1 U11373 ( .IN1(\mem1[40][11] ), .IN2(n948), .S(n7633), .Q(n14831) );
  MUX21X1 U11374 ( .IN1(\mem1[40][10] ), .IN2(n926), .S(n7633), .Q(n14830) );
  MUX21X1 U11375 ( .IN1(\mem1[40][9] ), .IN2(n904), .S(n7633), .Q(n14829) );
  MUX21X1 U11376 ( .IN1(\mem1[40][8] ), .IN2(n882), .S(n7633), .Q(n14828) );
  AND2X1 U11377 ( .IN1(n7626), .IN2(n7114), .Q(n7633) );
  MUX21X1 U11378 ( .IN1(\mem1[39][15] ), .IN2(n1037), .S(n7634), .Q(n14827) );
  MUX21X1 U11379 ( .IN1(\mem1[39][14] ), .IN2(n1015), .S(n7634), .Q(n14826) );
  MUX21X1 U11380 ( .IN1(\mem1[39][13] ), .IN2(n993), .S(n7634), .Q(n14825) );
  MUX21X1 U11381 ( .IN1(\mem1[39][12] ), .IN2(n971), .S(n7634), .Q(n14824) );
  MUX21X1 U11382 ( .IN1(\mem1[39][11] ), .IN2(n949), .S(n7634), .Q(n14823) );
  MUX21X1 U11383 ( .IN1(\mem1[39][10] ), .IN2(n927), .S(n7634), .Q(n14822) );
  MUX21X1 U11384 ( .IN1(\mem1[39][9] ), .IN2(n905), .S(n7634), .Q(n14821) );
  MUX21X1 U11385 ( .IN1(\mem1[39][8] ), .IN2(n883), .S(n7634), .Q(n14820) );
  AND2X1 U11386 ( .IN1(n7626), .IN2(n7116), .Q(n7634) );
  MUX21X1 U11387 ( .IN1(\mem1[38][15] ), .IN2(n1037), .S(n7635), .Q(n14819) );
  MUX21X1 U11388 ( .IN1(\mem1[38][14] ), .IN2(n1015), .S(n7635), .Q(n14818) );
  MUX21X1 U11389 ( .IN1(\mem1[38][13] ), .IN2(n993), .S(n7635), .Q(n14817) );
  MUX21X1 U11390 ( .IN1(\mem1[38][12] ), .IN2(n971), .S(n7635), .Q(n14816) );
  MUX21X1 U11391 ( .IN1(\mem1[38][11] ), .IN2(n949), .S(n7635), .Q(n14815) );
  MUX21X1 U11392 ( .IN1(\mem1[38][10] ), .IN2(n927), .S(n7635), .Q(n14814) );
  MUX21X1 U11393 ( .IN1(\mem1[38][9] ), .IN2(n905), .S(n7635), .Q(n14813) );
  MUX21X1 U11394 ( .IN1(\mem1[38][8] ), .IN2(n883), .S(n7635), .Q(n14812) );
  AND2X1 U11395 ( .IN1(n7626), .IN2(n7118), .Q(n7635) );
  MUX21X1 U11396 ( .IN1(\mem1[37][15] ), .IN2(n1037), .S(n7636), .Q(n14811) );
  MUX21X1 U11397 ( .IN1(\mem1[37][14] ), .IN2(n1015), .S(n7636), .Q(n14810) );
  MUX21X1 U11398 ( .IN1(\mem1[37][13] ), .IN2(n993), .S(n7636), .Q(n14809) );
  MUX21X1 U11399 ( .IN1(\mem1[37][12] ), .IN2(n971), .S(n7636), .Q(n14808) );
  MUX21X1 U11400 ( .IN1(\mem1[37][11] ), .IN2(n949), .S(n7636), .Q(n14807) );
  MUX21X1 U11401 ( .IN1(\mem1[37][10] ), .IN2(n927), .S(n7636), .Q(n14806) );
  MUX21X1 U11402 ( .IN1(\mem1[37][9] ), .IN2(n905), .S(n7636), .Q(n14805) );
  MUX21X1 U11403 ( .IN1(\mem1[37][8] ), .IN2(n883), .S(n7636), .Q(n14804) );
  AND2X1 U11404 ( .IN1(n7626), .IN2(n7120), .Q(n7636) );
  MUX21X1 U11405 ( .IN1(\mem1[36][15] ), .IN2(n1037), .S(n7637), .Q(n14803) );
  MUX21X1 U11406 ( .IN1(\mem1[36][14] ), .IN2(n1015), .S(n7637), .Q(n14802) );
  MUX21X1 U11407 ( .IN1(\mem1[36][13] ), .IN2(n993), .S(n7637), .Q(n14801) );
  MUX21X1 U11408 ( .IN1(\mem1[36][12] ), .IN2(n971), .S(n7637), .Q(n14800) );
  MUX21X1 U11409 ( .IN1(\mem1[36][11] ), .IN2(n949), .S(n7637), .Q(n14799) );
  MUX21X1 U11410 ( .IN1(\mem1[36][10] ), .IN2(n927), .S(n7637), .Q(n14798) );
  MUX21X1 U11411 ( .IN1(\mem1[36][9] ), .IN2(n905), .S(n7637), .Q(n14797) );
  MUX21X1 U11412 ( .IN1(\mem1[36][8] ), .IN2(n883), .S(n7637), .Q(n14796) );
  AND2X1 U11413 ( .IN1(n7626), .IN2(n7122), .Q(n7637) );
  MUX21X1 U11414 ( .IN1(\mem1[35][15] ), .IN2(n1037), .S(n7638), .Q(n14795) );
  MUX21X1 U11415 ( .IN1(\mem1[35][14] ), .IN2(n1015), .S(n7638), .Q(n14794) );
  MUX21X1 U11416 ( .IN1(\mem1[35][13] ), .IN2(n993), .S(n7638), .Q(n14793) );
  MUX21X1 U11417 ( .IN1(\mem1[35][12] ), .IN2(n971), .S(n7638), .Q(n14792) );
  MUX21X1 U11418 ( .IN1(\mem1[35][11] ), .IN2(n949), .S(n7638), .Q(n14791) );
  MUX21X1 U11419 ( .IN1(\mem1[35][10] ), .IN2(n927), .S(n7638), .Q(n14790) );
  MUX21X1 U11420 ( .IN1(\mem1[35][9] ), .IN2(n905), .S(n7638), .Q(n14789) );
  MUX21X1 U11421 ( .IN1(\mem1[35][8] ), .IN2(n883), .S(n7638), .Q(n14788) );
  AND2X1 U11422 ( .IN1(n7626), .IN2(n7124), .Q(n7638) );
  MUX21X1 U11423 ( .IN1(\mem1[34][15] ), .IN2(n1037), .S(n7639), .Q(n14787) );
  MUX21X1 U11424 ( .IN1(\mem1[34][14] ), .IN2(n1015), .S(n7639), .Q(n14786) );
  MUX21X1 U11425 ( .IN1(\mem1[34][13] ), .IN2(n993), .S(n7639), .Q(n14785) );
  MUX21X1 U11426 ( .IN1(\mem1[34][12] ), .IN2(n971), .S(n7639), .Q(n14784) );
  MUX21X1 U11427 ( .IN1(\mem1[34][11] ), .IN2(n949), .S(n7639), .Q(n14783) );
  MUX21X1 U11428 ( .IN1(\mem1[34][10] ), .IN2(n927), .S(n7639), .Q(n14782) );
  MUX21X1 U11429 ( .IN1(\mem1[34][9] ), .IN2(n905), .S(n7639), .Q(n14781) );
  MUX21X1 U11430 ( .IN1(\mem1[34][8] ), .IN2(n883), .S(n7639), .Q(n14780) );
  AND2X1 U11431 ( .IN1(n7626), .IN2(n7126), .Q(n7639) );
  MUX21X1 U11432 ( .IN1(\mem1[33][15] ), .IN2(n1037), .S(n7640), .Q(n14779) );
  MUX21X1 U11433 ( .IN1(\mem1[33][14] ), .IN2(n1015), .S(n7640), .Q(n14778) );
  MUX21X1 U11434 ( .IN1(\mem1[33][13] ), .IN2(n993), .S(n7640), .Q(n14777) );
  MUX21X1 U11435 ( .IN1(\mem1[33][12] ), .IN2(n971), .S(n7640), .Q(n14776) );
  MUX21X1 U11436 ( .IN1(\mem1[33][11] ), .IN2(n949), .S(n7640), .Q(n14775) );
  MUX21X1 U11437 ( .IN1(\mem1[33][10] ), .IN2(n927), .S(n7640), .Q(n14774) );
  MUX21X1 U11438 ( .IN1(\mem1[33][9] ), .IN2(n905), .S(n7640), .Q(n14773) );
  MUX21X1 U11439 ( .IN1(\mem1[33][8] ), .IN2(n883), .S(n7640), .Q(n14772) );
  AND2X1 U11440 ( .IN1(n7626), .IN2(n7128), .Q(n7640) );
  MUX21X1 U11441 ( .IN1(\mem1[32][15] ), .IN2(n1037), .S(n7641), .Q(n14771) );
  MUX21X1 U11442 ( .IN1(\mem1[32][14] ), .IN2(n1015), .S(n7641), .Q(n14770) );
  MUX21X1 U11443 ( .IN1(\mem1[32][13] ), .IN2(n993), .S(n7641), .Q(n14769) );
  MUX21X1 U11444 ( .IN1(\mem1[32][12] ), .IN2(n971), .S(n7641), .Q(n14768) );
  MUX21X1 U11445 ( .IN1(\mem1[32][11] ), .IN2(n949), .S(n7641), .Q(n14767) );
  MUX21X1 U11446 ( .IN1(\mem1[32][10] ), .IN2(n927), .S(n7641), .Q(n14766) );
  MUX21X1 U11447 ( .IN1(\mem1[32][9] ), .IN2(n905), .S(n7641), .Q(n14765) );
  MUX21X1 U11448 ( .IN1(\mem1[32][8] ), .IN2(n883), .S(n7641), .Q(n14764) );
  AND2X1 U11449 ( .IN1(n7626), .IN2(n7130), .Q(n7641) );
  AND2X1 U11450 ( .IN1(n7420), .IN2(n7366), .Q(n7626) );
  MUX21X1 U11451 ( .IN1(\mem1[31][15] ), .IN2(n1037), .S(n7642), .Q(n14763) );
  MUX21X1 U11452 ( .IN1(\mem1[31][14] ), .IN2(n1015), .S(n7642), .Q(n14762) );
  MUX21X1 U11453 ( .IN1(\mem1[31][13] ), .IN2(n993), .S(n7642), .Q(n14761) );
  MUX21X1 U11454 ( .IN1(\mem1[31][12] ), .IN2(n971), .S(n7642), .Q(n14760) );
  MUX21X1 U11455 ( .IN1(\mem1[31][11] ), .IN2(n949), .S(n7642), .Q(n14759) );
  MUX21X1 U11456 ( .IN1(\mem1[31][10] ), .IN2(n927), .S(n7642), .Q(n14758) );
  MUX21X1 U11457 ( .IN1(\mem1[31][9] ), .IN2(n905), .S(n7642), .Q(n14757) );
  MUX21X1 U11458 ( .IN1(\mem1[31][8] ), .IN2(n883), .S(n7642), .Q(n14756) );
  AND2X1 U11459 ( .IN1(n7643), .IN2(n7099), .Q(n7642) );
  MUX21X1 U11460 ( .IN1(\mem1[30][15] ), .IN2(n1037), .S(n7644), .Q(n14755) );
  MUX21X1 U11461 ( .IN1(\mem1[30][14] ), .IN2(n1015), .S(n7644), .Q(n14754) );
  MUX21X1 U11462 ( .IN1(\mem1[30][13] ), .IN2(n993), .S(n7644), .Q(n14753) );
  MUX21X1 U11463 ( .IN1(\mem1[30][12] ), .IN2(n971), .S(n7644), .Q(n14752) );
  MUX21X1 U11464 ( .IN1(\mem1[30][11] ), .IN2(n949), .S(n7644), .Q(n14751) );
  MUX21X1 U11465 ( .IN1(\mem1[30][10] ), .IN2(n927), .S(n7644), .Q(n14750) );
  MUX21X1 U11466 ( .IN1(\mem1[30][9] ), .IN2(n905), .S(n7644), .Q(n14749) );
  MUX21X1 U11467 ( .IN1(\mem1[30][8] ), .IN2(n883), .S(n7644), .Q(n14748) );
  AND2X1 U11468 ( .IN1(n7643), .IN2(n7102), .Q(n7644) );
  MUX21X1 U11469 ( .IN1(\mem1[29][15] ), .IN2(n1037), .S(n7645), .Q(n14747) );
  MUX21X1 U11470 ( .IN1(\mem1[29][14] ), .IN2(n1015), .S(n7645), .Q(n14746) );
  MUX21X1 U11471 ( .IN1(\mem1[29][13] ), .IN2(n993), .S(n7645), .Q(n14745) );
  MUX21X1 U11472 ( .IN1(\mem1[29][12] ), .IN2(n971), .S(n7645), .Q(n14744) );
  MUX21X1 U11473 ( .IN1(\mem1[29][11] ), .IN2(n949), .S(n7645), .Q(n14743) );
  MUX21X1 U11474 ( .IN1(\mem1[29][10] ), .IN2(n927), .S(n7645), .Q(n14742) );
  MUX21X1 U11475 ( .IN1(\mem1[29][9] ), .IN2(n905), .S(n7645), .Q(n14741) );
  MUX21X1 U11476 ( .IN1(\mem1[29][8] ), .IN2(n883), .S(n7645), .Q(n14740) );
  AND2X1 U11477 ( .IN1(n7643), .IN2(n7104), .Q(n7645) );
  MUX21X1 U11478 ( .IN1(\mem1[28][15] ), .IN2(n1037), .S(n7646), .Q(n14739) );
  MUX21X1 U11479 ( .IN1(\mem1[28][14] ), .IN2(n1015), .S(n7646), .Q(n14738) );
  MUX21X1 U11480 ( .IN1(\mem1[28][13] ), .IN2(n993), .S(n7646), .Q(n14737) );
  MUX21X1 U11481 ( .IN1(\mem1[28][12] ), .IN2(n971), .S(n7646), .Q(n14736) );
  MUX21X1 U11482 ( .IN1(\mem1[28][11] ), .IN2(n949), .S(n7646), .Q(n14735) );
  MUX21X1 U11483 ( .IN1(\mem1[28][10] ), .IN2(n927), .S(n7646), .Q(n14734) );
  MUX21X1 U11484 ( .IN1(\mem1[28][9] ), .IN2(n905), .S(n7646), .Q(n14733) );
  MUX21X1 U11485 ( .IN1(\mem1[28][8] ), .IN2(n883), .S(n7646), .Q(n14732) );
  AND2X1 U11486 ( .IN1(n7643), .IN2(n7106), .Q(n7646) );
  MUX21X1 U11487 ( .IN1(\mem1[27][15] ), .IN2(n1038), .S(n7647), .Q(n14731) );
  MUX21X1 U11488 ( .IN1(\mem1[27][14] ), .IN2(n1016), .S(n7647), .Q(n14730) );
  MUX21X1 U11489 ( .IN1(\mem1[27][13] ), .IN2(n994), .S(n7647), .Q(n14729) );
  MUX21X1 U11490 ( .IN1(\mem1[27][12] ), .IN2(n972), .S(n7647), .Q(n14728) );
  MUX21X1 U11491 ( .IN1(\mem1[27][11] ), .IN2(n950), .S(n7647), .Q(n14727) );
  MUX21X1 U11492 ( .IN1(\mem1[27][10] ), .IN2(n928), .S(n7647), .Q(n14726) );
  MUX21X1 U11493 ( .IN1(\mem1[27][9] ), .IN2(n906), .S(n7647), .Q(n14725) );
  MUX21X1 U11494 ( .IN1(\mem1[27][8] ), .IN2(n884), .S(n7647), .Q(n14724) );
  AND2X1 U11495 ( .IN1(n7643), .IN2(n7108), .Q(n7647) );
  MUX21X1 U11496 ( .IN1(\mem1[26][15] ), .IN2(n1038), .S(n7648), .Q(n14723) );
  MUX21X1 U11497 ( .IN1(\mem1[26][14] ), .IN2(n1016), .S(n7648), .Q(n14722) );
  MUX21X1 U11498 ( .IN1(\mem1[26][13] ), .IN2(n994), .S(n7648), .Q(n14721) );
  MUX21X1 U11499 ( .IN1(\mem1[26][12] ), .IN2(n972), .S(n7648), .Q(n14720) );
  MUX21X1 U11500 ( .IN1(\mem1[26][11] ), .IN2(n950), .S(n7648), .Q(n14719) );
  MUX21X1 U11501 ( .IN1(\mem1[26][10] ), .IN2(n928), .S(n7648), .Q(n14718) );
  MUX21X1 U11502 ( .IN1(\mem1[26][9] ), .IN2(n906), .S(n7648), .Q(n14717) );
  MUX21X1 U11503 ( .IN1(\mem1[26][8] ), .IN2(n884), .S(n7648), .Q(n14716) );
  AND2X1 U11504 ( .IN1(n7643), .IN2(n7110), .Q(n7648) );
  MUX21X1 U11505 ( .IN1(\mem1[25][15] ), .IN2(n1038), .S(n7649), .Q(n14715) );
  MUX21X1 U11506 ( .IN1(\mem1[25][14] ), .IN2(n1016), .S(n7649), .Q(n14714) );
  MUX21X1 U11507 ( .IN1(\mem1[25][13] ), .IN2(n994), .S(n7649), .Q(n14713) );
  MUX21X1 U11508 ( .IN1(\mem1[25][12] ), .IN2(n972), .S(n7649), .Q(n14712) );
  MUX21X1 U11509 ( .IN1(\mem1[25][11] ), .IN2(n950), .S(n7649), .Q(n14711) );
  MUX21X1 U11510 ( .IN1(\mem1[25][10] ), .IN2(n928), .S(n7649), .Q(n14710) );
  MUX21X1 U11511 ( .IN1(\mem1[25][9] ), .IN2(n906), .S(n7649), .Q(n14709) );
  MUX21X1 U11512 ( .IN1(\mem1[25][8] ), .IN2(n884), .S(n7649), .Q(n14708) );
  AND2X1 U11513 ( .IN1(n7643), .IN2(n7112), .Q(n7649) );
  MUX21X1 U11514 ( .IN1(\mem1[24][15] ), .IN2(n1038), .S(n7650), .Q(n14707) );
  MUX21X1 U11515 ( .IN1(\mem1[24][14] ), .IN2(n1016), .S(n7650), .Q(n14706) );
  MUX21X1 U11516 ( .IN1(\mem1[24][13] ), .IN2(n994), .S(n7650), .Q(n14705) );
  MUX21X1 U11517 ( .IN1(\mem1[24][12] ), .IN2(n972), .S(n7650), .Q(n14704) );
  MUX21X1 U11518 ( .IN1(\mem1[24][11] ), .IN2(n950), .S(n7650), .Q(n14703) );
  MUX21X1 U11519 ( .IN1(\mem1[24][10] ), .IN2(n928), .S(n7650), .Q(n14702) );
  MUX21X1 U11520 ( .IN1(\mem1[24][9] ), .IN2(n906), .S(n7650), .Q(n14701) );
  MUX21X1 U11521 ( .IN1(\mem1[24][8] ), .IN2(n884), .S(n7650), .Q(n14700) );
  AND2X1 U11522 ( .IN1(n7643), .IN2(n7114), .Q(n7650) );
  MUX21X1 U11523 ( .IN1(\mem1[23][15] ), .IN2(n1038), .S(n7651), .Q(n14699) );
  MUX21X1 U11524 ( .IN1(\mem1[23][14] ), .IN2(n1016), .S(n7651), .Q(n14698) );
  MUX21X1 U11525 ( .IN1(\mem1[23][13] ), .IN2(n994), .S(n7651), .Q(n14697) );
  MUX21X1 U11526 ( .IN1(\mem1[23][12] ), .IN2(n972), .S(n7651), .Q(n14696) );
  MUX21X1 U11527 ( .IN1(\mem1[23][11] ), .IN2(n950), .S(n7651), .Q(n14695) );
  MUX21X1 U11528 ( .IN1(\mem1[23][10] ), .IN2(n928), .S(n7651), .Q(n14694) );
  MUX21X1 U11529 ( .IN1(\mem1[23][9] ), .IN2(n906), .S(n7651), .Q(n14693) );
  MUX21X1 U11530 ( .IN1(\mem1[23][8] ), .IN2(n884), .S(n7651), .Q(n14692) );
  AND2X1 U11531 ( .IN1(n7643), .IN2(n7116), .Q(n7651) );
  MUX21X1 U11532 ( .IN1(\mem1[22][15] ), .IN2(n1038), .S(n7652), .Q(n14691) );
  MUX21X1 U11533 ( .IN1(\mem1[22][14] ), .IN2(n1016), .S(n7652), .Q(n14690) );
  MUX21X1 U11534 ( .IN1(\mem1[22][13] ), .IN2(n994), .S(n7652), .Q(n14689) );
  MUX21X1 U11535 ( .IN1(\mem1[22][12] ), .IN2(n972), .S(n7652), .Q(n14688) );
  MUX21X1 U11536 ( .IN1(\mem1[22][11] ), .IN2(n950), .S(n7652), .Q(n14687) );
  MUX21X1 U11537 ( .IN1(\mem1[22][10] ), .IN2(n928), .S(n7652), .Q(n14686) );
  MUX21X1 U11538 ( .IN1(\mem1[22][9] ), .IN2(n906), .S(n7652), .Q(n14685) );
  MUX21X1 U11539 ( .IN1(\mem1[22][8] ), .IN2(n884), .S(n7652), .Q(n14684) );
  AND2X1 U11540 ( .IN1(n7643), .IN2(n7118), .Q(n7652) );
  MUX21X1 U11541 ( .IN1(\mem1[21][15] ), .IN2(n1038), .S(n7653), .Q(n14683) );
  MUX21X1 U11542 ( .IN1(\mem1[21][14] ), .IN2(n1016), .S(n7653), .Q(n14682) );
  MUX21X1 U11543 ( .IN1(\mem1[21][13] ), .IN2(n994), .S(n7653), .Q(n14681) );
  MUX21X1 U11544 ( .IN1(\mem1[21][12] ), .IN2(n972), .S(n7653), .Q(n14680) );
  MUX21X1 U11545 ( .IN1(\mem1[21][11] ), .IN2(n950), .S(n7653), .Q(n14679) );
  MUX21X1 U11546 ( .IN1(\mem1[21][10] ), .IN2(n928), .S(n7653), .Q(n14678) );
  MUX21X1 U11547 ( .IN1(\mem1[21][9] ), .IN2(n906), .S(n7653), .Q(n14677) );
  MUX21X1 U11548 ( .IN1(\mem1[21][8] ), .IN2(n884), .S(n7653), .Q(n14676) );
  AND2X1 U11549 ( .IN1(n7643), .IN2(n7120), .Q(n7653) );
  MUX21X1 U11550 ( .IN1(\mem1[20][15] ), .IN2(n1038), .S(n7654), .Q(n14675) );
  MUX21X1 U11551 ( .IN1(\mem1[20][14] ), .IN2(n1016), .S(n7654), .Q(n14674) );
  MUX21X1 U11552 ( .IN1(\mem1[20][13] ), .IN2(n994), .S(n7654), .Q(n14673) );
  MUX21X1 U11553 ( .IN1(\mem1[20][12] ), .IN2(n972), .S(n7654), .Q(n14672) );
  MUX21X1 U11554 ( .IN1(\mem1[20][11] ), .IN2(n950), .S(n7654), .Q(n14671) );
  MUX21X1 U11555 ( .IN1(\mem1[20][10] ), .IN2(n928), .S(n7654), .Q(n14670) );
  MUX21X1 U11556 ( .IN1(\mem1[20][9] ), .IN2(n906), .S(n7654), .Q(n14669) );
  MUX21X1 U11557 ( .IN1(\mem1[20][8] ), .IN2(n884), .S(n7654), .Q(n14668) );
  AND2X1 U11558 ( .IN1(n7643), .IN2(n7122), .Q(n7654) );
  MUX21X1 U11559 ( .IN1(\mem1[19][15] ), .IN2(n1038), .S(n7655), .Q(n14667) );
  MUX21X1 U11560 ( .IN1(\mem1[19][14] ), .IN2(n1016), .S(n7655), .Q(n14666) );
  MUX21X1 U11561 ( .IN1(\mem1[19][13] ), .IN2(n994), .S(n7655), .Q(n14665) );
  MUX21X1 U11562 ( .IN1(\mem1[19][12] ), .IN2(n972), .S(n7655), .Q(n14664) );
  MUX21X1 U11563 ( .IN1(\mem1[19][11] ), .IN2(n950), .S(n7655), .Q(n14663) );
  MUX21X1 U11564 ( .IN1(\mem1[19][10] ), .IN2(n928), .S(n7655), .Q(n14662) );
  MUX21X1 U11565 ( .IN1(\mem1[19][9] ), .IN2(n906), .S(n7655), .Q(n14661) );
  MUX21X1 U11566 ( .IN1(\mem1[19][8] ), .IN2(n884), .S(n7655), .Q(n14660) );
  AND2X1 U11567 ( .IN1(n7643), .IN2(n7124), .Q(n7655) );
  MUX21X1 U11568 ( .IN1(\mem1[18][15] ), .IN2(n1038), .S(n7656), .Q(n14659) );
  MUX21X1 U11569 ( .IN1(\mem1[18][14] ), .IN2(n1016), .S(n7656), .Q(n14658) );
  MUX21X1 U11570 ( .IN1(\mem1[18][13] ), .IN2(n994), .S(n7656), .Q(n14657) );
  MUX21X1 U11571 ( .IN1(\mem1[18][12] ), .IN2(n972), .S(n7656), .Q(n14656) );
  MUX21X1 U11572 ( .IN1(\mem1[18][11] ), .IN2(n950), .S(n7656), .Q(n14655) );
  MUX21X1 U11573 ( .IN1(\mem1[18][10] ), .IN2(n928), .S(n7656), .Q(n14654) );
  MUX21X1 U11574 ( .IN1(\mem1[18][9] ), .IN2(n906), .S(n7656), .Q(n14653) );
  MUX21X1 U11575 ( .IN1(\mem1[18][8] ), .IN2(n884), .S(n7656), .Q(n14652) );
  AND2X1 U11576 ( .IN1(n7643), .IN2(n7126), .Q(n7656) );
  MUX21X1 U11577 ( .IN1(\mem1[17][15] ), .IN2(n1038), .S(n7657), .Q(n14651) );
  MUX21X1 U11578 ( .IN1(\mem1[17][14] ), .IN2(n1016), .S(n7657), .Q(n14650) );
  MUX21X1 U11579 ( .IN1(\mem1[17][13] ), .IN2(n994), .S(n7657), .Q(n14649) );
  MUX21X1 U11580 ( .IN1(\mem1[17][12] ), .IN2(n972), .S(n7657), .Q(n14648) );
  MUX21X1 U11581 ( .IN1(\mem1[17][11] ), .IN2(n950), .S(n7657), .Q(n14647) );
  MUX21X1 U11582 ( .IN1(\mem1[17][10] ), .IN2(n928), .S(n7657), .Q(n14646) );
  MUX21X1 U11583 ( .IN1(\mem1[17][9] ), .IN2(n906), .S(n7657), .Q(n14645) );
  MUX21X1 U11584 ( .IN1(\mem1[17][8] ), .IN2(n884), .S(n7657), .Q(n14644) );
  AND2X1 U11585 ( .IN1(n7643), .IN2(n7128), .Q(n7657) );
  MUX21X1 U11586 ( .IN1(\mem1[16][15] ), .IN2(n1038), .S(n7658), .Q(n14643) );
  MUX21X1 U11587 ( .IN1(\mem1[16][14] ), .IN2(n1016), .S(n7658), .Q(n14642) );
  MUX21X1 U11588 ( .IN1(\mem1[16][13] ), .IN2(n994), .S(n7658), .Q(n14641) );
  MUX21X1 U11589 ( .IN1(\mem1[16][12] ), .IN2(n972), .S(n7658), .Q(n14640) );
  MUX21X1 U11590 ( .IN1(\mem1[16][11] ), .IN2(n950), .S(n7658), .Q(n14639) );
  MUX21X1 U11591 ( .IN1(\mem1[16][10] ), .IN2(n928), .S(n7658), .Q(n14638) );
  MUX21X1 U11592 ( .IN1(\mem1[16][9] ), .IN2(n906), .S(n7658), .Q(n14637) );
  MUX21X1 U11593 ( .IN1(\mem1[16][8] ), .IN2(n884), .S(n7658), .Q(n14636) );
  AND2X1 U11594 ( .IN1(n7643), .IN2(n7130), .Q(n7658) );
  AND2X1 U11595 ( .IN1(n7420), .IN2(n7384), .Q(n7643) );
  MUX21X1 U11596 ( .IN1(\mem1[15][15] ), .IN2(n1039), .S(n7659), .Q(n14635) );
  MUX21X1 U11597 ( .IN1(\mem1[15][14] ), .IN2(n1017), .S(n7659), .Q(n14634) );
  MUX21X1 U11598 ( .IN1(\mem1[15][13] ), .IN2(n995), .S(n7659), .Q(n14633) );
  MUX21X1 U11599 ( .IN1(\mem1[15][12] ), .IN2(n973), .S(n7659), .Q(n14632) );
  MUX21X1 U11600 ( .IN1(\mem1[15][11] ), .IN2(n951), .S(n7659), .Q(n14631) );
  MUX21X1 U11601 ( .IN1(\mem1[15][10] ), .IN2(n929), .S(n7659), .Q(n14630) );
  MUX21X1 U11602 ( .IN1(\mem1[15][9] ), .IN2(n907), .S(n7659), .Q(n14629) );
  MUX21X1 U11603 ( .IN1(\mem1[15][8] ), .IN2(n885), .S(n7659), .Q(n14628) );
  AND2X1 U11604 ( .IN1(n7660), .IN2(n7099), .Q(n7659) );
  MUX21X1 U11605 ( .IN1(\mem1[14][15] ), .IN2(n1039), .S(n7661), .Q(n14627) );
  MUX21X1 U11606 ( .IN1(\mem1[14][14] ), .IN2(n1017), .S(n7661), .Q(n14626) );
  MUX21X1 U11607 ( .IN1(\mem1[14][13] ), .IN2(n995), .S(n7661), .Q(n14625) );
  MUX21X1 U11608 ( .IN1(\mem1[14][12] ), .IN2(n973), .S(n7661), .Q(n14624) );
  MUX21X1 U11609 ( .IN1(\mem1[14][11] ), .IN2(n951), .S(n7661), .Q(n14623) );
  MUX21X1 U11610 ( .IN1(\mem1[14][10] ), .IN2(n929), .S(n7661), .Q(n14622) );
  MUX21X1 U11611 ( .IN1(\mem1[14][9] ), .IN2(n907), .S(n7661), .Q(n14621) );
  MUX21X1 U11612 ( .IN1(\mem1[14][8] ), .IN2(n885), .S(n7661), .Q(n14620) );
  AND2X1 U11613 ( .IN1(n7660), .IN2(n7102), .Q(n7661) );
  MUX21X1 U11614 ( .IN1(\mem1[13][15] ), .IN2(n1039), .S(n7662), .Q(n14619) );
  MUX21X1 U11615 ( .IN1(\mem1[13][14] ), .IN2(n1017), .S(n7662), .Q(n14618) );
  MUX21X1 U11616 ( .IN1(\mem1[13][13] ), .IN2(n995), .S(n7662), .Q(n14617) );
  MUX21X1 U11617 ( .IN1(\mem1[13][12] ), .IN2(n973), .S(n7662), .Q(n14616) );
  MUX21X1 U11618 ( .IN1(\mem1[13][11] ), .IN2(n951), .S(n7662), .Q(n14615) );
  MUX21X1 U11619 ( .IN1(\mem1[13][10] ), .IN2(n929), .S(n7662), .Q(n14614) );
  MUX21X1 U11620 ( .IN1(\mem1[13][9] ), .IN2(n907), .S(n7662), .Q(n14613) );
  MUX21X1 U11621 ( .IN1(\mem1[13][8] ), .IN2(n885), .S(n7662), .Q(n14612) );
  AND2X1 U11622 ( .IN1(n7660), .IN2(n7104), .Q(n7662) );
  MUX21X1 U11623 ( .IN1(\mem1[12][15] ), .IN2(n1039), .S(n7663), .Q(n14611) );
  MUX21X1 U11624 ( .IN1(\mem1[12][14] ), .IN2(n1017), .S(n7663), .Q(n14610) );
  MUX21X1 U11625 ( .IN1(\mem1[12][13] ), .IN2(n995), .S(n7663), .Q(n14609) );
  MUX21X1 U11626 ( .IN1(\mem1[12][12] ), .IN2(n973), .S(n7663), .Q(n14608) );
  MUX21X1 U11627 ( .IN1(\mem1[12][11] ), .IN2(n951), .S(n7663), .Q(n14607) );
  MUX21X1 U11628 ( .IN1(\mem1[12][10] ), .IN2(n929), .S(n7663), .Q(n14606) );
  MUX21X1 U11629 ( .IN1(\mem1[12][9] ), .IN2(n907), .S(n7663), .Q(n14605) );
  MUX21X1 U11630 ( .IN1(\mem1[12][8] ), .IN2(n885), .S(n7663), .Q(n14604) );
  AND2X1 U11631 ( .IN1(n7660), .IN2(n7106), .Q(n7663) );
  MUX21X1 U11632 ( .IN1(\mem1[11][15] ), .IN2(n1039), .S(n7664), .Q(n14603) );
  MUX21X1 U11633 ( .IN1(\mem1[11][14] ), .IN2(n1017), .S(n7664), .Q(n14602) );
  MUX21X1 U11634 ( .IN1(\mem1[11][13] ), .IN2(n995), .S(n7664), .Q(n14601) );
  MUX21X1 U11635 ( .IN1(\mem1[11][12] ), .IN2(n973), .S(n7664), .Q(n14600) );
  MUX21X1 U11636 ( .IN1(\mem1[11][11] ), .IN2(n951), .S(n7664), .Q(n14599) );
  MUX21X1 U11637 ( .IN1(\mem1[11][10] ), .IN2(n929), .S(n7664), .Q(n14598) );
  MUX21X1 U11638 ( .IN1(\mem1[11][9] ), .IN2(n907), .S(n7664), .Q(n14597) );
  MUX21X1 U11639 ( .IN1(\mem1[11][8] ), .IN2(n885), .S(n7664), .Q(n14596) );
  AND2X1 U11640 ( .IN1(n7660), .IN2(n7108), .Q(n7664) );
  MUX21X1 U11641 ( .IN1(\mem1[10][15] ), .IN2(n1039), .S(n7665), .Q(n14595) );
  MUX21X1 U11642 ( .IN1(\mem1[10][14] ), .IN2(n1017), .S(n7665), .Q(n14594) );
  MUX21X1 U11643 ( .IN1(\mem1[10][13] ), .IN2(n995), .S(n7665), .Q(n14593) );
  MUX21X1 U11644 ( .IN1(\mem1[10][12] ), .IN2(n973), .S(n7665), .Q(n14592) );
  MUX21X1 U11645 ( .IN1(\mem1[10][11] ), .IN2(n951), .S(n7665), .Q(n14591) );
  MUX21X1 U11646 ( .IN1(\mem1[10][10] ), .IN2(n929), .S(n7665), .Q(n14590) );
  MUX21X1 U11647 ( .IN1(\mem1[10][9] ), .IN2(n907), .S(n7665), .Q(n14589) );
  MUX21X1 U11648 ( .IN1(\mem1[10][8] ), .IN2(n885), .S(n7665), .Q(n14588) );
  AND2X1 U11649 ( .IN1(n7660), .IN2(n7110), .Q(n7665) );
  MUX21X1 U11650 ( .IN1(\mem1[9][15] ), .IN2(n1039), .S(n7666), .Q(n14587) );
  MUX21X1 U11651 ( .IN1(\mem1[9][14] ), .IN2(n1017), .S(n7666), .Q(n14586) );
  MUX21X1 U11652 ( .IN1(\mem1[9][13] ), .IN2(n995), .S(n7666), .Q(n14585) );
  MUX21X1 U11653 ( .IN1(\mem1[9][12] ), .IN2(n973), .S(n7666), .Q(n14584) );
  MUX21X1 U11654 ( .IN1(\mem1[9][11] ), .IN2(n951), .S(n7666), .Q(n14583) );
  MUX21X1 U11655 ( .IN1(\mem1[9][10] ), .IN2(n929), .S(n7666), .Q(n14582) );
  MUX21X1 U11656 ( .IN1(\mem1[9][9] ), .IN2(n907), .S(n7666), .Q(n14581) );
  MUX21X1 U11657 ( .IN1(\mem1[9][8] ), .IN2(n885), .S(n7666), .Q(n14580) );
  AND2X1 U11658 ( .IN1(n7660), .IN2(n7112), .Q(n7666) );
  MUX21X1 U11659 ( .IN1(\mem1[8][15] ), .IN2(n1039), .S(n7667), .Q(n14579) );
  MUX21X1 U11660 ( .IN1(\mem1[8][14] ), .IN2(n1017), .S(n7667), .Q(n14578) );
  MUX21X1 U11661 ( .IN1(\mem1[8][13] ), .IN2(n995), .S(n7667), .Q(n14577) );
  MUX21X1 U11662 ( .IN1(\mem1[8][12] ), .IN2(n973), .S(n7667), .Q(n14576) );
  MUX21X1 U11663 ( .IN1(\mem1[8][11] ), .IN2(n951), .S(n7667), .Q(n14575) );
  MUX21X1 U11664 ( .IN1(\mem1[8][10] ), .IN2(n929), .S(n7667), .Q(n14574) );
  MUX21X1 U11665 ( .IN1(\mem1[8][9] ), .IN2(n907), .S(n7667), .Q(n14573) );
  MUX21X1 U11666 ( .IN1(\mem1[8][8] ), .IN2(n885), .S(n7667), .Q(n14572) );
  AND2X1 U11667 ( .IN1(n7660), .IN2(n7114), .Q(n7667) );
  MUX21X1 U11668 ( .IN1(\mem1[7][15] ), .IN2(n1039), .S(n7668), .Q(n14571) );
  MUX21X1 U11669 ( .IN1(\mem1[7][14] ), .IN2(n1017), .S(n7668), .Q(n14570) );
  MUX21X1 U11670 ( .IN1(\mem1[7][13] ), .IN2(n995), .S(n7668), .Q(n14569) );
  MUX21X1 U11671 ( .IN1(\mem1[7][12] ), .IN2(n973), .S(n7668), .Q(n14568) );
  MUX21X1 U11672 ( .IN1(\mem1[7][11] ), .IN2(n951), .S(n7668), .Q(n14567) );
  MUX21X1 U11673 ( .IN1(\mem1[7][10] ), .IN2(n929), .S(n7668), .Q(n14566) );
  MUX21X1 U11674 ( .IN1(\mem1[7][9] ), .IN2(n907), .S(n7668), .Q(n14565) );
  MUX21X1 U11675 ( .IN1(\mem1[7][8] ), .IN2(n885), .S(n7668), .Q(n14564) );
  AND2X1 U11676 ( .IN1(n7660), .IN2(n7116), .Q(n7668) );
  MUX21X1 U11677 ( .IN1(\mem1[6][15] ), .IN2(n1039), .S(n7669), .Q(n14563) );
  MUX21X1 U11678 ( .IN1(\mem1[6][14] ), .IN2(n1017), .S(n7669), .Q(n14562) );
  MUX21X1 U11679 ( .IN1(\mem1[6][13] ), .IN2(n995), .S(n7669), .Q(n14561) );
  MUX21X1 U11680 ( .IN1(\mem1[6][12] ), .IN2(n973), .S(n7669), .Q(n14560) );
  MUX21X1 U11681 ( .IN1(\mem1[6][11] ), .IN2(n951), .S(n7669), .Q(n14559) );
  MUX21X1 U11682 ( .IN1(\mem1[6][10] ), .IN2(n929), .S(n7669), .Q(n14558) );
  MUX21X1 U11683 ( .IN1(\mem1[6][9] ), .IN2(n907), .S(n7669), .Q(n14557) );
  MUX21X1 U11684 ( .IN1(\mem1[6][8] ), .IN2(n885), .S(n7669), .Q(n14556) );
  AND2X1 U11685 ( .IN1(n7660), .IN2(n7118), .Q(n7669) );
  MUX21X1 U11686 ( .IN1(\mem1[5][15] ), .IN2(n1039), .S(n7670), .Q(n14555) );
  MUX21X1 U11687 ( .IN1(\mem1[5][14] ), .IN2(n1017), .S(n7670), .Q(n14554) );
  MUX21X1 U11688 ( .IN1(\mem1[5][13] ), .IN2(n995), .S(n7670), .Q(n14553) );
  MUX21X1 U11689 ( .IN1(\mem1[5][12] ), .IN2(n973), .S(n7670), .Q(n14552) );
  MUX21X1 U11690 ( .IN1(\mem1[5][11] ), .IN2(n951), .S(n7670), .Q(n14551) );
  MUX21X1 U11691 ( .IN1(\mem1[5][10] ), .IN2(n929), .S(n7670), .Q(n14550) );
  MUX21X1 U11692 ( .IN1(\mem1[5][9] ), .IN2(n907), .S(n7670), .Q(n14549) );
  MUX21X1 U11693 ( .IN1(\mem1[5][8] ), .IN2(n885), .S(n7670), .Q(n14548) );
  AND2X1 U11694 ( .IN1(n7660), .IN2(n7120), .Q(n7670) );
  MUX21X1 U11695 ( .IN1(\mem1[4][15] ), .IN2(n1039), .S(n7671), .Q(n14547) );
  MUX21X1 U11696 ( .IN1(\mem1[4][14] ), .IN2(n1017), .S(n7671), .Q(n14546) );
  MUX21X1 U11697 ( .IN1(\mem1[4][13] ), .IN2(n995), .S(n7671), .Q(n14545) );
  MUX21X1 U11698 ( .IN1(\mem1[4][12] ), .IN2(n973), .S(n7671), .Q(n14544) );
  MUX21X1 U11699 ( .IN1(\mem1[4][11] ), .IN2(n951), .S(n7671), .Q(n14543) );
  MUX21X1 U11700 ( .IN1(\mem1[4][10] ), .IN2(n929), .S(n7671), .Q(n14542) );
  MUX21X1 U11701 ( .IN1(\mem1[4][9] ), .IN2(n907), .S(n7671), .Q(n14541) );
  MUX21X1 U11702 ( .IN1(\mem1[4][8] ), .IN2(n885), .S(n7671), .Q(n14540) );
  AND2X1 U11703 ( .IN1(n7660), .IN2(n7122), .Q(n7671) );
  MUX21X1 U11704 ( .IN1(\mem1[3][15] ), .IN2(n1040), .S(n7672), .Q(n14539) );
  MUX21X1 U11705 ( .IN1(\mem1[3][14] ), .IN2(n1018), .S(n7672), .Q(n14538) );
  MUX21X1 U11706 ( .IN1(\mem1[3][13] ), .IN2(n996), .S(n7672), .Q(n14537) );
  MUX21X1 U11707 ( .IN1(\mem1[3][12] ), .IN2(n974), .S(n7672), .Q(n14536) );
  MUX21X1 U11708 ( .IN1(\mem1[3][11] ), .IN2(n952), .S(n7672), .Q(n14535) );
  MUX21X1 U11709 ( .IN1(\mem1[3][10] ), .IN2(n930), .S(n7672), .Q(n14534) );
  MUX21X1 U11710 ( .IN1(\mem1[3][9] ), .IN2(n908), .S(n7672), .Q(n14533) );
  MUX21X1 U11711 ( .IN1(\mem1[3][8] ), .IN2(n886), .S(n7672), .Q(n14532) );
  AND2X1 U11712 ( .IN1(n7660), .IN2(n7124), .Q(n7672) );
  MUX21X1 U11713 ( .IN1(\mem1[2][15] ), .IN2(n1040), .S(n7673), .Q(n14531) );
  MUX21X1 U11714 ( .IN1(\mem1[2][14] ), .IN2(n1018), .S(n7673), .Q(n14530) );
  MUX21X1 U11715 ( .IN1(\mem1[2][13] ), .IN2(n996), .S(n7673), .Q(n14529) );
  MUX21X1 U11716 ( .IN1(\mem1[2][12] ), .IN2(n974), .S(n7673), .Q(n14528) );
  MUX21X1 U11717 ( .IN1(\mem1[2][11] ), .IN2(n952), .S(n7673), .Q(n14527) );
  MUX21X1 U11718 ( .IN1(\mem1[2][10] ), .IN2(n930), .S(n7673), .Q(n14526) );
  MUX21X1 U11719 ( .IN1(\mem1[2][9] ), .IN2(n908), .S(n7673), .Q(n14525) );
  MUX21X1 U11720 ( .IN1(\mem1[2][8] ), .IN2(n886), .S(n7673), .Q(n14524) );
  AND2X1 U11721 ( .IN1(n7660), .IN2(n7126), .Q(n7673) );
  MUX21X1 U11722 ( .IN1(\mem1[1][15] ), .IN2(n1040), .S(n7674), .Q(n14523) );
  MUX21X1 U11723 ( .IN1(\mem1[1][14] ), .IN2(n1018), .S(n7674), .Q(n14522) );
  MUX21X1 U11724 ( .IN1(\mem1[1][13] ), .IN2(n996), .S(n7674), .Q(n14521) );
  MUX21X1 U11725 ( .IN1(\mem1[1][12] ), .IN2(n974), .S(n7674), .Q(n14520) );
  MUX21X1 U11726 ( .IN1(\mem1[1][11] ), .IN2(n952), .S(n7674), .Q(n14519) );
  MUX21X1 U11727 ( .IN1(\mem1[1][10] ), .IN2(n930), .S(n7674), .Q(n14518) );
  MUX21X1 U11728 ( .IN1(\mem1[1][9] ), .IN2(n908), .S(n7674), .Q(n14517) );
  MUX21X1 U11729 ( .IN1(\mem1[1][8] ), .IN2(n886), .S(n7674), .Q(n14516) );
  AND2X1 U11730 ( .IN1(n7660), .IN2(n7128), .Q(n7674) );
  MUX21X1 U11731 ( .IN1(\mem1[0][15] ), .IN2(n1040), .S(n7675), .Q(n14515) );
  MUX21X1 U11732 ( .IN1(\mem1[0][14] ), .IN2(n1018), .S(n7675), .Q(n14514) );
  MUX21X1 U11733 ( .IN1(\mem1[0][13] ), .IN2(n996), .S(n7675), .Q(n14513) );
  MUX21X1 U11734 ( .IN1(\mem1[0][12] ), .IN2(n974), .S(n7675), .Q(n14512) );
  MUX21X1 U11735 ( .IN1(\mem1[0][11] ), .IN2(n952), .S(n7675), .Q(n14511) );
  MUX21X1 U11736 ( .IN1(\mem1[0][10] ), .IN2(n930), .S(n7675), .Q(n14510) );
  MUX21X1 U11737 ( .IN1(\mem1[0][9] ), .IN2(n908), .S(n7675), .Q(n14509) );
  MUX21X1 U11738 ( .IN1(\mem1[0][8] ), .IN2(n886), .S(n7675), .Q(n14508) );
  AND2X1 U11739 ( .IN1(n7660), .IN2(n7130), .Q(n7675) );
  AND2X1 U11740 ( .IN1(n7420), .IN2(n7402), .Q(n7660) );
  AND2X1 U11741 ( .IN1(we[1]), .IN2(ce), .Q(n7420) );
  MUX21X1 U11742 ( .IN1(\mem3[255][31] ), .IN2(n1371), .S(n7676), .Q(n14507)
         );
  MUX21X1 U11743 ( .IN1(\mem3[255][30] ), .IN2(n1349), .S(n7676), .Q(n14506)
         );
  MUX21X1 U11744 ( .IN1(\mem3[255][29] ), .IN2(n1327), .S(n7676), .Q(n14505)
         );
  MUX21X1 U11745 ( .IN1(\mem3[255][28] ), .IN2(n1305), .S(n7676), .Q(n14504)
         );
  MUX21X1 U11746 ( .IN1(\mem3[255][27] ), .IN2(n1283), .S(n7676), .Q(n14503)
         );
  MUX21X1 U11747 ( .IN1(\mem3[255][26] ), .IN2(n1261), .S(n7676), .Q(n14502)
         );
  MUX21X1 U11748 ( .IN1(\mem3[255][25] ), .IN2(n1239), .S(n7676), .Q(n14501)
         );
  MUX21X1 U11749 ( .IN1(\mem3[255][24] ), .IN2(n1217), .S(n7676), .Q(n14500)
         );
  AND2X1 U11750 ( .IN1(n7677), .IN2(n7099), .Q(n7676) );
  MUX21X1 U11751 ( .IN1(\mem3[254][31] ), .IN2(n1371), .S(n7678), .Q(n14499)
         );
  MUX21X1 U11752 ( .IN1(\mem3[254][30] ), .IN2(n1349), .S(n7678), .Q(n14498)
         );
  MUX21X1 U11753 ( .IN1(\mem3[254][29] ), .IN2(n1327), .S(n7678), .Q(n14497)
         );
  MUX21X1 U11754 ( .IN1(\mem3[254][28] ), .IN2(n1305), .S(n7678), .Q(n14496)
         );
  MUX21X1 U11755 ( .IN1(\mem3[254][27] ), .IN2(n1283), .S(n7678), .Q(n14495)
         );
  MUX21X1 U11756 ( .IN1(\mem3[254][26] ), .IN2(n1261), .S(n7678), .Q(n14494)
         );
  MUX21X1 U11757 ( .IN1(\mem3[254][25] ), .IN2(n1239), .S(n7678), .Q(n14493)
         );
  MUX21X1 U11758 ( .IN1(\mem3[254][24] ), .IN2(n1217), .S(n7678), .Q(n14492)
         );
  AND2X1 U11759 ( .IN1(n7677), .IN2(n7102), .Q(n7678) );
  MUX21X1 U11760 ( .IN1(\mem3[253][31] ), .IN2(n1371), .S(n7679), .Q(n14491)
         );
  MUX21X1 U11761 ( .IN1(\mem3[253][30] ), .IN2(n1349), .S(n7679), .Q(n14490)
         );
  MUX21X1 U11762 ( .IN1(\mem3[253][29] ), .IN2(n1327), .S(n7679), .Q(n14489)
         );
  MUX21X1 U11763 ( .IN1(\mem3[253][28] ), .IN2(n1305), .S(n7679), .Q(n14488)
         );
  MUX21X1 U11764 ( .IN1(\mem3[253][27] ), .IN2(n1283), .S(n7679), .Q(n14487)
         );
  MUX21X1 U11765 ( .IN1(\mem3[253][26] ), .IN2(n1261), .S(n7679), .Q(n14486)
         );
  MUX21X1 U11766 ( .IN1(\mem3[253][25] ), .IN2(n1239), .S(n7679), .Q(n14485)
         );
  MUX21X1 U11767 ( .IN1(\mem3[253][24] ), .IN2(n1217), .S(n7679), .Q(n14484)
         );
  AND2X1 U11768 ( .IN1(n7677), .IN2(n7104), .Q(n7679) );
  MUX21X1 U11769 ( .IN1(\mem3[252][31] ), .IN2(n1371), .S(n7680), .Q(n14483)
         );
  MUX21X1 U11770 ( .IN1(\mem3[252][30] ), .IN2(n1349), .S(n7680), .Q(n14482)
         );
  MUX21X1 U11771 ( .IN1(\mem3[252][29] ), .IN2(n1327), .S(n7680), .Q(n14481)
         );
  MUX21X1 U11772 ( .IN1(\mem3[252][28] ), .IN2(n1305), .S(n7680), .Q(n14480)
         );
  MUX21X1 U11773 ( .IN1(\mem3[252][27] ), .IN2(n1283), .S(n7680), .Q(n14479)
         );
  MUX21X1 U11774 ( .IN1(\mem3[252][26] ), .IN2(n1261), .S(n7680), .Q(n14478)
         );
  MUX21X1 U11775 ( .IN1(\mem3[252][25] ), .IN2(n1239), .S(n7680), .Q(n14477)
         );
  MUX21X1 U11776 ( .IN1(\mem3[252][24] ), .IN2(n1217), .S(n7680), .Q(n14476)
         );
  AND2X1 U11777 ( .IN1(n7677), .IN2(n7106), .Q(n7680) );
  MUX21X1 U11778 ( .IN1(\mem3[251][31] ), .IN2(n1371), .S(n7681), .Q(n14475)
         );
  MUX21X1 U11779 ( .IN1(\mem3[251][30] ), .IN2(n1349), .S(n7681), .Q(n14474)
         );
  MUX21X1 U11780 ( .IN1(\mem3[251][29] ), .IN2(n1327), .S(n7681), .Q(n14473)
         );
  MUX21X1 U11781 ( .IN1(\mem3[251][28] ), .IN2(n1305), .S(n7681), .Q(n14472)
         );
  MUX21X1 U11782 ( .IN1(\mem3[251][27] ), .IN2(n1283), .S(n7681), .Q(n14471)
         );
  MUX21X1 U11783 ( .IN1(\mem3[251][26] ), .IN2(n1261), .S(n7681), .Q(n14470)
         );
  MUX21X1 U11784 ( .IN1(\mem3[251][25] ), .IN2(n1239), .S(n7681), .Q(n14469)
         );
  MUX21X1 U11785 ( .IN1(\mem3[251][24] ), .IN2(n1217), .S(n7681), .Q(n14468)
         );
  AND2X1 U11786 ( .IN1(n7677), .IN2(n7108), .Q(n7681) );
  MUX21X1 U11787 ( .IN1(\mem3[250][31] ), .IN2(n1371), .S(n7682), .Q(n14467)
         );
  MUX21X1 U11788 ( .IN1(\mem3[250][30] ), .IN2(n1349), .S(n7682), .Q(n14466)
         );
  MUX21X1 U11789 ( .IN1(\mem3[250][29] ), .IN2(n1327), .S(n7682), .Q(n14465)
         );
  MUX21X1 U11790 ( .IN1(\mem3[250][28] ), .IN2(n1305), .S(n7682), .Q(n14464)
         );
  MUX21X1 U11791 ( .IN1(\mem3[250][27] ), .IN2(n1283), .S(n7682), .Q(n14463)
         );
  MUX21X1 U11792 ( .IN1(\mem3[250][26] ), .IN2(n1261), .S(n7682), .Q(n14462)
         );
  MUX21X1 U11793 ( .IN1(\mem3[250][25] ), .IN2(n1239), .S(n7682), .Q(n14461)
         );
  MUX21X1 U11794 ( .IN1(\mem3[250][24] ), .IN2(n1217), .S(n7682), .Q(n14460)
         );
  AND2X1 U11795 ( .IN1(n7677), .IN2(n7110), .Q(n7682) );
  MUX21X1 U11796 ( .IN1(\mem3[249][31] ), .IN2(n1371), .S(n7683), .Q(n14459)
         );
  MUX21X1 U11797 ( .IN1(\mem3[249][30] ), .IN2(n1349), .S(n7683), .Q(n14458)
         );
  MUX21X1 U11798 ( .IN1(\mem3[249][29] ), .IN2(n1327), .S(n7683), .Q(n14457)
         );
  MUX21X1 U11799 ( .IN1(\mem3[249][28] ), .IN2(n1305), .S(n7683), .Q(n14456)
         );
  MUX21X1 U11800 ( .IN1(\mem3[249][27] ), .IN2(n1283), .S(n7683), .Q(n14455)
         );
  MUX21X1 U11801 ( .IN1(\mem3[249][26] ), .IN2(n1261), .S(n7683), .Q(n14454)
         );
  MUX21X1 U11802 ( .IN1(\mem3[249][25] ), .IN2(n1239), .S(n7683), .Q(n14453)
         );
  MUX21X1 U11803 ( .IN1(\mem3[249][24] ), .IN2(n1217), .S(n7683), .Q(n14452)
         );
  AND2X1 U11804 ( .IN1(n7677), .IN2(n7112), .Q(n7683) );
  MUX21X1 U11805 ( .IN1(\mem3[248][31] ), .IN2(n1371), .S(n7684), .Q(n14451)
         );
  MUX21X1 U11806 ( .IN1(\mem3[248][30] ), .IN2(n1349), .S(n7684), .Q(n14450)
         );
  MUX21X1 U11807 ( .IN1(\mem3[248][29] ), .IN2(n1327), .S(n7684), .Q(n14449)
         );
  MUX21X1 U11808 ( .IN1(\mem3[248][28] ), .IN2(n1305), .S(n7684), .Q(n14448)
         );
  MUX21X1 U11809 ( .IN1(\mem3[248][27] ), .IN2(n1283), .S(n7684), .Q(n14447)
         );
  MUX21X1 U11810 ( .IN1(\mem3[248][26] ), .IN2(n1261), .S(n7684), .Q(n14446)
         );
  MUX21X1 U11811 ( .IN1(\mem3[248][25] ), .IN2(n1239), .S(n7684), .Q(n14445)
         );
  MUX21X1 U11812 ( .IN1(\mem3[248][24] ), .IN2(n1217), .S(n7684), .Q(n14444)
         );
  AND2X1 U11813 ( .IN1(n7677), .IN2(n7114), .Q(n7684) );
  MUX21X1 U11814 ( .IN1(\mem3[247][31] ), .IN2(n1371), .S(n7685), .Q(n14443)
         );
  MUX21X1 U11815 ( .IN1(\mem3[247][30] ), .IN2(n1349), .S(n7685), .Q(n14442)
         );
  MUX21X1 U11816 ( .IN1(\mem3[247][29] ), .IN2(n1327), .S(n7685), .Q(n14441)
         );
  MUX21X1 U11817 ( .IN1(\mem3[247][28] ), .IN2(n1305), .S(n7685), .Q(n14440)
         );
  MUX21X1 U11818 ( .IN1(\mem3[247][27] ), .IN2(n1283), .S(n7685), .Q(n14439)
         );
  MUX21X1 U11819 ( .IN1(\mem3[247][26] ), .IN2(n1261), .S(n7685), .Q(n14438)
         );
  MUX21X1 U11820 ( .IN1(\mem3[247][25] ), .IN2(n1239), .S(n7685), .Q(n14437)
         );
  MUX21X1 U11821 ( .IN1(\mem3[247][24] ), .IN2(n1217), .S(n7685), .Q(n14436)
         );
  AND2X1 U11822 ( .IN1(n7677), .IN2(n7116), .Q(n7685) );
  MUX21X1 U11823 ( .IN1(\mem3[246][31] ), .IN2(n1371), .S(n7686), .Q(n14435)
         );
  MUX21X1 U11824 ( .IN1(\mem3[246][30] ), .IN2(n1349), .S(n7686), .Q(n14434)
         );
  MUX21X1 U11825 ( .IN1(\mem3[246][29] ), .IN2(n1327), .S(n7686), .Q(n14433)
         );
  MUX21X1 U11826 ( .IN1(\mem3[246][28] ), .IN2(n1305), .S(n7686), .Q(n14432)
         );
  MUX21X1 U11827 ( .IN1(\mem3[246][27] ), .IN2(n1283), .S(n7686), .Q(n14431)
         );
  MUX21X1 U11828 ( .IN1(\mem3[246][26] ), .IN2(n1261), .S(n7686), .Q(n14430)
         );
  MUX21X1 U11829 ( .IN1(\mem3[246][25] ), .IN2(n1239), .S(n7686), .Q(n14429)
         );
  MUX21X1 U11830 ( .IN1(\mem3[246][24] ), .IN2(n1217), .S(n7686), .Q(n14428)
         );
  AND2X1 U11831 ( .IN1(n7677), .IN2(n7118), .Q(n7686) );
  MUX21X1 U11832 ( .IN1(\mem3[245][31] ), .IN2(n1371), .S(n7687), .Q(n14427)
         );
  MUX21X1 U11833 ( .IN1(\mem3[245][30] ), .IN2(n1349), .S(n7687), .Q(n14426)
         );
  MUX21X1 U11834 ( .IN1(\mem3[245][29] ), .IN2(n1327), .S(n7687), .Q(n14425)
         );
  MUX21X1 U11835 ( .IN1(\mem3[245][28] ), .IN2(n1305), .S(n7687), .Q(n14424)
         );
  MUX21X1 U11836 ( .IN1(\mem3[245][27] ), .IN2(n1283), .S(n7687), .Q(n14423)
         );
  MUX21X1 U11837 ( .IN1(\mem3[245][26] ), .IN2(n1261), .S(n7687), .Q(n14422)
         );
  MUX21X1 U11838 ( .IN1(\mem3[245][25] ), .IN2(n1239), .S(n7687), .Q(n14421)
         );
  MUX21X1 U11839 ( .IN1(\mem3[245][24] ), .IN2(n1217), .S(n7687), .Q(n14420)
         );
  AND2X1 U11840 ( .IN1(n7677), .IN2(n7120), .Q(n7687) );
  MUX21X1 U11841 ( .IN1(\mem3[244][31] ), .IN2(n1371), .S(n7688), .Q(n14419)
         );
  MUX21X1 U11842 ( .IN1(\mem3[244][30] ), .IN2(n1349), .S(n7688), .Q(n14418)
         );
  MUX21X1 U11843 ( .IN1(\mem3[244][29] ), .IN2(n1327), .S(n7688), .Q(n14417)
         );
  MUX21X1 U11844 ( .IN1(\mem3[244][28] ), .IN2(n1305), .S(n7688), .Q(n14416)
         );
  MUX21X1 U11845 ( .IN1(\mem3[244][27] ), .IN2(n1283), .S(n7688), .Q(n14415)
         );
  MUX21X1 U11846 ( .IN1(\mem3[244][26] ), .IN2(n1261), .S(n7688), .Q(n14414)
         );
  MUX21X1 U11847 ( .IN1(\mem3[244][25] ), .IN2(n1239), .S(n7688), .Q(n14413)
         );
  MUX21X1 U11848 ( .IN1(\mem3[244][24] ), .IN2(n1217), .S(n7688), .Q(n14412)
         );
  AND2X1 U11849 ( .IN1(n7677), .IN2(n7122), .Q(n7688) );
  MUX21X1 U11850 ( .IN1(\mem3[243][31] ), .IN2(n1372), .S(n7689), .Q(n14411)
         );
  MUX21X1 U11851 ( .IN1(\mem3[243][30] ), .IN2(n1350), .S(n7689), .Q(n14410)
         );
  MUX21X1 U11852 ( .IN1(\mem3[243][29] ), .IN2(n1328), .S(n7689), .Q(n14409)
         );
  MUX21X1 U11853 ( .IN1(\mem3[243][28] ), .IN2(n1306), .S(n7689), .Q(n14408)
         );
  MUX21X1 U11854 ( .IN1(\mem3[243][27] ), .IN2(n1284), .S(n7689), .Q(n14407)
         );
  MUX21X1 U11855 ( .IN1(\mem3[243][26] ), .IN2(n1262), .S(n7689), .Q(n14406)
         );
  MUX21X1 U11856 ( .IN1(\mem3[243][25] ), .IN2(n1240), .S(n7689), .Q(n14405)
         );
  MUX21X1 U11857 ( .IN1(\mem3[243][24] ), .IN2(n1218), .S(n7689), .Q(n14404)
         );
  AND2X1 U11858 ( .IN1(n7677), .IN2(n7124), .Q(n7689) );
  MUX21X1 U11859 ( .IN1(\mem3[242][31] ), .IN2(n1372), .S(n7690), .Q(n14403)
         );
  MUX21X1 U11860 ( .IN1(\mem3[242][30] ), .IN2(n1350), .S(n7690), .Q(n14402)
         );
  MUX21X1 U11861 ( .IN1(\mem3[242][29] ), .IN2(n1328), .S(n7690), .Q(n14401)
         );
  MUX21X1 U11862 ( .IN1(\mem3[242][28] ), .IN2(n1306), .S(n7690), .Q(n14400)
         );
  MUX21X1 U11863 ( .IN1(\mem3[242][27] ), .IN2(n1284), .S(n7690), .Q(n14399)
         );
  MUX21X1 U11864 ( .IN1(\mem3[242][26] ), .IN2(n1262), .S(n7690), .Q(n14398)
         );
  MUX21X1 U11865 ( .IN1(\mem3[242][25] ), .IN2(n1240), .S(n7690), .Q(n14397)
         );
  MUX21X1 U11866 ( .IN1(\mem3[242][24] ), .IN2(n1218), .S(n7690), .Q(n14396)
         );
  AND2X1 U11867 ( .IN1(n7677), .IN2(n7126), .Q(n7690) );
  MUX21X1 U11868 ( .IN1(\mem3[241][31] ), .IN2(n1372), .S(n7691), .Q(n14395)
         );
  MUX21X1 U11869 ( .IN1(\mem3[241][30] ), .IN2(n1350), .S(n7691), .Q(n14394)
         );
  MUX21X1 U11870 ( .IN1(\mem3[241][29] ), .IN2(n1328), .S(n7691), .Q(n14393)
         );
  MUX21X1 U11871 ( .IN1(\mem3[241][28] ), .IN2(n1306), .S(n7691), .Q(n14392)
         );
  MUX21X1 U11872 ( .IN1(\mem3[241][27] ), .IN2(n1284), .S(n7691), .Q(n14391)
         );
  MUX21X1 U11873 ( .IN1(\mem3[241][26] ), .IN2(n1262), .S(n7691), .Q(n14390)
         );
  MUX21X1 U11874 ( .IN1(\mem3[241][25] ), .IN2(n1240), .S(n7691), .Q(n14389)
         );
  MUX21X1 U11875 ( .IN1(\mem3[241][24] ), .IN2(n1218), .S(n7691), .Q(n14388)
         );
  AND2X1 U11876 ( .IN1(n7677), .IN2(n7128), .Q(n7691) );
  MUX21X1 U11877 ( .IN1(\mem3[240][31] ), .IN2(n1372), .S(n7692), .Q(n14387)
         );
  MUX21X1 U11878 ( .IN1(\mem3[240][30] ), .IN2(n1350), .S(n7692), .Q(n14386)
         );
  MUX21X1 U11879 ( .IN1(\mem3[240][29] ), .IN2(n1328), .S(n7692), .Q(n14385)
         );
  MUX21X1 U11880 ( .IN1(\mem3[240][28] ), .IN2(n1306), .S(n7692), .Q(n14384)
         );
  MUX21X1 U11881 ( .IN1(\mem3[240][27] ), .IN2(n1284), .S(n7692), .Q(n14383)
         );
  MUX21X1 U11882 ( .IN1(\mem3[240][26] ), .IN2(n1262), .S(n7692), .Q(n14382)
         );
  MUX21X1 U11883 ( .IN1(\mem3[240][25] ), .IN2(n1240), .S(n7692), .Q(n14381)
         );
  MUX21X1 U11884 ( .IN1(\mem3[240][24] ), .IN2(n1218), .S(n7692), .Q(n14380)
         );
  AND2X1 U11885 ( .IN1(n7677), .IN2(n7130), .Q(n7692) );
  AND2X1 U11886 ( .IN1(n7693), .IN2(n7131), .Q(n7677) );
  MUX21X1 U11887 ( .IN1(\mem3[239][31] ), .IN2(n1372), .S(n7694), .Q(n14379)
         );
  MUX21X1 U11888 ( .IN1(\mem3[239][30] ), .IN2(n1350), .S(n7694), .Q(n14378)
         );
  MUX21X1 U11889 ( .IN1(\mem3[239][29] ), .IN2(n1328), .S(n7694), .Q(n14377)
         );
  MUX21X1 U11890 ( .IN1(\mem3[239][28] ), .IN2(n1306), .S(n7694), .Q(n14376)
         );
  MUX21X1 U11891 ( .IN1(\mem3[239][27] ), .IN2(n1284), .S(n7694), .Q(n14375)
         );
  MUX21X1 U11892 ( .IN1(\mem3[239][26] ), .IN2(n1262), .S(n7694), .Q(n14374)
         );
  MUX21X1 U11893 ( .IN1(\mem3[239][25] ), .IN2(n1240), .S(n7694), .Q(n14373)
         );
  MUX21X1 U11894 ( .IN1(\mem3[239][24] ), .IN2(n1218), .S(n7694), .Q(n14372)
         );
  AND2X1 U11895 ( .IN1(n7695), .IN2(n7099), .Q(n7694) );
  MUX21X1 U11896 ( .IN1(\mem3[238][31] ), .IN2(n1372), .S(n7696), .Q(n14371)
         );
  MUX21X1 U11897 ( .IN1(\mem3[238][30] ), .IN2(n1350), .S(n7696), .Q(n14370)
         );
  MUX21X1 U11898 ( .IN1(\mem3[238][29] ), .IN2(n1328), .S(n7696), .Q(n14369)
         );
  MUX21X1 U11899 ( .IN1(\mem3[238][28] ), .IN2(n1306), .S(n7696), .Q(n14368)
         );
  MUX21X1 U11900 ( .IN1(\mem3[238][27] ), .IN2(n1284), .S(n7696), .Q(n14367)
         );
  MUX21X1 U11901 ( .IN1(\mem3[238][26] ), .IN2(n1262), .S(n7696), .Q(n14366)
         );
  MUX21X1 U11902 ( .IN1(\mem3[238][25] ), .IN2(n1240), .S(n7696), .Q(n14365)
         );
  MUX21X1 U11903 ( .IN1(\mem3[238][24] ), .IN2(n1218), .S(n7696), .Q(n14364)
         );
  AND2X1 U11904 ( .IN1(n7695), .IN2(n7102), .Q(n7696) );
  MUX21X1 U11905 ( .IN1(\mem3[237][31] ), .IN2(n1372), .S(n7697), .Q(n14363)
         );
  MUX21X1 U11906 ( .IN1(\mem3[237][30] ), .IN2(n1350), .S(n7697), .Q(n14362)
         );
  MUX21X1 U11907 ( .IN1(\mem3[237][29] ), .IN2(n1328), .S(n7697), .Q(n14361)
         );
  MUX21X1 U11908 ( .IN1(\mem3[237][28] ), .IN2(n1306), .S(n7697), .Q(n14360)
         );
  MUX21X1 U11909 ( .IN1(\mem3[237][27] ), .IN2(n1284), .S(n7697), .Q(n14359)
         );
  MUX21X1 U11910 ( .IN1(\mem3[237][26] ), .IN2(n1262), .S(n7697), .Q(n14358)
         );
  MUX21X1 U11911 ( .IN1(\mem3[237][25] ), .IN2(n1240), .S(n7697), .Q(n14357)
         );
  MUX21X1 U11912 ( .IN1(\mem3[237][24] ), .IN2(n1218), .S(n7697), .Q(n14356)
         );
  AND2X1 U11913 ( .IN1(n7695), .IN2(n7104), .Q(n7697) );
  MUX21X1 U11914 ( .IN1(\mem3[236][31] ), .IN2(n1372), .S(n7698), .Q(n14355)
         );
  MUX21X1 U11915 ( .IN1(\mem3[236][30] ), .IN2(n1350), .S(n7698), .Q(n14354)
         );
  MUX21X1 U11916 ( .IN1(\mem3[236][29] ), .IN2(n1328), .S(n7698), .Q(n14353)
         );
  MUX21X1 U11917 ( .IN1(\mem3[236][28] ), .IN2(n1306), .S(n7698), .Q(n14352)
         );
  MUX21X1 U11918 ( .IN1(\mem3[236][27] ), .IN2(n1284), .S(n7698), .Q(n14351)
         );
  MUX21X1 U11919 ( .IN1(\mem3[236][26] ), .IN2(n1262), .S(n7698), .Q(n14350)
         );
  MUX21X1 U11920 ( .IN1(\mem3[236][25] ), .IN2(n1240), .S(n7698), .Q(n14349)
         );
  MUX21X1 U11921 ( .IN1(\mem3[236][24] ), .IN2(n1218), .S(n7698), .Q(n14348)
         );
  AND2X1 U11922 ( .IN1(n7695), .IN2(n7106), .Q(n7698) );
  MUX21X1 U11923 ( .IN1(\mem3[235][31] ), .IN2(n1372), .S(n7699), .Q(n14347)
         );
  MUX21X1 U11924 ( .IN1(\mem3[235][30] ), .IN2(n1350), .S(n7699), .Q(n14346)
         );
  MUX21X1 U11925 ( .IN1(\mem3[235][29] ), .IN2(n1328), .S(n7699), .Q(n14345)
         );
  MUX21X1 U11926 ( .IN1(\mem3[235][28] ), .IN2(n1306), .S(n7699), .Q(n14344)
         );
  MUX21X1 U11927 ( .IN1(\mem3[235][27] ), .IN2(n1284), .S(n7699), .Q(n14343)
         );
  MUX21X1 U11928 ( .IN1(\mem3[235][26] ), .IN2(n1262), .S(n7699), .Q(n14342)
         );
  MUX21X1 U11929 ( .IN1(\mem3[235][25] ), .IN2(n1240), .S(n7699), .Q(n14341)
         );
  MUX21X1 U11930 ( .IN1(\mem3[235][24] ), .IN2(n1218), .S(n7699), .Q(n14340)
         );
  AND2X1 U11931 ( .IN1(n7695), .IN2(n7108), .Q(n7699) );
  MUX21X1 U11932 ( .IN1(\mem3[234][31] ), .IN2(n1372), .S(n7700), .Q(n14339)
         );
  MUX21X1 U11933 ( .IN1(\mem3[234][30] ), .IN2(n1350), .S(n7700), .Q(n14338)
         );
  MUX21X1 U11934 ( .IN1(\mem3[234][29] ), .IN2(n1328), .S(n7700), .Q(n14337)
         );
  MUX21X1 U11935 ( .IN1(\mem3[234][28] ), .IN2(n1306), .S(n7700), .Q(n14336)
         );
  MUX21X1 U11936 ( .IN1(\mem3[234][27] ), .IN2(n1284), .S(n7700), .Q(n14335)
         );
  MUX21X1 U11937 ( .IN1(\mem3[234][26] ), .IN2(n1262), .S(n7700), .Q(n14334)
         );
  MUX21X1 U11938 ( .IN1(\mem3[234][25] ), .IN2(n1240), .S(n7700), .Q(n14333)
         );
  MUX21X1 U11939 ( .IN1(\mem3[234][24] ), .IN2(n1218), .S(n7700), .Q(n14332)
         );
  AND2X1 U11940 ( .IN1(n7695), .IN2(n7110), .Q(n7700) );
  MUX21X1 U11941 ( .IN1(\mem3[233][31] ), .IN2(n1372), .S(n7701), .Q(n14331)
         );
  MUX21X1 U11942 ( .IN1(\mem3[233][30] ), .IN2(n1350), .S(n7701), .Q(n14330)
         );
  MUX21X1 U11943 ( .IN1(\mem3[233][29] ), .IN2(n1328), .S(n7701), .Q(n14329)
         );
  MUX21X1 U11944 ( .IN1(\mem3[233][28] ), .IN2(n1306), .S(n7701), .Q(n14328)
         );
  MUX21X1 U11945 ( .IN1(\mem3[233][27] ), .IN2(n1284), .S(n7701), .Q(n14327)
         );
  MUX21X1 U11946 ( .IN1(\mem3[233][26] ), .IN2(n1262), .S(n7701), .Q(n14326)
         );
  MUX21X1 U11947 ( .IN1(\mem3[233][25] ), .IN2(n1240), .S(n7701), .Q(n14325)
         );
  MUX21X1 U11948 ( .IN1(\mem3[233][24] ), .IN2(n1218), .S(n7701), .Q(n14324)
         );
  AND2X1 U11949 ( .IN1(n7695), .IN2(n7112), .Q(n7701) );
  MUX21X1 U11950 ( .IN1(\mem3[232][31] ), .IN2(n1372), .S(n7702), .Q(n14323)
         );
  MUX21X1 U11951 ( .IN1(\mem3[232][30] ), .IN2(n1350), .S(n7702), .Q(n14322)
         );
  MUX21X1 U11952 ( .IN1(\mem3[232][29] ), .IN2(n1328), .S(n7702), .Q(n14321)
         );
  MUX21X1 U11953 ( .IN1(\mem3[232][28] ), .IN2(n1306), .S(n7702), .Q(n14320)
         );
  MUX21X1 U11954 ( .IN1(\mem3[232][27] ), .IN2(n1284), .S(n7702), .Q(n14319)
         );
  MUX21X1 U11955 ( .IN1(\mem3[232][26] ), .IN2(n1262), .S(n7702), .Q(n14318)
         );
  MUX21X1 U11956 ( .IN1(\mem3[232][25] ), .IN2(n1240), .S(n7702), .Q(n14317)
         );
  MUX21X1 U11957 ( .IN1(\mem3[232][24] ), .IN2(n1218), .S(n7702), .Q(n14316)
         );
  AND2X1 U11958 ( .IN1(n7695), .IN2(n7114), .Q(n7702) );
  MUX21X1 U11959 ( .IN1(\mem3[231][31] ), .IN2(n1373), .S(n7703), .Q(n14315)
         );
  MUX21X1 U11960 ( .IN1(\mem3[231][30] ), .IN2(n1351), .S(n7703), .Q(n14314)
         );
  MUX21X1 U11961 ( .IN1(\mem3[231][29] ), .IN2(n1329), .S(n7703), .Q(n14313)
         );
  MUX21X1 U11962 ( .IN1(\mem3[231][28] ), .IN2(n1307), .S(n7703), .Q(n14312)
         );
  MUX21X1 U11963 ( .IN1(\mem3[231][27] ), .IN2(n1285), .S(n7703), .Q(n14311)
         );
  MUX21X1 U11964 ( .IN1(\mem3[231][26] ), .IN2(n1263), .S(n7703), .Q(n14310)
         );
  MUX21X1 U11965 ( .IN1(\mem3[231][25] ), .IN2(n1241), .S(n7703), .Q(n14309)
         );
  MUX21X1 U11966 ( .IN1(\mem3[231][24] ), .IN2(n1219), .S(n7703), .Q(n14308)
         );
  AND2X1 U11967 ( .IN1(n7695), .IN2(n7116), .Q(n7703) );
  MUX21X1 U11968 ( .IN1(\mem3[230][31] ), .IN2(n1373), .S(n7704), .Q(n14307)
         );
  MUX21X1 U11969 ( .IN1(\mem3[230][30] ), .IN2(n1351), .S(n7704), .Q(n14306)
         );
  MUX21X1 U11970 ( .IN1(\mem3[230][29] ), .IN2(n1329), .S(n7704), .Q(n14305)
         );
  MUX21X1 U11971 ( .IN1(\mem3[230][28] ), .IN2(n1307), .S(n7704), .Q(n14304)
         );
  MUX21X1 U11972 ( .IN1(\mem3[230][27] ), .IN2(n1285), .S(n7704), .Q(n14303)
         );
  MUX21X1 U11973 ( .IN1(\mem3[230][26] ), .IN2(n1263), .S(n7704), .Q(n14302)
         );
  MUX21X1 U11974 ( .IN1(\mem3[230][25] ), .IN2(n1241), .S(n7704), .Q(n14301)
         );
  MUX21X1 U11975 ( .IN1(\mem3[230][24] ), .IN2(n1219), .S(n7704), .Q(n14300)
         );
  AND2X1 U11976 ( .IN1(n7695), .IN2(n7118), .Q(n7704) );
  MUX21X1 U11977 ( .IN1(\mem3[229][31] ), .IN2(n1373), .S(n7705), .Q(n14299)
         );
  MUX21X1 U11978 ( .IN1(\mem3[229][30] ), .IN2(n1351), .S(n7705), .Q(n14298)
         );
  MUX21X1 U11979 ( .IN1(\mem3[229][29] ), .IN2(n1329), .S(n7705), .Q(n14297)
         );
  MUX21X1 U11980 ( .IN1(\mem3[229][28] ), .IN2(n1307), .S(n7705), .Q(n14296)
         );
  MUX21X1 U11981 ( .IN1(\mem3[229][27] ), .IN2(n1285), .S(n7705), .Q(n14295)
         );
  MUX21X1 U11982 ( .IN1(\mem3[229][26] ), .IN2(n1263), .S(n7705), .Q(n14294)
         );
  MUX21X1 U11983 ( .IN1(\mem3[229][25] ), .IN2(n1241), .S(n7705), .Q(n14293)
         );
  MUX21X1 U11984 ( .IN1(\mem3[229][24] ), .IN2(n1219), .S(n7705), .Q(n14292)
         );
  AND2X1 U11985 ( .IN1(n7695), .IN2(n7120), .Q(n7705) );
  MUX21X1 U11986 ( .IN1(\mem3[228][31] ), .IN2(n1373), .S(n7706), .Q(n14291)
         );
  MUX21X1 U11987 ( .IN1(\mem3[228][30] ), .IN2(n1351), .S(n7706), .Q(n14290)
         );
  MUX21X1 U11988 ( .IN1(\mem3[228][29] ), .IN2(n1329), .S(n7706), .Q(n14289)
         );
  MUX21X1 U11989 ( .IN1(\mem3[228][28] ), .IN2(n1307), .S(n7706), .Q(n14288)
         );
  MUX21X1 U11990 ( .IN1(\mem3[228][27] ), .IN2(n1285), .S(n7706), .Q(n14287)
         );
  MUX21X1 U11991 ( .IN1(\mem3[228][26] ), .IN2(n1263), .S(n7706), .Q(n14286)
         );
  MUX21X1 U11992 ( .IN1(\mem3[228][25] ), .IN2(n1241), .S(n7706), .Q(n14285)
         );
  MUX21X1 U11993 ( .IN1(\mem3[228][24] ), .IN2(n1219), .S(n7706), .Q(n14284)
         );
  AND2X1 U11994 ( .IN1(n7695), .IN2(n7122), .Q(n7706) );
  MUX21X1 U11995 ( .IN1(\mem3[227][31] ), .IN2(n1373), .S(n7707), .Q(n14283)
         );
  MUX21X1 U11996 ( .IN1(\mem3[227][30] ), .IN2(n1351), .S(n7707), .Q(n14282)
         );
  MUX21X1 U11997 ( .IN1(\mem3[227][29] ), .IN2(n1329), .S(n7707), .Q(n14281)
         );
  MUX21X1 U11998 ( .IN1(\mem3[227][28] ), .IN2(n1307), .S(n7707), .Q(n14280)
         );
  MUX21X1 U11999 ( .IN1(\mem3[227][27] ), .IN2(n1285), .S(n7707), .Q(n14279)
         );
  MUX21X1 U12000 ( .IN1(\mem3[227][26] ), .IN2(n1263), .S(n7707), .Q(n14278)
         );
  MUX21X1 U12001 ( .IN1(\mem3[227][25] ), .IN2(n1241), .S(n7707), .Q(n14277)
         );
  MUX21X1 U12002 ( .IN1(\mem3[227][24] ), .IN2(n1219), .S(n7707), .Q(n14276)
         );
  AND2X1 U12003 ( .IN1(n7695), .IN2(n7124), .Q(n7707) );
  MUX21X1 U12004 ( .IN1(\mem3[226][31] ), .IN2(n1373), .S(n7708), .Q(n14275)
         );
  MUX21X1 U12005 ( .IN1(\mem3[226][30] ), .IN2(n1351), .S(n7708), .Q(n14274)
         );
  MUX21X1 U12006 ( .IN1(\mem3[226][29] ), .IN2(n1329), .S(n7708), .Q(n14273)
         );
  MUX21X1 U12007 ( .IN1(\mem3[226][28] ), .IN2(n1307), .S(n7708), .Q(n14272)
         );
  MUX21X1 U12008 ( .IN1(\mem3[226][27] ), .IN2(n1285), .S(n7708), .Q(n14271)
         );
  MUX21X1 U12009 ( .IN1(\mem3[226][26] ), .IN2(n1263), .S(n7708), .Q(n14270)
         );
  MUX21X1 U12010 ( .IN1(\mem3[226][25] ), .IN2(n1241), .S(n7708), .Q(n14269)
         );
  MUX21X1 U12011 ( .IN1(\mem3[226][24] ), .IN2(n1219), .S(n7708), .Q(n14268)
         );
  AND2X1 U12012 ( .IN1(n7695), .IN2(n7126), .Q(n7708) );
  MUX21X1 U12013 ( .IN1(\mem3[225][31] ), .IN2(n1373), .S(n7709), .Q(n14267)
         );
  MUX21X1 U12014 ( .IN1(\mem3[225][30] ), .IN2(n1351), .S(n7709), .Q(n14266)
         );
  MUX21X1 U12015 ( .IN1(\mem3[225][29] ), .IN2(n1329), .S(n7709), .Q(n14265)
         );
  MUX21X1 U12016 ( .IN1(\mem3[225][28] ), .IN2(n1307), .S(n7709), .Q(n14264)
         );
  MUX21X1 U12017 ( .IN1(\mem3[225][27] ), .IN2(n1285), .S(n7709), .Q(n14263)
         );
  MUX21X1 U12018 ( .IN1(\mem3[225][26] ), .IN2(n1263), .S(n7709), .Q(n14262)
         );
  MUX21X1 U12019 ( .IN1(\mem3[225][25] ), .IN2(n1241), .S(n7709), .Q(n14261)
         );
  MUX21X1 U12020 ( .IN1(\mem3[225][24] ), .IN2(n1219), .S(n7709), .Q(n14260)
         );
  AND2X1 U12021 ( .IN1(n7695), .IN2(n7128), .Q(n7709) );
  MUX21X1 U12022 ( .IN1(\mem3[224][31] ), .IN2(n1373), .S(n7710), .Q(n14259)
         );
  MUX21X1 U12023 ( .IN1(\mem3[224][30] ), .IN2(n1351), .S(n7710), .Q(n14258)
         );
  MUX21X1 U12024 ( .IN1(\mem3[224][29] ), .IN2(n1329), .S(n7710), .Q(n14257)
         );
  MUX21X1 U12025 ( .IN1(\mem3[224][28] ), .IN2(n1307), .S(n7710), .Q(n14256)
         );
  MUX21X1 U12026 ( .IN1(\mem3[224][27] ), .IN2(n1285), .S(n7710), .Q(n14255)
         );
  MUX21X1 U12027 ( .IN1(\mem3[224][26] ), .IN2(n1263), .S(n7710), .Q(n14254)
         );
  MUX21X1 U12028 ( .IN1(\mem3[224][25] ), .IN2(n1241), .S(n7710), .Q(n14253)
         );
  MUX21X1 U12029 ( .IN1(\mem3[224][24] ), .IN2(n1219), .S(n7710), .Q(n14252)
         );
  AND2X1 U12030 ( .IN1(n7695), .IN2(n7130), .Q(n7710) );
  AND2X1 U12031 ( .IN1(n7693), .IN2(n7150), .Q(n7695) );
  MUX21X1 U12032 ( .IN1(\mem3[223][31] ), .IN2(n1373), .S(n7711), .Q(n14251)
         );
  MUX21X1 U12033 ( .IN1(\mem3[223][30] ), .IN2(n1351), .S(n7711), .Q(n14250)
         );
  MUX21X1 U12034 ( .IN1(\mem3[223][29] ), .IN2(n1329), .S(n7711), .Q(n14249)
         );
  MUX21X1 U12035 ( .IN1(\mem3[223][28] ), .IN2(n1307), .S(n7711), .Q(n14248)
         );
  MUX21X1 U12036 ( .IN1(\mem3[223][27] ), .IN2(n1285), .S(n7711), .Q(n14247)
         );
  MUX21X1 U12037 ( .IN1(\mem3[223][26] ), .IN2(n1263), .S(n7711), .Q(n14246)
         );
  MUX21X1 U12038 ( .IN1(\mem3[223][25] ), .IN2(n1241), .S(n7711), .Q(n14245)
         );
  MUX21X1 U12039 ( .IN1(\mem3[223][24] ), .IN2(n1219), .S(n7711), .Q(n14244)
         );
  AND2X1 U12040 ( .IN1(n7712), .IN2(n7099), .Q(n7711) );
  MUX21X1 U12041 ( .IN1(\mem3[222][31] ), .IN2(n1373), .S(n7713), .Q(n14243)
         );
  MUX21X1 U12042 ( .IN1(\mem3[222][30] ), .IN2(n1351), .S(n7713), .Q(n14242)
         );
  MUX21X1 U12043 ( .IN1(\mem3[222][29] ), .IN2(n1329), .S(n7713), .Q(n14241)
         );
  MUX21X1 U12044 ( .IN1(\mem3[222][28] ), .IN2(n1307), .S(n7713), .Q(n14240)
         );
  MUX21X1 U12045 ( .IN1(\mem3[222][27] ), .IN2(n1285), .S(n7713), .Q(n14239)
         );
  MUX21X1 U12046 ( .IN1(\mem3[222][26] ), .IN2(n1263), .S(n7713), .Q(n14238)
         );
  MUX21X1 U12047 ( .IN1(\mem3[222][25] ), .IN2(n1241), .S(n7713), .Q(n14237)
         );
  MUX21X1 U12048 ( .IN1(\mem3[222][24] ), .IN2(n1219), .S(n7713), .Q(n14236)
         );
  AND2X1 U12049 ( .IN1(n7712), .IN2(n7102), .Q(n7713) );
  MUX21X1 U12050 ( .IN1(\mem3[221][31] ), .IN2(n1373), .S(n7714), .Q(n14235)
         );
  MUX21X1 U12051 ( .IN1(\mem3[221][30] ), .IN2(n1351), .S(n7714), .Q(n14234)
         );
  MUX21X1 U12052 ( .IN1(\mem3[221][29] ), .IN2(n1329), .S(n7714), .Q(n14233)
         );
  MUX21X1 U12053 ( .IN1(\mem3[221][28] ), .IN2(n1307), .S(n7714), .Q(n14232)
         );
  MUX21X1 U12054 ( .IN1(\mem3[221][27] ), .IN2(n1285), .S(n7714), .Q(n14231)
         );
  MUX21X1 U12055 ( .IN1(\mem3[221][26] ), .IN2(n1263), .S(n7714), .Q(n14230)
         );
  MUX21X1 U12056 ( .IN1(\mem3[221][25] ), .IN2(n1241), .S(n7714), .Q(n14229)
         );
  MUX21X1 U12057 ( .IN1(\mem3[221][24] ), .IN2(n1219), .S(n7714), .Q(n14228)
         );
  AND2X1 U12058 ( .IN1(n7712), .IN2(n7104), .Q(n7714) );
  MUX21X1 U12059 ( .IN1(\mem3[220][31] ), .IN2(n1373), .S(n7715), .Q(n14227)
         );
  MUX21X1 U12060 ( .IN1(\mem3[220][30] ), .IN2(n1351), .S(n7715), .Q(n14226)
         );
  MUX21X1 U12061 ( .IN1(\mem3[220][29] ), .IN2(n1329), .S(n7715), .Q(n14225)
         );
  MUX21X1 U12062 ( .IN1(\mem3[220][28] ), .IN2(n1307), .S(n7715), .Q(n14224)
         );
  MUX21X1 U12063 ( .IN1(\mem3[220][27] ), .IN2(n1285), .S(n7715), .Q(n14223)
         );
  MUX21X1 U12064 ( .IN1(\mem3[220][26] ), .IN2(n1263), .S(n7715), .Q(n14222)
         );
  MUX21X1 U12065 ( .IN1(\mem3[220][25] ), .IN2(n1241), .S(n7715), .Q(n14221)
         );
  MUX21X1 U12066 ( .IN1(\mem3[220][24] ), .IN2(n1219), .S(n7715), .Q(n14220)
         );
  AND2X1 U12067 ( .IN1(n7712), .IN2(n7106), .Q(n7715) );
  MUX21X1 U12068 ( .IN1(\mem3[219][31] ), .IN2(n1374), .S(n7716), .Q(n14219)
         );
  MUX21X1 U12069 ( .IN1(\mem3[219][30] ), .IN2(n1352), .S(n7716), .Q(n14218)
         );
  MUX21X1 U12070 ( .IN1(\mem3[219][29] ), .IN2(n1330), .S(n7716), .Q(n14217)
         );
  MUX21X1 U12071 ( .IN1(\mem3[219][28] ), .IN2(n1308), .S(n7716), .Q(n14216)
         );
  MUX21X1 U12072 ( .IN1(\mem3[219][27] ), .IN2(n1286), .S(n7716), .Q(n14215)
         );
  MUX21X1 U12073 ( .IN1(\mem3[219][26] ), .IN2(n1264), .S(n7716), .Q(n14214)
         );
  MUX21X1 U12074 ( .IN1(\mem3[219][25] ), .IN2(n1242), .S(n7716), .Q(n14213)
         );
  MUX21X1 U12075 ( .IN1(\mem3[219][24] ), .IN2(n1220), .S(n7716), .Q(n14212)
         );
  AND2X1 U12076 ( .IN1(n7712), .IN2(n7108), .Q(n7716) );
  MUX21X1 U12077 ( .IN1(\mem3[218][31] ), .IN2(n1374), .S(n7717), .Q(n14211)
         );
  MUX21X1 U12078 ( .IN1(\mem3[218][30] ), .IN2(n1352), .S(n7717), .Q(n14210)
         );
  MUX21X1 U12079 ( .IN1(\mem3[218][29] ), .IN2(n1330), .S(n7717), .Q(n14209)
         );
  MUX21X1 U12080 ( .IN1(\mem3[218][28] ), .IN2(n1308), .S(n7717), .Q(n14208)
         );
  MUX21X1 U12081 ( .IN1(\mem3[218][27] ), .IN2(n1286), .S(n7717), .Q(n14207)
         );
  MUX21X1 U12082 ( .IN1(\mem3[218][26] ), .IN2(n1264), .S(n7717), .Q(n14206)
         );
  MUX21X1 U12083 ( .IN1(\mem3[218][25] ), .IN2(n1242), .S(n7717), .Q(n14205)
         );
  MUX21X1 U12084 ( .IN1(\mem3[218][24] ), .IN2(n1220), .S(n7717), .Q(n14204)
         );
  AND2X1 U12085 ( .IN1(n7712), .IN2(n7110), .Q(n7717) );
  MUX21X1 U12086 ( .IN1(\mem3[217][31] ), .IN2(n1374), .S(n7718), .Q(n14203)
         );
  MUX21X1 U12087 ( .IN1(\mem3[217][30] ), .IN2(n1352), .S(n7718), .Q(n14202)
         );
  MUX21X1 U12088 ( .IN1(\mem3[217][29] ), .IN2(n1330), .S(n7718), .Q(n14201)
         );
  MUX21X1 U12089 ( .IN1(\mem3[217][28] ), .IN2(n1308), .S(n7718), .Q(n14200)
         );
  MUX21X1 U12090 ( .IN1(\mem3[217][27] ), .IN2(n1286), .S(n7718), .Q(n14199)
         );
  MUX21X1 U12091 ( .IN1(\mem3[217][26] ), .IN2(n1264), .S(n7718), .Q(n14198)
         );
  MUX21X1 U12092 ( .IN1(\mem3[217][25] ), .IN2(n1242), .S(n7718), .Q(n14197)
         );
  MUX21X1 U12093 ( .IN1(\mem3[217][24] ), .IN2(n1220), .S(n7718), .Q(n14196)
         );
  AND2X1 U12094 ( .IN1(n7712), .IN2(n7112), .Q(n7718) );
  MUX21X1 U12095 ( .IN1(\mem3[216][31] ), .IN2(n1374), .S(n7719), .Q(n14195)
         );
  MUX21X1 U12096 ( .IN1(\mem3[216][30] ), .IN2(n1352), .S(n7719), .Q(n14194)
         );
  MUX21X1 U12097 ( .IN1(\mem3[216][29] ), .IN2(n1330), .S(n7719), .Q(n14193)
         );
  MUX21X1 U12098 ( .IN1(\mem3[216][28] ), .IN2(n1308), .S(n7719), .Q(n14192)
         );
  MUX21X1 U12099 ( .IN1(\mem3[216][27] ), .IN2(n1286), .S(n7719), .Q(n14191)
         );
  MUX21X1 U12100 ( .IN1(\mem3[216][26] ), .IN2(n1264), .S(n7719), .Q(n14190)
         );
  MUX21X1 U12101 ( .IN1(\mem3[216][25] ), .IN2(n1242), .S(n7719), .Q(n14189)
         );
  MUX21X1 U12102 ( .IN1(\mem3[216][24] ), .IN2(n1220), .S(n7719), .Q(n14188)
         );
  AND2X1 U12103 ( .IN1(n7712), .IN2(n7114), .Q(n7719) );
  MUX21X1 U12104 ( .IN1(\mem3[215][31] ), .IN2(n1374), .S(n7720), .Q(n14187)
         );
  MUX21X1 U12105 ( .IN1(\mem3[215][30] ), .IN2(n1352), .S(n7720), .Q(n14186)
         );
  MUX21X1 U12106 ( .IN1(\mem3[215][29] ), .IN2(n1330), .S(n7720), .Q(n14185)
         );
  MUX21X1 U12107 ( .IN1(\mem3[215][28] ), .IN2(n1308), .S(n7720), .Q(n14184)
         );
  MUX21X1 U12108 ( .IN1(\mem3[215][27] ), .IN2(n1286), .S(n7720), .Q(n14183)
         );
  MUX21X1 U12109 ( .IN1(\mem3[215][26] ), .IN2(n1264), .S(n7720), .Q(n14182)
         );
  MUX21X1 U12110 ( .IN1(\mem3[215][25] ), .IN2(n1242), .S(n7720), .Q(n14181)
         );
  MUX21X1 U12111 ( .IN1(\mem3[215][24] ), .IN2(n1220), .S(n7720), .Q(n14180)
         );
  AND2X1 U12112 ( .IN1(n7712), .IN2(n7116), .Q(n7720) );
  MUX21X1 U12113 ( .IN1(\mem3[214][31] ), .IN2(n1374), .S(n7721), .Q(n14179)
         );
  MUX21X1 U12114 ( .IN1(\mem3[214][30] ), .IN2(n1352), .S(n7721), .Q(n14178)
         );
  MUX21X1 U12115 ( .IN1(\mem3[214][29] ), .IN2(n1330), .S(n7721), .Q(n14177)
         );
  MUX21X1 U12116 ( .IN1(\mem3[214][28] ), .IN2(n1308), .S(n7721), .Q(n14176)
         );
  MUX21X1 U12117 ( .IN1(\mem3[214][27] ), .IN2(n1286), .S(n7721), .Q(n14175)
         );
  MUX21X1 U12118 ( .IN1(\mem3[214][26] ), .IN2(n1264), .S(n7721), .Q(n14174)
         );
  MUX21X1 U12119 ( .IN1(\mem3[214][25] ), .IN2(n1242), .S(n7721), .Q(n14173)
         );
  MUX21X1 U12120 ( .IN1(\mem3[214][24] ), .IN2(n1220), .S(n7721), .Q(n14172)
         );
  AND2X1 U12121 ( .IN1(n7712), .IN2(n7118), .Q(n7721) );
  MUX21X1 U12122 ( .IN1(\mem3[213][31] ), .IN2(n1374), .S(n7722), .Q(n14171)
         );
  MUX21X1 U12123 ( .IN1(\mem3[213][30] ), .IN2(n1352), .S(n7722), .Q(n14170)
         );
  MUX21X1 U12124 ( .IN1(\mem3[213][29] ), .IN2(n1330), .S(n7722), .Q(n14169)
         );
  MUX21X1 U12125 ( .IN1(\mem3[213][28] ), .IN2(n1308), .S(n7722), .Q(n14168)
         );
  MUX21X1 U12126 ( .IN1(\mem3[213][27] ), .IN2(n1286), .S(n7722), .Q(n14167)
         );
  MUX21X1 U12127 ( .IN1(\mem3[213][26] ), .IN2(n1264), .S(n7722), .Q(n14166)
         );
  MUX21X1 U12128 ( .IN1(\mem3[213][25] ), .IN2(n1242), .S(n7722), .Q(n14165)
         );
  MUX21X1 U12129 ( .IN1(\mem3[213][24] ), .IN2(n1220), .S(n7722), .Q(n14164)
         );
  AND2X1 U12130 ( .IN1(n7712), .IN2(n7120), .Q(n7722) );
  MUX21X1 U12131 ( .IN1(\mem3[212][31] ), .IN2(n1374), .S(n7723), .Q(n14163)
         );
  MUX21X1 U12132 ( .IN1(\mem3[212][30] ), .IN2(n1352), .S(n7723), .Q(n14162)
         );
  MUX21X1 U12133 ( .IN1(\mem3[212][29] ), .IN2(n1330), .S(n7723), .Q(n14161)
         );
  MUX21X1 U12134 ( .IN1(\mem3[212][28] ), .IN2(n1308), .S(n7723), .Q(n14160)
         );
  MUX21X1 U12135 ( .IN1(\mem3[212][27] ), .IN2(n1286), .S(n7723), .Q(n14159)
         );
  MUX21X1 U12136 ( .IN1(\mem3[212][26] ), .IN2(n1264), .S(n7723), .Q(n14158)
         );
  MUX21X1 U12137 ( .IN1(\mem3[212][25] ), .IN2(n1242), .S(n7723), .Q(n14157)
         );
  MUX21X1 U12138 ( .IN1(\mem3[212][24] ), .IN2(n1220), .S(n7723), .Q(n14156)
         );
  AND2X1 U12139 ( .IN1(n7712), .IN2(n7122), .Q(n7723) );
  MUX21X1 U12140 ( .IN1(\mem3[211][31] ), .IN2(n1374), .S(n7724), .Q(n14155)
         );
  MUX21X1 U12141 ( .IN1(\mem3[211][30] ), .IN2(n1352), .S(n7724), .Q(n14154)
         );
  MUX21X1 U12142 ( .IN1(\mem3[211][29] ), .IN2(n1330), .S(n7724), .Q(n14153)
         );
  MUX21X1 U12143 ( .IN1(\mem3[211][28] ), .IN2(n1308), .S(n7724), .Q(n14152)
         );
  MUX21X1 U12144 ( .IN1(\mem3[211][27] ), .IN2(n1286), .S(n7724), .Q(n14151)
         );
  MUX21X1 U12145 ( .IN1(\mem3[211][26] ), .IN2(n1264), .S(n7724), .Q(n14150)
         );
  MUX21X1 U12146 ( .IN1(\mem3[211][25] ), .IN2(n1242), .S(n7724), .Q(n14149)
         );
  MUX21X1 U12147 ( .IN1(\mem3[211][24] ), .IN2(n1220), .S(n7724), .Q(n14148)
         );
  AND2X1 U12148 ( .IN1(n7712), .IN2(n7124), .Q(n7724) );
  MUX21X1 U12149 ( .IN1(\mem3[210][31] ), .IN2(n1374), .S(n7725), .Q(n14147)
         );
  MUX21X1 U12150 ( .IN1(\mem3[210][30] ), .IN2(n1352), .S(n7725), .Q(n14146)
         );
  MUX21X1 U12151 ( .IN1(\mem3[210][29] ), .IN2(n1330), .S(n7725), .Q(n14145)
         );
  MUX21X1 U12152 ( .IN1(\mem3[210][28] ), .IN2(n1308), .S(n7725), .Q(n14144)
         );
  MUX21X1 U12153 ( .IN1(\mem3[210][27] ), .IN2(n1286), .S(n7725), .Q(n14143)
         );
  MUX21X1 U12154 ( .IN1(\mem3[210][26] ), .IN2(n1264), .S(n7725), .Q(n14142)
         );
  MUX21X1 U12155 ( .IN1(\mem3[210][25] ), .IN2(n1242), .S(n7725), .Q(n14141)
         );
  MUX21X1 U12156 ( .IN1(\mem3[210][24] ), .IN2(n1220), .S(n7725), .Q(n14140)
         );
  AND2X1 U12157 ( .IN1(n7712), .IN2(n7126), .Q(n7725) );
  MUX21X1 U12158 ( .IN1(\mem3[209][31] ), .IN2(n1374), .S(n7726), .Q(n14139)
         );
  MUX21X1 U12159 ( .IN1(\mem3[209][30] ), .IN2(n1352), .S(n7726), .Q(n14138)
         );
  MUX21X1 U12160 ( .IN1(\mem3[209][29] ), .IN2(n1330), .S(n7726), .Q(n14137)
         );
  MUX21X1 U12161 ( .IN1(\mem3[209][28] ), .IN2(n1308), .S(n7726), .Q(n14136)
         );
  MUX21X1 U12162 ( .IN1(\mem3[209][27] ), .IN2(n1286), .S(n7726), .Q(n14135)
         );
  MUX21X1 U12163 ( .IN1(\mem3[209][26] ), .IN2(n1264), .S(n7726), .Q(n14134)
         );
  MUX21X1 U12164 ( .IN1(\mem3[209][25] ), .IN2(n1242), .S(n7726), .Q(n14133)
         );
  MUX21X1 U12165 ( .IN1(\mem3[209][24] ), .IN2(n1220), .S(n7726), .Q(n14132)
         );
  AND2X1 U12166 ( .IN1(n7712), .IN2(n7128), .Q(n7726) );
  MUX21X1 U12167 ( .IN1(\mem3[208][31] ), .IN2(n1374), .S(n7727), .Q(n14131)
         );
  MUX21X1 U12168 ( .IN1(\mem3[208][30] ), .IN2(n1352), .S(n7727), .Q(n14130)
         );
  MUX21X1 U12169 ( .IN1(\mem3[208][29] ), .IN2(n1330), .S(n7727), .Q(n14129)
         );
  MUX21X1 U12170 ( .IN1(\mem3[208][28] ), .IN2(n1308), .S(n7727), .Q(n14128)
         );
  MUX21X1 U12171 ( .IN1(\mem3[208][27] ), .IN2(n1286), .S(n7727), .Q(n14127)
         );
  MUX21X1 U12172 ( .IN1(\mem3[208][26] ), .IN2(n1264), .S(n7727), .Q(n14126)
         );
  MUX21X1 U12173 ( .IN1(\mem3[208][25] ), .IN2(n1242), .S(n7727), .Q(n14125)
         );
  MUX21X1 U12174 ( .IN1(\mem3[208][24] ), .IN2(n1220), .S(n7727), .Q(n14124)
         );
  AND2X1 U12175 ( .IN1(n7712), .IN2(n7130), .Q(n7727) );
  AND2X1 U12176 ( .IN1(n7693), .IN2(n7168), .Q(n7712) );
  MUX21X1 U12177 ( .IN1(\mem3[207][31] ), .IN2(n1375), .S(n7728), .Q(n14123)
         );
  MUX21X1 U12178 ( .IN1(\mem3[207][30] ), .IN2(n1353), .S(n7728), .Q(n14122)
         );
  MUX21X1 U12179 ( .IN1(\mem3[207][29] ), .IN2(n1331), .S(n7728), .Q(n14121)
         );
  MUX21X1 U12180 ( .IN1(\mem3[207][28] ), .IN2(n1309), .S(n7728), .Q(n14120)
         );
  MUX21X1 U12181 ( .IN1(\mem3[207][27] ), .IN2(n1287), .S(n7728), .Q(n14119)
         );
  MUX21X1 U12182 ( .IN1(\mem3[207][26] ), .IN2(n1265), .S(n7728), .Q(n14118)
         );
  MUX21X1 U12183 ( .IN1(\mem3[207][25] ), .IN2(n1243), .S(n7728), .Q(n14117)
         );
  MUX21X1 U12184 ( .IN1(\mem3[207][24] ), .IN2(n1221), .S(n7728), .Q(n14116)
         );
  AND2X1 U12185 ( .IN1(n7729), .IN2(n7099), .Q(n7728) );
  MUX21X1 U12186 ( .IN1(\mem3[206][31] ), .IN2(n1375), .S(n7730), .Q(n14115)
         );
  MUX21X1 U12187 ( .IN1(\mem3[206][30] ), .IN2(n1353), .S(n7730), .Q(n14114)
         );
  MUX21X1 U12188 ( .IN1(\mem3[206][29] ), .IN2(n1331), .S(n7730), .Q(n14113)
         );
  MUX21X1 U12189 ( .IN1(\mem3[206][28] ), .IN2(n1309), .S(n7730), .Q(n14112)
         );
  MUX21X1 U12190 ( .IN1(\mem3[206][27] ), .IN2(n1287), .S(n7730), .Q(n14111)
         );
  MUX21X1 U12191 ( .IN1(\mem3[206][26] ), .IN2(n1265), .S(n7730), .Q(n14110)
         );
  MUX21X1 U12192 ( .IN1(\mem3[206][25] ), .IN2(n1243), .S(n7730), .Q(n14109)
         );
  MUX21X1 U12193 ( .IN1(\mem3[206][24] ), .IN2(n1221), .S(n7730), .Q(n14108)
         );
  AND2X1 U12194 ( .IN1(n7729), .IN2(n7102), .Q(n7730) );
  MUX21X1 U12195 ( .IN1(\mem3[205][31] ), .IN2(n1375), .S(n7731), .Q(n14107)
         );
  MUX21X1 U12196 ( .IN1(\mem3[205][30] ), .IN2(n1353), .S(n7731), .Q(n14106)
         );
  MUX21X1 U12197 ( .IN1(\mem3[205][29] ), .IN2(n1331), .S(n7731), .Q(n14105)
         );
  MUX21X1 U12198 ( .IN1(\mem3[205][28] ), .IN2(n1309), .S(n7731), .Q(n14104)
         );
  MUX21X1 U12199 ( .IN1(\mem3[205][27] ), .IN2(n1287), .S(n7731), .Q(n14103)
         );
  MUX21X1 U12200 ( .IN1(\mem3[205][26] ), .IN2(n1265), .S(n7731), .Q(n14102)
         );
  MUX21X1 U12201 ( .IN1(\mem3[205][25] ), .IN2(n1243), .S(n7731), .Q(n14101)
         );
  MUX21X1 U12202 ( .IN1(\mem3[205][24] ), .IN2(n1221), .S(n7731), .Q(n14100)
         );
  AND2X1 U12203 ( .IN1(n7729), .IN2(n7104), .Q(n7731) );
  MUX21X1 U12204 ( .IN1(\mem3[204][31] ), .IN2(n1375), .S(n7732), .Q(n14099)
         );
  MUX21X1 U12205 ( .IN1(\mem3[204][30] ), .IN2(n1353), .S(n7732), .Q(n14098)
         );
  MUX21X1 U12206 ( .IN1(\mem3[204][29] ), .IN2(n1331), .S(n7732), .Q(n14097)
         );
  MUX21X1 U12207 ( .IN1(\mem3[204][28] ), .IN2(n1309), .S(n7732), .Q(n14096)
         );
  MUX21X1 U12208 ( .IN1(\mem3[204][27] ), .IN2(n1287), .S(n7732), .Q(n14095)
         );
  MUX21X1 U12209 ( .IN1(\mem3[204][26] ), .IN2(n1265), .S(n7732), .Q(n14094)
         );
  MUX21X1 U12210 ( .IN1(\mem3[204][25] ), .IN2(n1243), .S(n7732), .Q(n14093)
         );
  MUX21X1 U12211 ( .IN1(\mem3[204][24] ), .IN2(n1221), .S(n7732), .Q(n14092)
         );
  AND2X1 U12212 ( .IN1(n7729), .IN2(n7106), .Q(n7732) );
  MUX21X1 U12213 ( .IN1(\mem3[203][31] ), .IN2(n1375), .S(n7733), .Q(n14091)
         );
  MUX21X1 U12214 ( .IN1(\mem3[203][30] ), .IN2(n1353), .S(n7733), .Q(n14090)
         );
  MUX21X1 U12215 ( .IN1(\mem3[203][29] ), .IN2(n1331), .S(n7733), .Q(n14089)
         );
  MUX21X1 U12216 ( .IN1(\mem3[203][28] ), .IN2(n1309), .S(n7733), .Q(n14088)
         );
  MUX21X1 U12217 ( .IN1(\mem3[203][27] ), .IN2(n1287), .S(n7733), .Q(n14087)
         );
  MUX21X1 U12218 ( .IN1(\mem3[203][26] ), .IN2(n1265), .S(n7733), .Q(n14086)
         );
  MUX21X1 U12219 ( .IN1(\mem3[203][25] ), .IN2(n1243), .S(n7733), .Q(n14085)
         );
  MUX21X1 U12220 ( .IN1(\mem3[203][24] ), .IN2(n1221), .S(n7733), .Q(n14084)
         );
  AND2X1 U12221 ( .IN1(n7729), .IN2(n7108), .Q(n7733) );
  MUX21X1 U12222 ( .IN1(\mem3[202][31] ), .IN2(n1375), .S(n7734), .Q(n14083)
         );
  MUX21X1 U12223 ( .IN1(\mem3[202][30] ), .IN2(n1353), .S(n7734), .Q(n14082)
         );
  MUX21X1 U12224 ( .IN1(\mem3[202][29] ), .IN2(n1331), .S(n7734), .Q(n14081)
         );
  MUX21X1 U12225 ( .IN1(\mem3[202][28] ), .IN2(n1309), .S(n7734), .Q(n14080)
         );
  MUX21X1 U12226 ( .IN1(\mem3[202][27] ), .IN2(n1287), .S(n7734), .Q(n14079)
         );
  MUX21X1 U12227 ( .IN1(\mem3[202][26] ), .IN2(n1265), .S(n7734), .Q(n14078)
         );
  MUX21X1 U12228 ( .IN1(\mem3[202][25] ), .IN2(n1243), .S(n7734), .Q(n14077)
         );
  MUX21X1 U12229 ( .IN1(\mem3[202][24] ), .IN2(n1221), .S(n7734), .Q(n14076)
         );
  AND2X1 U12230 ( .IN1(n7729), .IN2(n7110), .Q(n7734) );
  MUX21X1 U12231 ( .IN1(\mem3[201][31] ), .IN2(n1375), .S(n7735), .Q(n14075)
         );
  MUX21X1 U12232 ( .IN1(\mem3[201][30] ), .IN2(n1353), .S(n7735), .Q(n14074)
         );
  MUX21X1 U12233 ( .IN1(\mem3[201][29] ), .IN2(n1331), .S(n7735), .Q(n14073)
         );
  MUX21X1 U12234 ( .IN1(\mem3[201][28] ), .IN2(n1309), .S(n7735), .Q(n14072)
         );
  MUX21X1 U12235 ( .IN1(\mem3[201][27] ), .IN2(n1287), .S(n7735), .Q(n14071)
         );
  MUX21X1 U12236 ( .IN1(\mem3[201][26] ), .IN2(n1265), .S(n7735), .Q(n14070)
         );
  MUX21X1 U12237 ( .IN1(\mem3[201][25] ), .IN2(n1243), .S(n7735), .Q(n14069)
         );
  MUX21X1 U12238 ( .IN1(\mem3[201][24] ), .IN2(n1221), .S(n7735), .Q(n14068)
         );
  AND2X1 U12239 ( .IN1(n7729), .IN2(n7112), .Q(n7735) );
  MUX21X1 U12240 ( .IN1(\mem3[200][31] ), .IN2(n1375), .S(n7736), .Q(n14067)
         );
  MUX21X1 U12241 ( .IN1(\mem3[200][30] ), .IN2(n1353), .S(n7736), .Q(n14066)
         );
  MUX21X1 U12242 ( .IN1(\mem3[200][29] ), .IN2(n1331), .S(n7736), .Q(n14065)
         );
  MUX21X1 U12243 ( .IN1(\mem3[200][28] ), .IN2(n1309), .S(n7736), .Q(n14064)
         );
  MUX21X1 U12244 ( .IN1(\mem3[200][27] ), .IN2(n1287), .S(n7736), .Q(n14063)
         );
  MUX21X1 U12245 ( .IN1(\mem3[200][26] ), .IN2(n1265), .S(n7736), .Q(n14062)
         );
  MUX21X1 U12246 ( .IN1(\mem3[200][25] ), .IN2(n1243), .S(n7736), .Q(n14061)
         );
  MUX21X1 U12247 ( .IN1(\mem3[200][24] ), .IN2(n1221), .S(n7736), .Q(n14060)
         );
  AND2X1 U12248 ( .IN1(n7729), .IN2(n7114), .Q(n7736) );
  MUX21X1 U12249 ( .IN1(\mem3[199][31] ), .IN2(n1375), .S(n7737), .Q(n14059)
         );
  MUX21X1 U12250 ( .IN1(\mem3[199][30] ), .IN2(n1353), .S(n7737), .Q(n14058)
         );
  MUX21X1 U12251 ( .IN1(\mem3[199][29] ), .IN2(n1331), .S(n7737), .Q(n14057)
         );
  MUX21X1 U12252 ( .IN1(\mem3[199][28] ), .IN2(n1309), .S(n7737), .Q(n14056)
         );
  MUX21X1 U12253 ( .IN1(\mem3[199][27] ), .IN2(n1287), .S(n7737), .Q(n14055)
         );
  MUX21X1 U12254 ( .IN1(\mem3[199][26] ), .IN2(n1265), .S(n7737), .Q(n14054)
         );
  MUX21X1 U12255 ( .IN1(\mem3[199][25] ), .IN2(n1243), .S(n7737), .Q(n14053)
         );
  MUX21X1 U12256 ( .IN1(\mem3[199][24] ), .IN2(n1221), .S(n7737), .Q(n14052)
         );
  AND2X1 U12257 ( .IN1(n7729), .IN2(n7116), .Q(n7737) );
  MUX21X1 U12258 ( .IN1(\mem3[198][31] ), .IN2(n1375), .S(n7738), .Q(n14051)
         );
  MUX21X1 U12259 ( .IN1(\mem3[198][30] ), .IN2(n1353), .S(n7738), .Q(n14050)
         );
  MUX21X1 U12260 ( .IN1(\mem3[198][29] ), .IN2(n1331), .S(n7738), .Q(n14049)
         );
  MUX21X1 U12261 ( .IN1(\mem3[198][28] ), .IN2(n1309), .S(n7738), .Q(n14048)
         );
  MUX21X1 U12262 ( .IN1(\mem3[198][27] ), .IN2(n1287), .S(n7738), .Q(n14047)
         );
  MUX21X1 U12263 ( .IN1(\mem3[198][26] ), .IN2(n1265), .S(n7738), .Q(n14046)
         );
  MUX21X1 U12264 ( .IN1(\mem3[198][25] ), .IN2(n1243), .S(n7738), .Q(n14045)
         );
  MUX21X1 U12265 ( .IN1(\mem3[198][24] ), .IN2(n1221), .S(n7738), .Q(n14044)
         );
  AND2X1 U12266 ( .IN1(n7729), .IN2(n7118), .Q(n7738) );
  MUX21X1 U12267 ( .IN1(\mem3[197][31] ), .IN2(n1375), .S(n7739), .Q(n14043)
         );
  MUX21X1 U12268 ( .IN1(\mem3[197][30] ), .IN2(n1353), .S(n7739), .Q(n14042)
         );
  MUX21X1 U12269 ( .IN1(\mem3[197][29] ), .IN2(n1331), .S(n7739), .Q(n14041)
         );
  MUX21X1 U12270 ( .IN1(\mem3[197][28] ), .IN2(n1309), .S(n7739), .Q(n14040)
         );
  MUX21X1 U12271 ( .IN1(\mem3[197][27] ), .IN2(n1287), .S(n7739), .Q(n14039)
         );
  MUX21X1 U12272 ( .IN1(\mem3[197][26] ), .IN2(n1265), .S(n7739), .Q(n14038)
         );
  MUX21X1 U12273 ( .IN1(\mem3[197][25] ), .IN2(n1243), .S(n7739), .Q(n14037)
         );
  MUX21X1 U12274 ( .IN1(\mem3[197][24] ), .IN2(n1221), .S(n7739), .Q(n14036)
         );
  AND2X1 U12275 ( .IN1(n7729), .IN2(n7120), .Q(n7739) );
  MUX21X1 U12276 ( .IN1(\mem3[196][31] ), .IN2(n1375), .S(n7740), .Q(n14035)
         );
  MUX21X1 U12277 ( .IN1(\mem3[196][30] ), .IN2(n1353), .S(n7740), .Q(n14034)
         );
  MUX21X1 U12278 ( .IN1(\mem3[196][29] ), .IN2(n1331), .S(n7740), .Q(n14033)
         );
  MUX21X1 U12279 ( .IN1(\mem3[196][28] ), .IN2(n1309), .S(n7740), .Q(n14032)
         );
  MUX21X1 U12280 ( .IN1(\mem3[196][27] ), .IN2(n1287), .S(n7740), .Q(n14031)
         );
  MUX21X1 U12281 ( .IN1(\mem3[196][26] ), .IN2(n1265), .S(n7740), .Q(n14030)
         );
  MUX21X1 U12282 ( .IN1(\mem3[196][25] ), .IN2(n1243), .S(n7740), .Q(n14029)
         );
  MUX21X1 U12283 ( .IN1(\mem3[196][24] ), .IN2(n1221), .S(n7740), .Q(n14028)
         );
  AND2X1 U12284 ( .IN1(n7729), .IN2(n7122), .Q(n7740) );
  MUX21X1 U12285 ( .IN1(\mem3[195][31] ), .IN2(n1376), .S(n7741), .Q(n14027)
         );
  MUX21X1 U12286 ( .IN1(\mem3[195][30] ), .IN2(n1354), .S(n7741), .Q(n14026)
         );
  MUX21X1 U12287 ( .IN1(\mem3[195][29] ), .IN2(n1332), .S(n7741), .Q(n14025)
         );
  MUX21X1 U12288 ( .IN1(\mem3[195][28] ), .IN2(n1310), .S(n7741), .Q(n14024)
         );
  MUX21X1 U12289 ( .IN1(\mem3[195][27] ), .IN2(n1288), .S(n7741), .Q(n14023)
         );
  MUX21X1 U12290 ( .IN1(\mem3[195][26] ), .IN2(n1266), .S(n7741), .Q(n14022)
         );
  MUX21X1 U12291 ( .IN1(\mem3[195][25] ), .IN2(n1244), .S(n7741), .Q(n14021)
         );
  MUX21X1 U12292 ( .IN1(\mem3[195][24] ), .IN2(n1222), .S(n7741), .Q(n14020)
         );
  AND2X1 U12293 ( .IN1(n7729), .IN2(n7124), .Q(n7741) );
  MUX21X1 U12294 ( .IN1(\mem3[194][31] ), .IN2(n1376), .S(n7742), .Q(n14019)
         );
  MUX21X1 U12295 ( .IN1(\mem3[194][30] ), .IN2(n1354), .S(n7742), .Q(n14018)
         );
  MUX21X1 U12296 ( .IN1(\mem3[194][29] ), .IN2(n1332), .S(n7742), .Q(n14017)
         );
  MUX21X1 U12297 ( .IN1(\mem3[194][28] ), .IN2(n1310), .S(n7742), .Q(n14016)
         );
  MUX21X1 U12298 ( .IN1(\mem3[194][27] ), .IN2(n1288), .S(n7742), .Q(n14015)
         );
  MUX21X1 U12299 ( .IN1(\mem3[194][26] ), .IN2(n1266), .S(n7742), .Q(n14014)
         );
  MUX21X1 U12300 ( .IN1(\mem3[194][25] ), .IN2(n1244), .S(n7742), .Q(n14013)
         );
  MUX21X1 U12301 ( .IN1(\mem3[194][24] ), .IN2(n1222), .S(n7742), .Q(n14012)
         );
  AND2X1 U12302 ( .IN1(n7729), .IN2(n7126), .Q(n7742) );
  MUX21X1 U12303 ( .IN1(\mem3[193][31] ), .IN2(n1376), .S(n7743), .Q(n14011)
         );
  MUX21X1 U12304 ( .IN1(\mem3[193][30] ), .IN2(n1354), .S(n7743), .Q(n14010)
         );
  MUX21X1 U12305 ( .IN1(\mem3[193][29] ), .IN2(n1332), .S(n7743), .Q(n14009)
         );
  MUX21X1 U12306 ( .IN1(\mem3[193][28] ), .IN2(n1310), .S(n7743), .Q(n14008)
         );
  MUX21X1 U12307 ( .IN1(\mem3[193][27] ), .IN2(n1288), .S(n7743), .Q(n14007)
         );
  MUX21X1 U12308 ( .IN1(\mem3[193][26] ), .IN2(n1266), .S(n7743), .Q(n14006)
         );
  MUX21X1 U12309 ( .IN1(\mem3[193][25] ), .IN2(n1244), .S(n7743), .Q(n14005)
         );
  MUX21X1 U12310 ( .IN1(\mem3[193][24] ), .IN2(n1222), .S(n7743), .Q(n14004)
         );
  AND2X1 U12311 ( .IN1(n7729), .IN2(n7128), .Q(n7743) );
  MUX21X1 U12312 ( .IN1(\mem3[192][31] ), .IN2(n1376), .S(n7744), .Q(n14003)
         );
  MUX21X1 U12313 ( .IN1(\mem3[192][30] ), .IN2(n1354), .S(n7744), .Q(n14002)
         );
  MUX21X1 U12314 ( .IN1(\mem3[192][29] ), .IN2(n1332), .S(n7744), .Q(n14001)
         );
  MUX21X1 U12315 ( .IN1(\mem3[192][28] ), .IN2(n1310), .S(n7744), .Q(n14000)
         );
  MUX21X1 U12316 ( .IN1(\mem3[192][27] ), .IN2(n1288), .S(n7744), .Q(n13999)
         );
  MUX21X1 U12317 ( .IN1(\mem3[192][26] ), .IN2(n1266), .S(n7744), .Q(n13998)
         );
  MUX21X1 U12318 ( .IN1(\mem3[192][25] ), .IN2(n1244), .S(n7744), .Q(n13997)
         );
  MUX21X1 U12319 ( .IN1(\mem3[192][24] ), .IN2(n1222), .S(n7744), .Q(n13996)
         );
  AND2X1 U12320 ( .IN1(n7729), .IN2(n7130), .Q(n7744) );
  AND2X1 U12321 ( .IN1(n7693), .IN2(n7186), .Q(n7729) );
  MUX21X1 U12322 ( .IN1(\mem3[191][31] ), .IN2(n1376), .S(n7745), .Q(n13995)
         );
  MUX21X1 U12323 ( .IN1(\mem3[191][30] ), .IN2(n1354), .S(n7745), .Q(n13994)
         );
  MUX21X1 U12324 ( .IN1(\mem3[191][29] ), .IN2(n1332), .S(n7745), .Q(n13993)
         );
  MUX21X1 U12325 ( .IN1(\mem3[191][28] ), .IN2(n1310), .S(n7745), .Q(n13992)
         );
  MUX21X1 U12326 ( .IN1(\mem3[191][27] ), .IN2(n1288), .S(n7745), .Q(n13991)
         );
  MUX21X1 U12327 ( .IN1(\mem3[191][26] ), .IN2(n1266), .S(n7745), .Q(n13990)
         );
  MUX21X1 U12328 ( .IN1(\mem3[191][25] ), .IN2(n1244), .S(n7745), .Q(n13989)
         );
  MUX21X1 U12329 ( .IN1(\mem3[191][24] ), .IN2(n1222), .S(n7745), .Q(n13988)
         );
  AND2X1 U12330 ( .IN1(n7746), .IN2(n7099), .Q(n7745) );
  MUX21X1 U12331 ( .IN1(\mem3[190][31] ), .IN2(n1376), .S(n7747), .Q(n13987)
         );
  MUX21X1 U12332 ( .IN1(\mem3[190][30] ), .IN2(n1354), .S(n7747), .Q(n13986)
         );
  MUX21X1 U12333 ( .IN1(\mem3[190][29] ), .IN2(n1332), .S(n7747), .Q(n13985)
         );
  MUX21X1 U12334 ( .IN1(\mem3[190][28] ), .IN2(n1310), .S(n7747), .Q(n13984)
         );
  MUX21X1 U12335 ( .IN1(\mem3[190][27] ), .IN2(n1288), .S(n7747), .Q(n13983)
         );
  MUX21X1 U12336 ( .IN1(\mem3[190][26] ), .IN2(n1266), .S(n7747), .Q(n13982)
         );
  MUX21X1 U12337 ( .IN1(\mem3[190][25] ), .IN2(n1244), .S(n7747), .Q(n13981)
         );
  MUX21X1 U12338 ( .IN1(\mem3[190][24] ), .IN2(n1222), .S(n7747), .Q(n13980)
         );
  AND2X1 U12339 ( .IN1(n7746), .IN2(n7102), .Q(n7747) );
  MUX21X1 U12340 ( .IN1(\mem3[189][31] ), .IN2(n1376), .S(n7748), .Q(n13979)
         );
  MUX21X1 U12341 ( .IN1(\mem3[189][30] ), .IN2(n1354), .S(n7748), .Q(n13978)
         );
  MUX21X1 U12342 ( .IN1(\mem3[189][29] ), .IN2(n1332), .S(n7748), .Q(n13977)
         );
  MUX21X1 U12343 ( .IN1(\mem3[189][28] ), .IN2(n1310), .S(n7748), .Q(n13976)
         );
  MUX21X1 U12344 ( .IN1(\mem3[189][27] ), .IN2(n1288), .S(n7748), .Q(n13975)
         );
  MUX21X1 U12345 ( .IN1(\mem3[189][26] ), .IN2(n1266), .S(n7748), .Q(n13974)
         );
  MUX21X1 U12346 ( .IN1(\mem3[189][25] ), .IN2(n1244), .S(n7748), .Q(n13973)
         );
  MUX21X1 U12347 ( .IN1(\mem3[189][24] ), .IN2(n1222), .S(n7748), .Q(n13972)
         );
  AND2X1 U12348 ( .IN1(n7746), .IN2(n7104), .Q(n7748) );
  MUX21X1 U12349 ( .IN1(\mem3[188][31] ), .IN2(n1376), .S(n7749), .Q(n13971)
         );
  MUX21X1 U12350 ( .IN1(\mem3[188][30] ), .IN2(n1354), .S(n7749), .Q(n13970)
         );
  MUX21X1 U12351 ( .IN1(\mem3[188][29] ), .IN2(n1332), .S(n7749), .Q(n13969)
         );
  MUX21X1 U12352 ( .IN1(\mem3[188][28] ), .IN2(n1310), .S(n7749), .Q(n13968)
         );
  MUX21X1 U12353 ( .IN1(\mem3[188][27] ), .IN2(n1288), .S(n7749), .Q(n13967)
         );
  MUX21X1 U12354 ( .IN1(\mem3[188][26] ), .IN2(n1266), .S(n7749), .Q(n13966)
         );
  MUX21X1 U12355 ( .IN1(\mem3[188][25] ), .IN2(n1244), .S(n7749), .Q(n13965)
         );
  MUX21X1 U12356 ( .IN1(\mem3[188][24] ), .IN2(n1222), .S(n7749), .Q(n13964)
         );
  AND2X1 U12357 ( .IN1(n7746), .IN2(n7106), .Q(n7749) );
  MUX21X1 U12358 ( .IN1(\mem3[187][31] ), .IN2(n1376), .S(n7750), .Q(n13963)
         );
  MUX21X1 U12359 ( .IN1(\mem3[187][30] ), .IN2(n1354), .S(n7750), .Q(n13962)
         );
  MUX21X1 U12360 ( .IN1(\mem3[187][29] ), .IN2(n1332), .S(n7750), .Q(n13961)
         );
  MUX21X1 U12361 ( .IN1(\mem3[187][28] ), .IN2(n1310), .S(n7750), .Q(n13960)
         );
  MUX21X1 U12362 ( .IN1(\mem3[187][27] ), .IN2(n1288), .S(n7750), .Q(n13959)
         );
  MUX21X1 U12363 ( .IN1(\mem3[187][26] ), .IN2(n1266), .S(n7750), .Q(n13958)
         );
  MUX21X1 U12364 ( .IN1(\mem3[187][25] ), .IN2(n1244), .S(n7750), .Q(n13957)
         );
  MUX21X1 U12365 ( .IN1(\mem3[187][24] ), .IN2(n1222), .S(n7750), .Q(n13956)
         );
  AND2X1 U12366 ( .IN1(n7746), .IN2(n7108), .Q(n7750) );
  MUX21X1 U12367 ( .IN1(\mem3[186][31] ), .IN2(n1376), .S(n7751), .Q(n13955)
         );
  MUX21X1 U12368 ( .IN1(\mem3[186][30] ), .IN2(n1354), .S(n7751), .Q(n13954)
         );
  MUX21X1 U12369 ( .IN1(\mem3[186][29] ), .IN2(n1332), .S(n7751), .Q(n13953)
         );
  MUX21X1 U12370 ( .IN1(\mem3[186][28] ), .IN2(n1310), .S(n7751), .Q(n13952)
         );
  MUX21X1 U12371 ( .IN1(\mem3[186][27] ), .IN2(n1288), .S(n7751), .Q(n13951)
         );
  MUX21X1 U12372 ( .IN1(\mem3[186][26] ), .IN2(n1266), .S(n7751), .Q(n13950)
         );
  MUX21X1 U12373 ( .IN1(\mem3[186][25] ), .IN2(n1244), .S(n7751), .Q(n13949)
         );
  MUX21X1 U12374 ( .IN1(\mem3[186][24] ), .IN2(n1222), .S(n7751), .Q(n13948)
         );
  AND2X1 U12375 ( .IN1(n7746), .IN2(n7110), .Q(n7751) );
  MUX21X1 U12376 ( .IN1(\mem3[185][31] ), .IN2(n1376), .S(n7752), .Q(n13947)
         );
  MUX21X1 U12377 ( .IN1(\mem3[185][30] ), .IN2(n1354), .S(n7752), .Q(n13946)
         );
  MUX21X1 U12378 ( .IN1(\mem3[185][29] ), .IN2(n1332), .S(n7752), .Q(n13945)
         );
  MUX21X1 U12379 ( .IN1(\mem3[185][28] ), .IN2(n1310), .S(n7752), .Q(n13944)
         );
  MUX21X1 U12380 ( .IN1(\mem3[185][27] ), .IN2(n1288), .S(n7752), .Q(n13943)
         );
  MUX21X1 U12381 ( .IN1(\mem3[185][26] ), .IN2(n1266), .S(n7752), .Q(n13942)
         );
  MUX21X1 U12382 ( .IN1(\mem3[185][25] ), .IN2(n1244), .S(n7752), .Q(n13941)
         );
  MUX21X1 U12383 ( .IN1(\mem3[185][24] ), .IN2(n1222), .S(n7752), .Q(n13940)
         );
  AND2X1 U12384 ( .IN1(n7746), .IN2(n7112), .Q(n7752) );
  MUX21X1 U12385 ( .IN1(\mem3[184][31] ), .IN2(n1376), .S(n7753), .Q(n13939)
         );
  MUX21X1 U12386 ( .IN1(\mem3[184][30] ), .IN2(n1354), .S(n7753), .Q(n13938)
         );
  MUX21X1 U12387 ( .IN1(\mem3[184][29] ), .IN2(n1332), .S(n7753), .Q(n13937)
         );
  MUX21X1 U12388 ( .IN1(\mem3[184][28] ), .IN2(n1310), .S(n7753), .Q(n13936)
         );
  MUX21X1 U12389 ( .IN1(\mem3[184][27] ), .IN2(n1288), .S(n7753), .Q(n13935)
         );
  MUX21X1 U12390 ( .IN1(\mem3[184][26] ), .IN2(n1266), .S(n7753), .Q(n13934)
         );
  MUX21X1 U12391 ( .IN1(\mem3[184][25] ), .IN2(n1244), .S(n7753), .Q(n13933)
         );
  MUX21X1 U12392 ( .IN1(\mem3[184][24] ), .IN2(n1222), .S(n7753), .Q(n13932)
         );
  AND2X1 U12393 ( .IN1(n7746), .IN2(n7114), .Q(n7753) );
  MUX21X1 U12394 ( .IN1(\mem3[183][31] ), .IN2(n1377), .S(n7754), .Q(n13931)
         );
  MUX21X1 U12395 ( .IN1(\mem3[183][30] ), .IN2(n1355), .S(n7754), .Q(n13930)
         );
  MUX21X1 U12396 ( .IN1(\mem3[183][29] ), .IN2(n1333), .S(n7754), .Q(n13929)
         );
  MUX21X1 U12397 ( .IN1(\mem3[183][28] ), .IN2(n1311), .S(n7754), .Q(n13928)
         );
  MUX21X1 U12398 ( .IN1(\mem3[183][27] ), .IN2(n1289), .S(n7754), .Q(n13927)
         );
  MUX21X1 U12399 ( .IN1(\mem3[183][26] ), .IN2(n1267), .S(n7754), .Q(n13926)
         );
  MUX21X1 U12400 ( .IN1(\mem3[183][25] ), .IN2(n1245), .S(n7754), .Q(n13925)
         );
  MUX21X1 U12401 ( .IN1(\mem3[183][24] ), .IN2(n1223), .S(n7754), .Q(n13924)
         );
  AND2X1 U12402 ( .IN1(n7746), .IN2(n7116), .Q(n7754) );
  MUX21X1 U12403 ( .IN1(\mem3[182][31] ), .IN2(n1377), .S(n7755), .Q(n13923)
         );
  MUX21X1 U12404 ( .IN1(\mem3[182][30] ), .IN2(n1355), .S(n7755), .Q(n13922)
         );
  MUX21X1 U12405 ( .IN1(\mem3[182][29] ), .IN2(n1333), .S(n7755), .Q(n13921)
         );
  MUX21X1 U12406 ( .IN1(\mem3[182][28] ), .IN2(n1311), .S(n7755), .Q(n13920)
         );
  MUX21X1 U12407 ( .IN1(\mem3[182][27] ), .IN2(n1289), .S(n7755), .Q(n13919)
         );
  MUX21X1 U12408 ( .IN1(\mem3[182][26] ), .IN2(n1267), .S(n7755), .Q(n13918)
         );
  MUX21X1 U12409 ( .IN1(\mem3[182][25] ), .IN2(n1245), .S(n7755), .Q(n13917)
         );
  MUX21X1 U12410 ( .IN1(\mem3[182][24] ), .IN2(n1223), .S(n7755), .Q(n13916)
         );
  AND2X1 U12411 ( .IN1(n7746), .IN2(n7118), .Q(n7755) );
  MUX21X1 U12412 ( .IN1(\mem3[181][31] ), .IN2(n1377), .S(n7756), .Q(n13915)
         );
  MUX21X1 U12413 ( .IN1(\mem3[181][30] ), .IN2(n1355), .S(n7756), .Q(n13914)
         );
  MUX21X1 U12414 ( .IN1(\mem3[181][29] ), .IN2(n1333), .S(n7756), .Q(n13913)
         );
  MUX21X1 U12415 ( .IN1(\mem3[181][28] ), .IN2(n1311), .S(n7756), .Q(n13912)
         );
  MUX21X1 U12416 ( .IN1(\mem3[181][27] ), .IN2(n1289), .S(n7756), .Q(n13911)
         );
  MUX21X1 U12417 ( .IN1(\mem3[181][26] ), .IN2(n1267), .S(n7756), .Q(n13910)
         );
  MUX21X1 U12418 ( .IN1(\mem3[181][25] ), .IN2(n1245), .S(n7756), .Q(n13909)
         );
  MUX21X1 U12419 ( .IN1(\mem3[181][24] ), .IN2(n1223), .S(n7756), .Q(n13908)
         );
  AND2X1 U12420 ( .IN1(n7746), .IN2(n7120), .Q(n7756) );
  MUX21X1 U12421 ( .IN1(\mem3[180][31] ), .IN2(n1377), .S(n7757), .Q(n13907)
         );
  MUX21X1 U12422 ( .IN1(\mem3[180][30] ), .IN2(n1355), .S(n7757), .Q(n13906)
         );
  MUX21X1 U12423 ( .IN1(\mem3[180][29] ), .IN2(n1333), .S(n7757), .Q(n13905)
         );
  MUX21X1 U12424 ( .IN1(\mem3[180][28] ), .IN2(n1311), .S(n7757), .Q(n13904)
         );
  MUX21X1 U12425 ( .IN1(\mem3[180][27] ), .IN2(n1289), .S(n7757), .Q(n13903)
         );
  MUX21X1 U12426 ( .IN1(\mem3[180][26] ), .IN2(n1267), .S(n7757), .Q(n13902)
         );
  MUX21X1 U12427 ( .IN1(\mem3[180][25] ), .IN2(n1245), .S(n7757), .Q(n13901)
         );
  MUX21X1 U12428 ( .IN1(\mem3[180][24] ), .IN2(n1223), .S(n7757), .Q(n13900)
         );
  AND2X1 U12429 ( .IN1(n7746), .IN2(n7122), .Q(n7757) );
  MUX21X1 U12430 ( .IN1(\mem3[179][31] ), .IN2(n1377), .S(n7758), .Q(n13899)
         );
  MUX21X1 U12431 ( .IN1(\mem3[179][30] ), .IN2(n1355), .S(n7758), .Q(n13898)
         );
  MUX21X1 U12432 ( .IN1(\mem3[179][29] ), .IN2(n1333), .S(n7758), .Q(n13897)
         );
  MUX21X1 U12433 ( .IN1(\mem3[179][28] ), .IN2(n1311), .S(n7758), .Q(n13896)
         );
  MUX21X1 U12434 ( .IN1(\mem3[179][27] ), .IN2(n1289), .S(n7758), .Q(n13895)
         );
  MUX21X1 U12435 ( .IN1(\mem3[179][26] ), .IN2(n1267), .S(n7758), .Q(n13894)
         );
  MUX21X1 U12436 ( .IN1(\mem3[179][25] ), .IN2(n1245), .S(n7758), .Q(n13893)
         );
  MUX21X1 U12437 ( .IN1(\mem3[179][24] ), .IN2(n1223), .S(n7758), .Q(n13892)
         );
  AND2X1 U12438 ( .IN1(n7746), .IN2(n7124), .Q(n7758) );
  MUX21X1 U12439 ( .IN1(\mem3[178][31] ), .IN2(n1377), .S(n7759), .Q(n13891)
         );
  MUX21X1 U12440 ( .IN1(\mem3[178][30] ), .IN2(n1355), .S(n7759), .Q(n13890)
         );
  MUX21X1 U12441 ( .IN1(\mem3[178][29] ), .IN2(n1333), .S(n7759), .Q(n13889)
         );
  MUX21X1 U12442 ( .IN1(\mem3[178][28] ), .IN2(n1311), .S(n7759), .Q(n13888)
         );
  MUX21X1 U12443 ( .IN1(\mem3[178][27] ), .IN2(n1289), .S(n7759), .Q(n13887)
         );
  MUX21X1 U12444 ( .IN1(\mem3[178][26] ), .IN2(n1267), .S(n7759), .Q(n13886)
         );
  MUX21X1 U12445 ( .IN1(\mem3[178][25] ), .IN2(n1245), .S(n7759), .Q(n13885)
         );
  MUX21X1 U12446 ( .IN1(\mem3[178][24] ), .IN2(n1223), .S(n7759), .Q(n13884)
         );
  AND2X1 U12447 ( .IN1(n7746), .IN2(n7126), .Q(n7759) );
  MUX21X1 U12448 ( .IN1(\mem3[177][31] ), .IN2(n1377), .S(n7760), .Q(n13883)
         );
  MUX21X1 U12449 ( .IN1(\mem3[177][30] ), .IN2(n1355), .S(n7760), .Q(n13882)
         );
  MUX21X1 U12450 ( .IN1(\mem3[177][29] ), .IN2(n1333), .S(n7760), .Q(n13881)
         );
  MUX21X1 U12451 ( .IN1(\mem3[177][28] ), .IN2(n1311), .S(n7760), .Q(n13880)
         );
  MUX21X1 U12452 ( .IN1(\mem3[177][27] ), .IN2(n1289), .S(n7760), .Q(n13879)
         );
  MUX21X1 U12453 ( .IN1(\mem3[177][26] ), .IN2(n1267), .S(n7760), .Q(n13878)
         );
  MUX21X1 U12454 ( .IN1(\mem3[177][25] ), .IN2(n1245), .S(n7760), .Q(n13877)
         );
  MUX21X1 U12455 ( .IN1(\mem3[177][24] ), .IN2(n1223), .S(n7760), .Q(n13876)
         );
  AND2X1 U12456 ( .IN1(n7746), .IN2(n7128), .Q(n7760) );
  MUX21X1 U12457 ( .IN1(\mem3[176][31] ), .IN2(n1377), .S(n7761), .Q(n13875)
         );
  MUX21X1 U12458 ( .IN1(\mem3[176][30] ), .IN2(n1355), .S(n7761), .Q(n13874)
         );
  MUX21X1 U12459 ( .IN1(\mem3[176][29] ), .IN2(n1333), .S(n7761), .Q(n13873)
         );
  MUX21X1 U12460 ( .IN1(\mem3[176][28] ), .IN2(n1311), .S(n7761), .Q(n13872)
         );
  MUX21X1 U12461 ( .IN1(\mem3[176][27] ), .IN2(n1289), .S(n7761), .Q(n13871)
         );
  MUX21X1 U12462 ( .IN1(\mem3[176][26] ), .IN2(n1267), .S(n7761), .Q(n13870)
         );
  MUX21X1 U12463 ( .IN1(\mem3[176][25] ), .IN2(n1245), .S(n7761), .Q(n13869)
         );
  MUX21X1 U12464 ( .IN1(\mem3[176][24] ), .IN2(n1223), .S(n7761), .Q(n13868)
         );
  AND2X1 U12465 ( .IN1(n7746), .IN2(n7130), .Q(n7761) );
  AND2X1 U12466 ( .IN1(n7693), .IN2(n7204), .Q(n7746) );
  MUX21X1 U12467 ( .IN1(\mem3[175][31] ), .IN2(n1377), .S(n7762), .Q(n13867)
         );
  MUX21X1 U12468 ( .IN1(\mem3[175][30] ), .IN2(n1355), .S(n7762), .Q(n13866)
         );
  MUX21X1 U12469 ( .IN1(\mem3[175][29] ), .IN2(n1333), .S(n7762), .Q(n13865)
         );
  MUX21X1 U12470 ( .IN1(\mem3[175][28] ), .IN2(n1311), .S(n7762), .Q(n13864)
         );
  MUX21X1 U12471 ( .IN1(\mem3[175][27] ), .IN2(n1289), .S(n7762), .Q(n13863)
         );
  MUX21X1 U12472 ( .IN1(\mem3[175][26] ), .IN2(n1267), .S(n7762), .Q(n13862)
         );
  MUX21X1 U12473 ( .IN1(\mem3[175][25] ), .IN2(n1245), .S(n7762), .Q(n13861)
         );
  MUX21X1 U12474 ( .IN1(\mem3[175][24] ), .IN2(n1223), .S(n7762), .Q(n13860)
         );
  AND2X1 U12475 ( .IN1(n7763), .IN2(n7099), .Q(n7762) );
  MUX21X1 U12476 ( .IN1(\mem3[174][31] ), .IN2(n1377), .S(n7764), .Q(n13859)
         );
  MUX21X1 U12477 ( .IN1(\mem3[174][30] ), .IN2(n1355), .S(n7764), .Q(n13858)
         );
  MUX21X1 U12478 ( .IN1(\mem3[174][29] ), .IN2(n1333), .S(n7764), .Q(n13857)
         );
  MUX21X1 U12479 ( .IN1(\mem3[174][28] ), .IN2(n1311), .S(n7764), .Q(n13856)
         );
  MUX21X1 U12480 ( .IN1(\mem3[174][27] ), .IN2(n1289), .S(n7764), .Q(n13855)
         );
  MUX21X1 U12481 ( .IN1(\mem3[174][26] ), .IN2(n1267), .S(n7764), .Q(n13854)
         );
  MUX21X1 U12482 ( .IN1(\mem3[174][25] ), .IN2(n1245), .S(n7764), .Q(n13853)
         );
  MUX21X1 U12483 ( .IN1(\mem3[174][24] ), .IN2(n1223), .S(n7764), .Q(n13852)
         );
  AND2X1 U12484 ( .IN1(n7763), .IN2(n7102), .Q(n7764) );
  MUX21X1 U12485 ( .IN1(\mem3[173][31] ), .IN2(n1377), .S(n7765), .Q(n13851)
         );
  MUX21X1 U12486 ( .IN1(\mem3[173][30] ), .IN2(n1355), .S(n7765), .Q(n13850)
         );
  MUX21X1 U12487 ( .IN1(\mem3[173][29] ), .IN2(n1333), .S(n7765), .Q(n13849)
         );
  MUX21X1 U12488 ( .IN1(\mem3[173][28] ), .IN2(n1311), .S(n7765), .Q(n13848)
         );
  MUX21X1 U12489 ( .IN1(\mem3[173][27] ), .IN2(n1289), .S(n7765), .Q(n13847)
         );
  MUX21X1 U12490 ( .IN1(\mem3[173][26] ), .IN2(n1267), .S(n7765), .Q(n13846)
         );
  MUX21X1 U12491 ( .IN1(\mem3[173][25] ), .IN2(n1245), .S(n7765), .Q(n13845)
         );
  MUX21X1 U12492 ( .IN1(\mem3[173][24] ), .IN2(n1223), .S(n7765), .Q(n13844)
         );
  AND2X1 U12493 ( .IN1(n7763), .IN2(n7104), .Q(n7765) );
  MUX21X1 U12494 ( .IN1(\mem3[172][31] ), .IN2(n1377), .S(n7766), .Q(n13843)
         );
  MUX21X1 U12495 ( .IN1(\mem3[172][30] ), .IN2(n1355), .S(n7766), .Q(n13842)
         );
  MUX21X1 U12496 ( .IN1(\mem3[172][29] ), .IN2(n1333), .S(n7766), .Q(n13841)
         );
  MUX21X1 U12497 ( .IN1(\mem3[172][28] ), .IN2(n1311), .S(n7766), .Q(n13840)
         );
  MUX21X1 U12498 ( .IN1(\mem3[172][27] ), .IN2(n1289), .S(n7766), .Q(n13839)
         );
  MUX21X1 U12499 ( .IN1(\mem3[172][26] ), .IN2(n1267), .S(n7766), .Q(n13838)
         );
  MUX21X1 U12500 ( .IN1(\mem3[172][25] ), .IN2(n1245), .S(n7766), .Q(n13837)
         );
  MUX21X1 U12501 ( .IN1(\mem3[172][24] ), .IN2(n1223), .S(n7766), .Q(n13836)
         );
  AND2X1 U12502 ( .IN1(n7763), .IN2(n7106), .Q(n7766) );
  MUX21X1 U12503 ( .IN1(\mem3[171][31] ), .IN2(n1378), .S(n7767), .Q(n13835)
         );
  MUX21X1 U12504 ( .IN1(\mem3[171][30] ), .IN2(n1356), .S(n7767), .Q(n13834)
         );
  MUX21X1 U12505 ( .IN1(\mem3[171][29] ), .IN2(n1334), .S(n7767), .Q(n13833)
         );
  MUX21X1 U12506 ( .IN1(\mem3[171][28] ), .IN2(n1312), .S(n7767), .Q(n13832)
         );
  MUX21X1 U12507 ( .IN1(\mem3[171][27] ), .IN2(n1290), .S(n7767), .Q(n13831)
         );
  MUX21X1 U12508 ( .IN1(\mem3[171][26] ), .IN2(n1268), .S(n7767), .Q(n13830)
         );
  MUX21X1 U12509 ( .IN1(\mem3[171][25] ), .IN2(n1246), .S(n7767), .Q(n13829)
         );
  MUX21X1 U12510 ( .IN1(\mem3[171][24] ), .IN2(n1224), .S(n7767), .Q(n13828)
         );
  AND2X1 U12511 ( .IN1(n7763), .IN2(n7108), .Q(n7767) );
  MUX21X1 U12512 ( .IN1(\mem3[170][31] ), .IN2(n1378), .S(n7768), .Q(n13827)
         );
  MUX21X1 U12513 ( .IN1(\mem3[170][30] ), .IN2(n1356), .S(n7768), .Q(n13826)
         );
  MUX21X1 U12514 ( .IN1(\mem3[170][29] ), .IN2(n1334), .S(n7768), .Q(n13825)
         );
  MUX21X1 U12515 ( .IN1(\mem3[170][28] ), .IN2(n1312), .S(n7768), .Q(n13824)
         );
  MUX21X1 U12516 ( .IN1(\mem3[170][27] ), .IN2(n1290), .S(n7768), .Q(n13823)
         );
  MUX21X1 U12517 ( .IN1(\mem3[170][26] ), .IN2(n1268), .S(n7768), .Q(n13822)
         );
  MUX21X1 U12518 ( .IN1(\mem3[170][25] ), .IN2(n1246), .S(n7768), .Q(n13821)
         );
  MUX21X1 U12519 ( .IN1(\mem3[170][24] ), .IN2(n1224), .S(n7768), .Q(n13820)
         );
  AND2X1 U12520 ( .IN1(n7763), .IN2(n7110), .Q(n7768) );
  MUX21X1 U12521 ( .IN1(\mem3[169][31] ), .IN2(n1378), .S(n7769), .Q(n13819)
         );
  MUX21X1 U12522 ( .IN1(\mem3[169][30] ), .IN2(n1356), .S(n7769), .Q(n13818)
         );
  MUX21X1 U12523 ( .IN1(\mem3[169][29] ), .IN2(n1334), .S(n7769), .Q(n13817)
         );
  MUX21X1 U12524 ( .IN1(\mem3[169][28] ), .IN2(n1312), .S(n7769), .Q(n13816)
         );
  MUX21X1 U12525 ( .IN1(\mem3[169][27] ), .IN2(n1290), .S(n7769), .Q(n13815)
         );
  MUX21X1 U12526 ( .IN1(\mem3[169][26] ), .IN2(n1268), .S(n7769), .Q(n13814)
         );
  MUX21X1 U12527 ( .IN1(\mem3[169][25] ), .IN2(n1246), .S(n7769), .Q(n13813)
         );
  MUX21X1 U12528 ( .IN1(\mem3[169][24] ), .IN2(n1224), .S(n7769), .Q(n13812)
         );
  AND2X1 U12529 ( .IN1(n7763), .IN2(n7112), .Q(n7769) );
  MUX21X1 U12530 ( .IN1(\mem3[168][31] ), .IN2(n1378), .S(n7770), .Q(n13811)
         );
  MUX21X1 U12531 ( .IN1(\mem3[168][30] ), .IN2(n1356), .S(n7770), .Q(n13810)
         );
  MUX21X1 U12532 ( .IN1(\mem3[168][29] ), .IN2(n1334), .S(n7770), .Q(n13809)
         );
  MUX21X1 U12533 ( .IN1(\mem3[168][28] ), .IN2(n1312), .S(n7770), .Q(n13808)
         );
  MUX21X1 U12534 ( .IN1(\mem3[168][27] ), .IN2(n1290), .S(n7770), .Q(n13807)
         );
  MUX21X1 U12535 ( .IN1(\mem3[168][26] ), .IN2(n1268), .S(n7770), .Q(n13806)
         );
  MUX21X1 U12536 ( .IN1(\mem3[168][25] ), .IN2(n1246), .S(n7770), .Q(n13805)
         );
  MUX21X1 U12537 ( .IN1(\mem3[168][24] ), .IN2(n1224), .S(n7770), .Q(n13804)
         );
  AND2X1 U12538 ( .IN1(n7763), .IN2(n7114), .Q(n7770) );
  MUX21X1 U12539 ( .IN1(\mem3[167][31] ), .IN2(n1378), .S(n7771), .Q(n13803)
         );
  MUX21X1 U12540 ( .IN1(\mem3[167][30] ), .IN2(n1356), .S(n7771), .Q(n13802)
         );
  MUX21X1 U12541 ( .IN1(\mem3[167][29] ), .IN2(n1334), .S(n7771), .Q(n13801)
         );
  MUX21X1 U12542 ( .IN1(\mem3[167][28] ), .IN2(n1312), .S(n7771), .Q(n13800)
         );
  MUX21X1 U12543 ( .IN1(\mem3[167][27] ), .IN2(n1290), .S(n7771), .Q(n13799)
         );
  MUX21X1 U12544 ( .IN1(\mem3[167][26] ), .IN2(n1268), .S(n7771), .Q(n13798)
         );
  MUX21X1 U12545 ( .IN1(\mem3[167][25] ), .IN2(n1246), .S(n7771), .Q(n13797)
         );
  MUX21X1 U12546 ( .IN1(\mem3[167][24] ), .IN2(n1224), .S(n7771), .Q(n13796)
         );
  AND2X1 U12547 ( .IN1(n7763), .IN2(n7116), .Q(n7771) );
  MUX21X1 U12548 ( .IN1(\mem3[166][31] ), .IN2(n1378), .S(n7772), .Q(n13795)
         );
  MUX21X1 U12549 ( .IN1(\mem3[166][30] ), .IN2(n1356), .S(n7772), .Q(n13794)
         );
  MUX21X1 U12550 ( .IN1(\mem3[166][29] ), .IN2(n1334), .S(n7772), .Q(n13793)
         );
  MUX21X1 U12551 ( .IN1(\mem3[166][28] ), .IN2(n1312), .S(n7772), .Q(n13792)
         );
  MUX21X1 U12552 ( .IN1(\mem3[166][27] ), .IN2(n1290), .S(n7772), .Q(n13791)
         );
  MUX21X1 U12553 ( .IN1(\mem3[166][26] ), .IN2(n1268), .S(n7772), .Q(n13790)
         );
  MUX21X1 U12554 ( .IN1(\mem3[166][25] ), .IN2(n1246), .S(n7772), .Q(n13789)
         );
  MUX21X1 U12555 ( .IN1(\mem3[166][24] ), .IN2(n1224), .S(n7772), .Q(n13788)
         );
  AND2X1 U12556 ( .IN1(n7763), .IN2(n7118), .Q(n7772) );
  MUX21X1 U12557 ( .IN1(\mem3[165][31] ), .IN2(n1378), .S(n7773), .Q(n13787)
         );
  MUX21X1 U12558 ( .IN1(\mem3[165][30] ), .IN2(n1356), .S(n7773), .Q(n13786)
         );
  MUX21X1 U12559 ( .IN1(\mem3[165][29] ), .IN2(n1334), .S(n7773), .Q(n13785)
         );
  MUX21X1 U12560 ( .IN1(\mem3[165][28] ), .IN2(n1312), .S(n7773), .Q(n13784)
         );
  MUX21X1 U12561 ( .IN1(\mem3[165][27] ), .IN2(n1290), .S(n7773), .Q(n13783)
         );
  MUX21X1 U12562 ( .IN1(\mem3[165][26] ), .IN2(n1268), .S(n7773), .Q(n13782)
         );
  MUX21X1 U12563 ( .IN1(\mem3[165][25] ), .IN2(n1246), .S(n7773), .Q(n13781)
         );
  MUX21X1 U12564 ( .IN1(\mem3[165][24] ), .IN2(n1224), .S(n7773), .Q(n13780)
         );
  AND2X1 U12565 ( .IN1(n7763), .IN2(n7120), .Q(n7773) );
  MUX21X1 U12566 ( .IN1(\mem3[164][31] ), .IN2(n1378), .S(n7774), .Q(n13779)
         );
  MUX21X1 U12567 ( .IN1(\mem3[164][30] ), .IN2(n1356), .S(n7774), .Q(n13778)
         );
  MUX21X1 U12568 ( .IN1(\mem3[164][29] ), .IN2(n1334), .S(n7774), .Q(n13777)
         );
  MUX21X1 U12569 ( .IN1(\mem3[164][28] ), .IN2(n1312), .S(n7774), .Q(n13776)
         );
  MUX21X1 U12570 ( .IN1(\mem3[164][27] ), .IN2(n1290), .S(n7774), .Q(n13775)
         );
  MUX21X1 U12571 ( .IN1(\mem3[164][26] ), .IN2(n1268), .S(n7774), .Q(n13774)
         );
  MUX21X1 U12572 ( .IN1(\mem3[164][25] ), .IN2(n1246), .S(n7774), .Q(n13773)
         );
  MUX21X1 U12573 ( .IN1(\mem3[164][24] ), .IN2(n1224), .S(n7774), .Q(n13772)
         );
  AND2X1 U12574 ( .IN1(n7763), .IN2(n7122), .Q(n7774) );
  MUX21X1 U12575 ( .IN1(\mem3[163][31] ), .IN2(n1378), .S(n7775), .Q(n13771)
         );
  MUX21X1 U12576 ( .IN1(\mem3[163][30] ), .IN2(n1356), .S(n7775), .Q(n13770)
         );
  MUX21X1 U12577 ( .IN1(\mem3[163][29] ), .IN2(n1334), .S(n7775), .Q(n13769)
         );
  MUX21X1 U12578 ( .IN1(\mem3[163][28] ), .IN2(n1312), .S(n7775), .Q(n13768)
         );
  MUX21X1 U12579 ( .IN1(\mem3[163][27] ), .IN2(n1290), .S(n7775), .Q(n13767)
         );
  MUX21X1 U12580 ( .IN1(\mem3[163][26] ), .IN2(n1268), .S(n7775), .Q(n13766)
         );
  MUX21X1 U12581 ( .IN1(\mem3[163][25] ), .IN2(n1246), .S(n7775), .Q(n13765)
         );
  MUX21X1 U12582 ( .IN1(\mem3[163][24] ), .IN2(n1224), .S(n7775), .Q(n13764)
         );
  AND2X1 U12583 ( .IN1(n7763), .IN2(n7124), .Q(n7775) );
  MUX21X1 U12584 ( .IN1(\mem3[162][31] ), .IN2(n1378), .S(n7776), .Q(n13763)
         );
  MUX21X1 U12585 ( .IN1(\mem3[162][30] ), .IN2(n1356), .S(n7776), .Q(n13762)
         );
  MUX21X1 U12586 ( .IN1(\mem3[162][29] ), .IN2(n1334), .S(n7776), .Q(n13761)
         );
  MUX21X1 U12587 ( .IN1(\mem3[162][28] ), .IN2(n1312), .S(n7776), .Q(n13760)
         );
  MUX21X1 U12588 ( .IN1(\mem3[162][27] ), .IN2(n1290), .S(n7776), .Q(n13759)
         );
  MUX21X1 U12589 ( .IN1(\mem3[162][26] ), .IN2(n1268), .S(n7776), .Q(n13758)
         );
  MUX21X1 U12590 ( .IN1(\mem3[162][25] ), .IN2(n1246), .S(n7776), .Q(n13757)
         );
  MUX21X1 U12591 ( .IN1(\mem3[162][24] ), .IN2(n1224), .S(n7776), .Q(n13756)
         );
  AND2X1 U12592 ( .IN1(n7763), .IN2(n7126), .Q(n7776) );
  MUX21X1 U12593 ( .IN1(\mem3[161][31] ), .IN2(n1378), .S(n7777), .Q(n13755)
         );
  MUX21X1 U12594 ( .IN1(\mem3[161][30] ), .IN2(n1356), .S(n7777), .Q(n13754)
         );
  MUX21X1 U12595 ( .IN1(\mem3[161][29] ), .IN2(n1334), .S(n7777), .Q(n13753)
         );
  MUX21X1 U12596 ( .IN1(\mem3[161][28] ), .IN2(n1312), .S(n7777), .Q(n13752)
         );
  MUX21X1 U12597 ( .IN1(\mem3[161][27] ), .IN2(n1290), .S(n7777), .Q(n13751)
         );
  MUX21X1 U12598 ( .IN1(\mem3[161][26] ), .IN2(n1268), .S(n7777), .Q(n13750)
         );
  MUX21X1 U12599 ( .IN1(\mem3[161][25] ), .IN2(n1246), .S(n7777), .Q(n13749)
         );
  MUX21X1 U12600 ( .IN1(\mem3[161][24] ), .IN2(n1224), .S(n7777), .Q(n13748)
         );
  AND2X1 U12601 ( .IN1(n7763), .IN2(n7128), .Q(n7777) );
  MUX21X1 U12602 ( .IN1(\mem3[160][31] ), .IN2(n1378), .S(n7778), .Q(n13747)
         );
  MUX21X1 U12603 ( .IN1(\mem3[160][30] ), .IN2(n1356), .S(n7778), .Q(n13746)
         );
  MUX21X1 U12604 ( .IN1(\mem3[160][29] ), .IN2(n1334), .S(n7778), .Q(n13745)
         );
  MUX21X1 U12605 ( .IN1(\mem3[160][28] ), .IN2(n1312), .S(n7778), .Q(n13744)
         );
  MUX21X1 U12606 ( .IN1(\mem3[160][27] ), .IN2(n1290), .S(n7778), .Q(n13743)
         );
  MUX21X1 U12607 ( .IN1(\mem3[160][26] ), .IN2(n1268), .S(n7778), .Q(n13742)
         );
  MUX21X1 U12608 ( .IN1(\mem3[160][25] ), .IN2(n1246), .S(n7778), .Q(n13741)
         );
  MUX21X1 U12609 ( .IN1(\mem3[160][24] ), .IN2(n1224), .S(n7778), .Q(n13740)
         );
  AND2X1 U12610 ( .IN1(n7763), .IN2(n7130), .Q(n7778) );
  AND2X1 U12611 ( .IN1(n7693), .IN2(n7222), .Q(n7763) );
  MUX21X1 U12612 ( .IN1(\mem3[159][31] ), .IN2(n1379), .S(n7779), .Q(n13739)
         );
  MUX21X1 U12613 ( .IN1(\mem3[159][30] ), .IN2(n1357), .S(n7779), .Q(n13738)
         );
  MUX21X1 U12614 ( .IN1(\mem3[159][29] ), .IN2(n1335), .S(n7779), .Q(n13737)
         );
  MUX21X1 U12615 ( .IN1(\mem3[159][28] ), .IN2(n1313), .S(n7779), .Q(n13736)
         );
  MUX21X1 U12616 ( .IN1(\mem3[159][27] ), .IN2(n1291), .S(n7779), .Q(n13735)
         );
  MUX21X1 U12617 ( .IN1(\mem3[159][26] ), .IN2(n1269), .S(n7779), .Q(n13734)
         );
  MUX21X1 U12618 ( .IN1(\mem3[159][25] ), .IN2(n1247), .S(n7779), .Q(n13733)
         );
  MUX21X1 U12619 ( .IN1(\mem3[159][24] ), .IN2(n1225), .S(n7779), .Q(n13732)
         );
  AND2X1 U12620 ( .IN1(n7780), .IN2(n7099), .Q(n7779) );
  MUX21X1 U12621 ( .IN1(\mem3[158][31] ), .IN2(n1379), .S(n7781), .Q(n13731)
         );
  MUX21X1 U12622 ( .IN1(\mem3[158][30] ), .IN2(n1357), .S(n7781), .Q(n13730)
         );
  MUX21X1 U12623 ( .IN1(\mem3[158][29] ), .IN2(n1335), .S(n7781), .Q(n13729)
         );
  MUX21X1 U12624 ( .IN1(\mem3[158][28] ), .IN2(n1313), .S(n7781), .Q(n13728)
         );
  MUX21X1 U12625 ( .IN1(\mem3[158][27] ), .IN2(n1291), .S(n7781), .Q(n13727)
         );
  MUX21X1 U12626 ( .IN1(\mem3[158][26] ), .IN2(n1269), .S(n7781), .Q(n13726)
         );
  MUX21X1 U12627 ( .IN1(\mem3[158][25] ), .IN2(n1247), .S(n7781), .Q(n13725)
         );
  MUX21X1 U12628 ( .IN1(\mem3[158][24] ), .IN2(n1225), .S(n7781), .Q(n13724)
         );
  AND2X1 U12629 ( .IN1(n7780), .IN2(n7102), .Q(n7781) );
  MUX21X1 U12630 ( .IN1(\mem3[157][31] ), .IN2(n1379), .S(n7782), .Q(n13723)
         );
  MUX21X1 U12631 ( .IN1(\mem3[157][30] ), .IN2(n1357), .S(n7782), .Q(n13722)
         );
  MUX21X1 U12632 ( .IN1(\mem3[157][29] ), .IN2(n1335), .S(n7782), .Q(n13721)
         );
  MUX21X1 U12633 ( .IN1(\mem3[157][28] ), .IN2(n1313), .S(n7782), .Q(n13720)
         );
  MUX21X1 U12634 ( .IN1(\mem3[157][27] ), .IN2(n1291), .S(n7782), .Q(n13719)
         );
  MUX21X1 U12635 ( .IN1(\mem3[157][26] ), .IN2(n1269), .S(n7782), .Q(n13718)
         );
  MUX21X1 U12636 ( .IN1(\mem3[157][25] ), .IN2(n1247), .S(n7782), .Q(n13717)
         );
  MUX21X1 U12637 ( .IN1(\mem3[157][24] ), .IN2(n1225), .S(n7782), .Q(n13716)
         );
  AND2X1 U12638 ( .IN1(n7780), .IN2(n7104), .Q(n7782) );
  MUX21X1 U12639 ( .IN1(\mem3[156][31] ), .IN2(n1379), .S(n7783), .Q(n13715)
         );
  MUX21X1 U12640 ( .IN1(\mem3[156][30] ), .IN2(n1357), .S(n7783), .Q(n13714)
         );
  MUX21X1 U12641 ( .IN1(\mem3[156][29] ), .IN2(n1335), .S(n7783), .Q(n13713)
         );
  MUX21X1 U12642 ( .IN1(\mem3[156][28] ), .IN2(n1313), .S(n7783), .Q(n13712)
         );
  MUX21X1 U12643 ( .IN1(\mem3[156][27] ), .IN2(n1291), .S(n7783), .Q(n13711)
         );
  MUX21X1 U12644 ( .IN1(\mem3[156][26] ), .IN2(n1269), .S(n7783), .Q(n13710)
         );
  MUX21X1 U12645 ( .IN1(\mem3[156][25] ), .IN2(n1247), .S(n7783), .Q(n13709)
         );
  MUX21X1 U12646 ( .IN1(\mem3[156][24] ), .IN2(n1225), .S(n7783), .Q(n13708)
         );
  AND2X1 U12647 ( .IN1(n7780), .IN2(n7106), .Q(n7783) );
  MUX21X1 U12648 ( .IN1(\mem3[155][31] ), .IN2(n1379), .S(n7784), .Q(n13707)
         );
  MUX21X1 U12649 ( .IN1(\mem3[155][30] ), .IN2(n1357), .S(n7784), .Q(n13706)
         );
  MUX21X1 U12650 ( .IN1(\mem3[155][29] ), .IN2(n1335), .S(n7784), .Q(n13705)
         );
  MUX21X1 U12651 ( .IN1(\mem3[155][28] ), .IN2(n1313), .S(n7784), .Q(n13704)
         );
  MUX21X1 U12652 ( .IN1(\mem3[155][27] ), .IN2(n1291), .S(n7784), .Q(n13703)
         );
  MUX21X1 U12653 ( .IN1(\mem3[155][26] ), .IN2(n1269), .S(n7784), .Q(n13702)
         );
  MUX21X1 U12654 ( .IN1(\mem3[155][25] ), .IN2(n1247), .S(n7784), .Q(n13701)
         );
  MUX21X1 U12655 ( .IN1(\mem3[155][24] ), .IN2(n1225), .S(n7784), .Q(n13700)
         );
  AND2X1 U12656 ( .IN1(n7780), .IN2(n7108), .Q(n7784) );
  MUX21X1 U12657 ( .IN1(\mem3[154][31] ), .IN2(n1379), .S(n7785), .Q(n13699)
         );
  MUX21X1 U12658 ( .IN1(\mem3[154][30] ), .IN2(n1357), .S(n7785), .Q(n13698)
         );
  MUX21X1 U12659 ( .IN1(\mem3[154][29] ), .IN2(n1335), .S(n7785), .Q(n13697)
         );
  MUX21X1 U12660 ( .IN1(\mem3[154][28] ), .IN2(n1313), .S(n7785), .Q(n13696)
         );
  MUX21X1 U12661 ( .IN1(\mem3[154][27] ), .IN2(n1291), .S(n7785), .Q(n13695)
         );
  MUX21X1 U12662 ( .IN1(\mem3[154][26] ), .IN2(n1269), .S(n7785), .Q(n13694)
         );
  MUX21X1 U12663 ( .IN1(\mem3[154][25] ), .IN2(n1247), .S(n7785), .Q(n13693)
         );
  MUX21X1 U12664 ( .IN1(\mem3[154][24] ), .IN2(n1225), .S(n7785), .Q(n13692)
         );
  AND2X1 U12665 ( .IN1(n7780), .IN2(n7110), .Q(n7785) );
  MUX21X1 U12666 ( .IN1(\mem3[153][31] ), .IN2(n1379), .S(n7786), .Q(n13691)
         );
  MUX21X1 U12667 ( .IN1(\mem3[153][30] ), .IN2(n1357), .S(n7786), .Q(n13690)
         );
  MUX21X1 U12668 ( .IN1(\mem3[153][29] ), .IN2(n1335), .S(n7786), .Q(n13689)
         );
  MUX21X1 U12669 ( .IN1(\mem3[153][28] ), .IN2(n1313), .S(n7786), .Q(n13688)
         );
  MUX21X1 U12670 ( .IN1(\mem3[153][27] ), .IN2(n1291), .S(n7786), .Q(n13687)
         );
  MUX21X1 U12671 ( .IN1(\mem3[153][26] ), .IN2(n1269), .S(n7786), .Q(n13686)
         );
  MUX21X1 U12672 ( .IN1(\mem3[153][25] ), .IN2(n1247), .S(n7786), .Q(n13685)
         );
  MUX21X1 U12673 ( .IN1(\mem3[153][24] ), .IN2(n1225), .S(n7786), .Q(n13684)
         );
  AND2X1 U12674 ( .IN1(n7780), .IN2(n7112), .Q(n7786) );
  MUX21X1 U12675 ( .IN1(\mem3[152][31] ), .IN2(n1379), .S(n7787), .Q(n13683)
         );
  MUX21X1 U12676 ( .IN1(\mem3[152][30] ), .IN2(n1357), .S(n7787), .Q(n13682)
         );
  MUX21X1 U12677 ( .IN1(\mem3[152][29] ), .IN2(n1335), .S(n7787), .Q(n13681)
         );
  MUX21X1 U12678 ( .IN1(\mem3[152][28] ), .IN2(n1313), .S(n7787), .Q(n13680)
         );
  MUX21X1 U12679 ( .IN1(\mem3[152][27] ), .IN2(n1291), .S(n7787), .Q(n13679)
         );
  MUX21X1 U12680 ( .IN1(\mem3[152][26] ), .IN2(n1269), .S(n7787), .Q(n13678)
         );
  MUX21X1 U12681 ( .IN1(\mem3[152][25] ), .IN2(n1247), .S(n7787), .Q(n13677)
         );
  MUX21X1 U12682 ( .IN1(\mem3[152][24] ), .IN2(n1225), .S(n7787), .Q(n13676)
         );
  AND2X1 U12683 ( .IN1(n7780), .IN2(n7114), .Q(n7787) );
  MUX21X1 U12684 ( .IN1(\mem3[151][31] ), .IN2(n1379), .S(n7788), .Q(n13675)
         );
  MUX21X1 U12685 ( .IN1(\mem3[151][30] ), .IN2(n1357), .S(n7788), .Q(n13674)
         );
  MUX21X1 U12686 ( .IN1(\mem3[151][29] ), .IN2(n1335), .S(n7788), .Q(n13673)
         );
  MUX21X1 U12687 ( .IN1(\mem3[151][28] ), .IN2(n1313), .S(n7788), .Q(n13672)
         );
  MUX21X1 U12688 ( .IN1(\mem3[151][27] ), .IN2(n1291), .S(n7788), .Q(n13671)
         );
  MUX21X1 U12689 ( .IN1(\mem3[151][26] ), .IN2(n1269), .S(n7788), .Q(n13670)
         );
  MUX21X1 U12690 ( .IN1(\mem3[151][25] ), .IN2(n1247), .S(n7788), .Q(n13669)
         );
  MUX21X1 U12691 ( .IN1(\mem3[151][24] ), .IN2(n1225), .S(n7788), .Q(n13668)
         );
  AND2X1 U12692 ( .IN1(n7780), .IN2(n7116), .Q(n7788) );
  MUX21X1 U12693 ( .IN1(\mem3[150][31] ), .IN2(n1379), .S(n7789), .Q(n13667)
         );
  MUX21X1 U12694 ( .IN1(\mem3[150][30] ), .IN2(n1357), .S(n7789), .Q(n13666)
         );
  MUX21X1 U12695 ( .IN1(\mem3[150][29] ), .IN2(n1335), .S(n7789), .Q(n13665)
         );
  MUX21X1 U12696 ( .IN1(\mem3[150][28] ), .IN2(n1313), .S(n7789), .Q(n13664)
         );
  MUX21X1 U12697 ( .IN1(\mem3[150][27] ), .IN2(n1291), .S(n7789), .Q(n13663)
         );
  MUX21X1 U12698 ( .IN1(\mem3[150][26] ), .IN2(n1269), .S(n7789), .Q(n13662)
         );
  MUX21X1 U12699 ( .IN1(\mem3[150][25] ), .IN2(n1247), .S(n7789), .Q(n13661)
         );
  MUX21X1 U12700 ( .IN1(\mem3[150][24] ), .IN2(n1225), .S(n7789), .Q(n13660)
         );
  AND2X1 U12701 ( .IN1(n7780), .IN2(n7118), .Q(n7789) );
  MUX21X1 U12702 ( .IN1(\mem3[149][31] ), .IN2(n1379), .S(n7790), .Q(n13659)
         );
  MUX21X1 U12703 ( .IN1(\mem3[149][30] ), .IN2(n1357), .S(n7790), .Q(n13658)
         );
  MUX21X1 U12704 ( .IN1(\mem3[149][29] ), .IN2(n1335), .S(n7790), .Q(n13657)
         );
  MUX21X1 U12705 ( .IN1(\mem3[149][28] ), .IN2(n1313), .S(n7790), .Q(n13656)
         );
  MUX21X1 U12706 ( .IN1(\mem3[149][27] ), .IN2(n1291), .S(n7790), .Q(n13655)
         );
  MUX21X1 U12707 ( .IN1(\mem3[149][26] ), .IN2(n1269), .S(n7790), .Q(n13654)
         );
  MUX21X1 U12708 ( .IN1(\mem3[149][25] ), .IN2(n1247), .S(n7790), .Q(n13653)
         );
  MUX21X1 U12709 ( .IN1(\mem3[149][24] ), .IN2(n1225), .S(n7790), .Q(n13652)
         );
  AND2X1 U12710 ( .IN1(n7780), .IN2(n7120), .Q(n7790) );
  MUX21X1 U12711 ( .IN1(\mem3[148][31] ), .IN2(n1379), .S(n7791), .Q(n13651)
         );
  MUX21X1 U12712 ( .IN1(\mem3[148][30] ), .IN2(n1357), .S(n7791), .Q(n13650)
         );
  MUX21X1 U12713 ( .IN1(\mem3[148][29] ), .IN2(n1335), .S(n7791), .Q(n13649)
         );
  MUX21X1 U12714 ( .IN1(\mem3[148][28] ), .IN2(n1313), .S(n7791), .Q(n13648)
         );
  MUX21X1 U12715 ( .IN1(\mem3[148][27] ), .IN2(n1291), .S(n7791), .Q(n13647)
         );
  MUX21X1 U12716 ( .IN1(\mem3[148][26] ), .IN2(n1269), .S(n7791), .Q(n13646)
         );
  MUX21X1 U12717 ( .IN1(\mem3[148][25] ), .IN2(n1247), .S(n7791), .Q(n13645)
         );
  MUX21X1 U12718 ( .IN1(\mem3[148][24] ), .IN2(n1225), .S(n7791), .Q(n13644)
         );
  AND2X1 U12719 ( .IN1(n7780), .IN2(n7122), .Q(n7791) );
  MUX21X1 U12720 ( .IN1(\mem3[147][31] ), .IN2(n1380), .S(n7792), .Q(n13643)
         );
  MUX21X1 U12721 ( .IN1(\mem3[147][30] ), .IN2(n1358), .S(n7792), .Q(n13642)
         );
  MUX21X1 U12722 ( .IN1(\mem3[147][29] ), .IN2(n1336), .S(n7792), .Q(n13641)
         );
  MUX21X1 U12723 ( .IN1(\mem3[147][28] ), .IN2(n1314), .S(n7792), .Q(n13640)
         );
  MUX21X1 U12724 ( .IN1(\mem3[147][27] ), .IN2(n1292), .S(n7792), .Q(n13639)
         );
  MUX21X1 U12725 ( .IN1(\mem3[147][26] ), .IN2(n1270), .S(n7792), .Q(n13638)
         );
  MUX21X1 U12726 ( .IN1(\mem3[147][25] ), .IN2(n1248), .S(n7792), .Q(n13637)
         );
  MUX21X1 U12727 ( .IN1(\mem3[147][24] ), .IN2(n1226), .S(n7792), .Q(n13636)
         );
  AND2X1 U12728 ( .IN1(n7780), .IN2(n7124), .Q(n7792) );
  MUX21X1 U12729 ( .IN1(\mem3[146][31] ), .IN2(n1380), .S(n7793), .Q(n13635)
         );
  MUX21X1 U12730 ( .IN1(\mem3[146][30] ), .IN2(n1358), .S(n7793), .Q(n13634)
         );
  MUX21X1 U12731 ( .IN1(\mem3[146][29] ), .IN2(n1336), .S(n7793), .Q(n13633)
         );
  MUX21X1 U12732 ( .IN1(\mem3[146][28] ), .IN2(n1314), .S(n7793), .Q(n13632)
         );
  MUX21X1 U12733 ( .IN1(\mem3[146][27] ), .IN2(n1292), .S(n7793), .Q(n13631)
         );
  MUX21X1 U12734 ( .IN1(\mem3[146][26] ), .IN2(n1270), .S(n7793), .Q(n13630)
         );
  MUX21X1 U12735 ( .IN1(\mem3[146][25] ), .IN2(n1248), .S(n7793), .Q(n13629)
         );
  MUX21X1 U12736 ( .IN1(\mem3[146][24] ), .IN2(n1226), .S(n7793), .Q(n13628)
         );
  AND2X1 U12737 ( .IN1(n7780), .IN2(n7126), .Q(n7793) );
  MUX21X1 U12738 ( .IN1(\mem3[145][31] ), .IN2(n1380), .S(n7794), .Q(n13627)
         );
  MUX21X1 U12739 ( .IN1(\mem3[145][30] ), .IN2(n1358), .S(n7794), .Q(n13626)
         );
  MUX21X1 U12740 ( .IN1(\mem3[145][29] ), .IN2(n1336), .S(n7794), .Q(n13625)
         );
  MUX21X1 U12741 ( .IN1(\mem3[145][28] ), .IN2(n1314), .S(n7794), .Q(n13624)
         );
  MUX21X1 U12742 ( .IN1(\mem3[145][27] ), .IN2(n1292), .S(n7794), .Q(n13623)
         );
  MUX21X1 U12743 ( .IN1(\mem3[145][26] ), .IN2(n1270), .S(n7794), .Q(n13622)
         );
  MUX21X1 U12744 ( .IN1(\mem3[145][25] ), .IN2(n1248), .S(n7794), .Q(n13621)
         );
  MUX21X1 U12745 ( .IN1(\mem3[145][24] ), .IN2(n1226), .S(n7794), .Q(n13620)
         );
  AND2X1 U12746 ( .IN1(n7780), .IN2(n7128), .Q(n7794) );
  MUX21X1 U12747 ( .IN1(\mem3[144][31] ), .IN2(n1380), .S(n7795), .Q(n13619)
         );
  MUX21X1 U12748 ( .IN1(\mem3[144][30] ), .IN2(n1358), .S(n7795), .Q(n13618)
         );
  MUX21X1 U12749 ( .IN1(\mem3[144][29] ), .IN2(n1336), .S(n7795), .Q(n13617)
         );
  MUX21X1 U12750 ( .IN1(\mem3[144][28] ), .IN2(n1314), .S(n7795), .Q(n13616)
         );
  MUX21X1 U12751 ( .IN1(\mem3[144][27] ), .IN2(n1292), .S(n7795), .Q(n13615)
         );
  MUX21X1 U12752 ( .IN1(\mem3[144][26] ), .IN2(n1270), .S(n7795), .Q(n13614)
         );
  MUX21X1 U12753 ( .IN1(\mem3[144][25] ), .IN2(n1248), .S(n7795), .Q(n13613)
         );
  MUX21X1 U12754 ( .IN1(\mem3[144][24] ), .IN2(n1226), .S(n7795), .Q(n13612)
         );
  AND2X1 U12755 ( .IN1(n7780), .IN2(n7130), .Q(n7795) );
  AND2X1 U12756 ( .IN1(n7693), .IN2(n7240), .Q(n7780) );
  MUX21X1 U12757 ( .IN1(\mem3[143][31] ), .IN2(n1380), .S(n7796), .Q(n13611)
         );
  MUX21X1 U12758 ( .IN1(\mem3[143][30] ), .IN2(n1358), .S(n7796), .Q(n13610)
         );
  MUX21X1 U12759 ( .IN1(\mem3[143][29] ), .IN2(n1336), .S(n7796), .Q(n13609)
         );
  MUX21X1 U12760 ( .IN1(\mem3[143][28] ), .IN2(n1314), .S(n7796), .Q(n13608)
         );
  MUX21X1 U12761 ( .IN1(\mem3[143][27] ), .IN2(n1292), .S(n7796), .Q(n13607)
         );
  MUX21X1 U12762 ( .IN1(\mem3[143][26] ), .IN2(n1270), .S(n7796), .Q(n13606)
         );
  MUX21X1 U12763 ( .IN1(\mem3[143][25] ), .IN2(n1248), .S(n7796), .Q(n13605)
         );
  MUX21X1 U12764 ( .IN1(\mem3[143][24] ), .IN2(n1226), .S(n7796), .Q(n13604)
         );
  AND2X1 U12765 ( .IN1(n7797), .IN2(n7099), .Q(n7796) );
  MUX21X1 U12766 ( .IN1(\mem3[142][31] ), .IN2(n1380), .S(n7798), .Q(n13603)
         );
  MUX21X1 U12767 ( .IN1(\mem3[142][30] ), .IN2(n1358), .S(n7798), .Q(n13602)
         );
  MUX21X1 U12768 ( .IN1(\mem3[142][29] ), .IN2(n1336), .S(n7798), .Q(n13601)
         );
  MUX21X1 U12769 ( .IN1(\mem3[142][28] ), .IN2(n1314), .S(n7798), .Q(n13600)
         );
  MUX21X1 U12770 ( .IN1(\mem3[142][27] ), .IN2(n1292), .S(n7798), .Q(n13599)
         );
  MUX21X1 U12771 ( .IN1(\mem3[142][26] ), .IN2(n1270), .S(n7798), .Q(n13598)
         );
  MUX21X1 U12772 ( .IN1(\mem3[142][25] ), .IN2(n1248), .S(n7798), .Q(n13597)
         );
  MUX21X1 U12773 ( .IN1(\mem3[142][24] ), .IN2(n1226), .S(n7798), .Q(n13596)
         );
  AND2X1 U12774 ( .IN1(n7797), .IN2(n7102), .Q(n7798) );
  MUX21X1 U12775 ( .IN1(\mem3[141][31] ), .IN2(n1380), .S(n7799), .Q(n13595)
         );
  MUX21X1 U12776 ( .IN1(\mem3[141][30] ), .IN2(n1358), .S(n7799), .Q(n13594)
         );
  MUX21X1 U12777 ( .IN1(\mem3[141][29] ), .IN2(n1336), .S(n7799), .Q(n13593)
         );
  MUX21X1 U12778 ( .IN1(\mem3[141][28] ), .IN2(n1314), .S(n7799), .Q(n13592)
         );
  MUX21X1 U12779 ( .IN1(\mem3[141][27] ), .IN2(n1292), .S(n7799), .Q(n13591)
         );
  MUX21X1 U12780 ( .IN1(\mem3[141][26] ), .IN2(n1270), .S(n7799), .Q(n13590)
         );
  MUX21X1 U12781 ( .IN1(\mem3[141][25] ), .IN2(n1248), .S(n7799), .Q(n13589)
         );
  MUX21X1 U12782 ( .IN1(\mem3[141][24] ), .IN2(n1226), .S(n7799), .Q(n13588)
         );
  AND2X1 U12783 ( .IN1(n7797), .IN2(n7104), .Q(n7799) );
  MUX21X1 U12784 ( .IN1(\mem3[140][31] ), .IN2(n1380), .S(n7800), .Q(n13587)
         );
  MUX21X1 U12785 ( .IN1(\mem3[140][30] ), .IN2(n1358), .S(n7800), .Q(n13586)
         );
  MUX21X1 U12786 ( .IN1(\mem3[140][29] ), .IN2(n1336), .S(n7800), .Q(n13585)
         );
  MUX21X1 U12787 ( .IN1(\mem3[140][28] ), .IN2(n1314), .S(n7800), .Q(n13584)
         );
  MUX21X1 U12788 ( .IN1(\mem3[140][27] ), .IN2(n1292), .S(n7800), .Q(n13583)
         );
  MUX21X1 U12789 ( .IN1(\mem3[140][26] ), .IN2(n1270), .S(n7800), .Q(n13582)
         );
  MUX21X1 U12790 ( .IN1(\mem3[140][25] ), .IN2(n1248), .S(n7800), .Q(n13581)
         );
  MUX21X1 U12791 ( .IN1(\mem3[140][24] ), .IN2(n1226), .S(n7800), .Q(n13580)
         );
  AND2X1 U12792 ( .IN1(n7797), .IN2(n7106), .Q(n7800) );
  MUX21X1 U12793 ( .IN1(\mem3[139][31] ), .IN2(n1380), .S(n7801), .Q(n13579)
         );
  MUX21X1 U12794 ( .IN1(\mem3[139][30] ), .IN2(n1358), .S(n7801), .Q(n13578)
         );
  MUX21X1 U12795 ( .IN1(\mem3[139][29] ), .IN2(n1336), .S(n7801), .Q(n13577)
         );
  MUX21X1 U12796 ( .IN1(\mem3[139][28] ), .IN2(n1314), .S(n7801), .Q(n13576)
         );
  MUX21X1 U12797 ( .IN1(\mem3[139][27] ), .IN2(n1292), .S(n7801), .Q(n13575)
         );
  MUX21X1 U12798 ( .IN1(\mem3[139][26] ), .IN2(n1270), .S(n7801), .Q(n13574)
         );
  MUX21X1 U12799 ( .IN1(\mem3[139][25] ), .IN2(n1248), .S(n7801), .Q(n13573)
         );
  MUX21X1 U12800 ( .IN1(\mem3[139][24] ), .IN2(n1226), .S(n7801), .Q(n13572)
         );
  AND2X1 U12801 ( .IN1(n7797), .IN2(n7108), .Q(n7801) );
  MUX21X1 U12802 ( .IN1(\mem3[138][31] ), .IN2(n1380), .S(n7802), .Q(n13571)
         );
  MUX21X1 U12803 ( .IN1(\mem3[138][30] ), .IN2(n1358), .S(n7802), .Q(n13570)
         );
  MUX21X1 U12804 ( .IN1(\mem3[138][29] ), .IN2(n1336), .S(n7802), .Q(n13569)
         );
  MUX21X1 U12805 ( .IN1(\mem3[138][28] ), .IN2(n1314), .S(n7802), .Q(n13568)
         );
  MUX21X1 U12806 ( .IN1(\mem3[138][27] ), .IN2(n1292), .S(n7802), .Q(n13567)
         );
  MUX21X1 U12807 ( .IN1(\mem3[138][26] ), .IN2(n1270), .S(n7802), .Q(n13566)
         );
  MUX21X1 U12808 ( .IN1(\mem3[138][25] ), .IN2(n1248), .S(n7802), .Q(n13565)
         );
  MUX21X1 U12809 ( .IN1(\mem3[138][24] ), .IN2(n1226), .S(n7802), .Q(n13564)
         );
  AND2X1 U12810 ( .IN1(n7797), .IN2(n7110), .Q(n7802) );
  MUX21X1 U12811 ( .IN1(\mem3[137][31] ), .IN2(n1380), .S(n7803), .Q(n13563)
         );
  MUX21X1 U12812 ( .IN1(\mem3[137][30] ), .IN2(n1358), .S(n7803), .Q(n13562)
         );
  MUX21X1 U12813 ( .IN1(\mem3[137][29] ), .IN2(n1336), .S(n7803), .Q(n13561)
         );
  MUX21X1 U12814 ( .IN1(\mem3[137][28] ), .IN2(n1314), .S(n7803), .Q(n13560)
         );
  MUX21X1 U12815 ( .IN1(\mem3[137][27] ), .IN2(n1292), .S(n7803), .Q(n13559)
         );
  MUX21X1 U12816 ( .IN1(\mem3[137][26] ), .IN2(n1270), .S(n7803), .Q(n13558)
         );
  MUX21X1 U12817 ( .IN1(\mem3[137][25] ), .IN2(n1248), .S(n7803), .Q(n13557)
         );
  MUX21X1 U12818 ( .IN1(\mem3[137][24] ), .IN2(n1226), .S(n7803), .Q(n13556)
         );
  AND2X1 U12819 ( .IN1(n7797), .IN2(n7112), .Q(n7803) );
  MUX21X1 U12820 ( .IN1(\mem3[136][31] ), .IN2(n1380), .S(n7804), .Q(n13555)
         );
  MUX21X1 U12821 ( .IN1(\mem3[136][30] ), .IN2(n1358), .S(n7804), .Q(n13554)
         );
  MUX21X1 U12822 ( .IN1(\mem3[136][29] ), .IN2(n1336), .S(n7804), .Q(n13553)
         );
  MUX21X1 U12823 ( .IN1(\mem3[136][28] ), .IN2(n1314), .S(n7804), .Q(n13552)
         );
  MUX21X1 U12824 ( .IN1(\mem3[136][27] ), .IN2(n1292), .S(n7804), .Q(n13551)
         );
  MUX21X1 U12825 ( .IN1(\mem3[136][26] ), .IN2(n1270), .S(n7804), .Q(n13550)
         );
  MUX21X1 U12826 ( .IN1(\mem3[136][25] ), .IN2(n1248), .S(n7804), .Q(n13549)
         );
  MUX21X1 U12827 ( .IN1(\mem3[136][24] ), .IN2(n1226), .S(n7804), .Q(n13548)
         );
  AND2X1 U12828 ( .IN1(n7797), .IN2(n7114), .Q(n7804) );
  MUX21X1 U12829 ( .IN1(\mem3[135][31] ), .IN2(n1381), .S(n7805), .Q(n13547)
         );
  MUX21X1 U12830 ( .IN1(\mem3[135][30] ), .IN2(n1359), .S(n7805), .Q(n13546)
         );
  MUX21X1 U12831 ( .IN1(\mem3[135][29] ), .IN2(n1337), .S(n7805), .Q(n13545)
         );
  MUX21X1 U12832 ( .IN1(\mem3[135][28] ), .IN2(n1315), .S(n7805), .Q(n13544)
         );
  MUX21X1 U12833 ( .IN1(\mem3[135][27] ), .IN2(n1293), .S(n7805), .Q(n13543)
         );
  MUX21X1 U12834 ( .IN1(\mem3[135][26] ), .IN2(n1271), .S(n7805), .Q(n13542)
         );
  MUX21X1 U12835 ( .IN1(\mem3[135][25] ), .IN2(n1249), .S(n7805), .Q(n13541)
         );
  MUX21X1 U12836 ( .IN1(\mem3[135][24] ), .IN2(n1227), .S(n7805), .Q(n13540)
         );
  AND2X1 U12837 ( .IN1(n7797), .IN2(n7116), .Q(n7805) );
  MUX21X1 U12838 ( .IN1(\mem3[134][31] ), .IN2(n1381), .S(n7806), .Q(n13539)
         );
  MUX21X1 U12839 ( .IN1(\mem3[134][30] ), .IN2(n1359), .S(n7806), .Q(n13538)
         );
  MUX21X1 U12840 ( .IN1(\mem3[134][29] ), .IN2(n1337), .S(n7806), .Q(n13537)
         );
  MUX21X1 U12841 ( .IN1(\mem3[134][28] ), .IN2(n1315), .S(n7806), .Q(n13536)
         );
  MUX21X1 U12842 ( .IN1(\mem3[134][27] ), .IN2(n1293), .S(n7806), .Q(n13535)
         );
  MUX21X1 U12843 ( .IN1(\mem3[134][26] ), .IN2(n1271), .S(n7806), .Q(n13534)
         );
  MUX21X1 U12844 ( .IN1(\mem3[134][25] ), .IN2(n1249), .S(n7806), .Q(n13533)
         );
  MUX21X1 U12845 ( .IN1(\mem3[134][24] ), .IN2(n1227), .S(n7806), .Q(n13532)
         );
  AND2X1 U12846 ( .IN1(n7797), .IN2(n7118), .Q(n7806) );
  MUX21X1 U12847 ( .IN1(\mem3[133][31] ), .IN2(n1381), .S(n7807), .Q(n13531)
         );
  MUX21X1 U12848 ( .IN1(\mem3[133][30] ), .IN2(n1359), .S(n7807), .Q(n13530)
         );
  MUX21X1 U12849 ( .IN1(\mem3[133][29] ), .IN2(n1337), .S(n7807), .Q(n13529)
         );
  MUX21X1 U12850 ( .IN1(\mem3[133][28] ), .IN2(n1315), .S(n7807), .Q(n13528)
         );
  MUX21X1 U12851 ( .IN1(\mem3[133][27] ), .IN2(n1293), .S(n7807), .Q(n13527)
         );
  MUX21X1 U12852 ( .IN1(\mem3[133][26] ), .IN2(n1271), .S(n7807), .Q(n13526)
         );
  MUX21X1 U12853 ( .IN1(\mem3[133][25] ), .IN2(n1249), .S(n7807), .Q(n13525)
         );
  MUX21X1 U12854 ( .IN1(\mem3[133][24] ), .IN2(n1227), .S(n7807), .Q(n13524)
         );
  AND2X1 U12855 ( .IN1(n7797), .IN2(n7120), .Q(n7807) );
  MUX21X1 U12856 ( .IN1(\mem3[132][31] ), .IN2(n1381), .S(n7808), .Q(n13523)
         );
  MUX21X1 U12857 ( .IN1(\mem3[132][30] ), .IN2(n1359), .S(n7808), .Q(n13522)
         );
  MUX21X1 U12858 ( .IN1(\mem3[132][29] ), .IN2(n1337), .S(n7808), .Q(n13521)
         );
  MUX21X1 U12859 ( .IN1(\mem3[132][28] ), .IN2(n1315), .S(n7808), .Q(n13520)
         );
  MUX21X1 U12860 ( .IN1(\mem3[132][27] ), .IN2(n1293), .S(n7808), .Q(n13519)
         );
  MUX21X1 U12861 ( .IN1(\mem3[132][26] ), .IN2(n1271), .S(n7808), .Q(n13518)
         );
  MUX21X1 U12862 ( .IN1(\mem3[132][25] ), .IN2(n1249), .S(n7808), .Q(n13517)
         );
  MUX21X1 U12863 ( .IN1(\mem3[132][24] ), .IN2(n1227), .S(n7808), .Q(n13516)
         );
  AND2X1 U12864 ( .IN1(n7797), .IN2(n7122), .Q(n7808) );
  MUX21X1 U12865 ( .IN1(\mem3[131][31] ), .IN2(n1381), .S(n7809), .Q(n13515)
         );
  MUX21X1 U12866 ( .IN1(\mem3[131][30] ), .IN2(n1359), .S(n7809), .Q(n13514)
         );
  MUX21X1 U12867 ( .IN1(\mem3[131][29] ), .IN2(n1337), .S(n7809), .Q(n13513)
         );
  MUX21X1 U12868 ( .IN1(\mem3[131][28] ), .IN2(n1315), .S(n7809), .Q(n13512)
         );
  MUX21X1 U12869 ( .IN1(\mem3[131][27] ), .IN2(n1293), .S(n7809), .Q(n13511)
         );
  MUX21X1 U12870 ( .IN1(\mem3[131][26] ), .IN2(n1271), .S(n7809), .Q(n13510)
         );
  MUX21X1 U12871 ( .IN1(\mem3[131][25] ), .IN2(n1249), .S(n7809), .Q(n13509)
         );
  MUX21X1 U12872 ( .IN1(\mem3[131][24] ), .IN2(n1227), .S(n7809), .Q(n13508)
         );
  AND2X1 U12873 ( .IN1(n7797), .IN2(n7124), .Q(n7809) );
  MUX21X1 U12874 ( .IN1(\mem3[130][31] ), .IN2(n1381), .S(n7810), .Q(n13507)
         );
  MUX21X1 U12875 ( .IN1(\mem3[130][30] ), .IN2(n1359), .S(n7810), .Q(n13506)
         );
  MUX21X1 U12876 ( .IN1(\mem3[130][29] ), .IN2(n1337), .S(n7810), .Q(n13505)
         );
  MUX21X1 U12877 ( .IN1(\mem3[130][28] ), .IN2(n1315), .S(n7810), .Q(n13504)
         );
  MUX21X1 U12878 ( .IN1(\mem3[130][27] ), .IN2(n1293), .S(n7810), .Q(n13503)
         );
  MUX21X1 U12879 ( .IN1(\mem3[130][26] ), .IN2(n1271), .S(n7810), .Q(n13502)
         );
  MUX21X1 U12880 ( .IN1(\mem3[130][25] ), .IN2(n1249), .S(n7810), .Q(n13501)
         );
  MUX21X1 U12881 ( .IN1(\mem3[130][24] ), .IN2(n1227), .S(n7810), .Q(n13500)
         );
  AND2X1 U12882 ( .IN1(n7797), .IN2(n7126), .Q(n7810) );
  MUX21X1 U12883 ( .IN1(\mem3[129][31] ), .IN2(n1381), .S(n7811), .Q(n13499)
         );
  MUX21X1 U12884 ( .IN1(\mem3[129][30] ), .IN2(n1359), .S(n7811), .Q(n13498)
         );
  MUX21X1 U12885 ( .IN1(\mem3[129][29] ), .IN2(n1337), .S(n7811), .Q(n13497)
         );
  MUX21X1 U12886 ( .IN1(\mem3[129][28] ), .IN2(n1315), .S(n7811), .Q(n13496)
         );
  MUX21X1 U12887 ( .IN1(\mem3[129][27] ), .IN2(n1293), .S(n7811), .Q(n13495)
         );
  MUX21X1 U12888 ( .IN1(\mem3[129][26] ), .IN2(n1271), .S(n7811), .Q(n13494)
         );
  MUX21X1 U12889 ( .IN1(\mem3[129][25] ), .IN2(n1249), .S(n7811), .Q(n13493)
         );
  MUX21X1 U12890 ( .IN1(\mem3[129][24] ), .IN2(n1227), .S(n7811), .Q(n13492)
         );
  AND2X1 U12891 ( .IN1(n7797), .IN2(n7128), .Q(n7811) );
  MUX21X1 U12892 ( .IN1(\mem3[128][31] ), .IN2(n1381), .S(n7812), .Q(n13491)
         );
  MUX21X1 U12893 ( .IN1(\mem3[128][30] ), .IN2(n1359), .S(n7812), .Q(n13490)
         );
  MUX21X1 U12894 ( .IN1(\mem3[128][29] ), .IN2(n1337), .S(n7812), .Q(n13489)
         );
  MUX21X1 U12895 ( .IN1(\mem3[128][28] ), .IN2(n1315), .S(n7812), .Q(n13488)
         );
  MUX21X1 U12896 ( .IN1(\mem3[128][27] ), .IN2(n1293), .S(n7812), .Q(n13487)
         );
  MUX21X1 U12897 ( .IN1(\mem3[128][26] ), .IN2(n1271), .S(n7812), .Q(n13486)
         );
  MUX21X1 U12898 ( .IN1(\mem3[128][25] ), .IN2(n1249), .S(n7812), .Q(n13485)
         );
  MUX21X1 U12899 ( .IN1(\mem3[128][24] ), .IN2(n1227), .S(n7812), .Q(n13484)
         );
  AND2X1 U12900 ( .IN1(n7797), .IN2(n7130), .Q(n7812) );
  AND2X1 U12901 ( .IN1(n7693), .IN2(n7258), .Q(n7797) );
  MUX21X1 U12902 ( .IN1(\mem3[127][31] ), .IN2(n1381), .S(n7813), .Q(n13483)
         );
  MUX21X1 U12903 ( .IN1(\mem3[127][30] ), .IN2(n1359), .S(n7813), .Q(n13482)
         );
  MUX21X1 U12904 ( .IN1(\mem3[127][29] ), .IN2(n1337), .S(n7813), .Q(n13481)
         );
  MUX21X1 U12905 ( .IN1(\mem3[127][28] ), .IN2(n1315), .S(n7813), .Q(n13480)
         );
  MUX21X1 U12906 ( .IN1(\mem3[127][27] ), .IN2(n1293), .S(n7813), .Q(n13479)
         );
  MUX21X1 U12907 ( .IN1(\mem3[127][26] ), .IN2(n1271), .S(n7813), .Q(n13478)
         );
  MUX21X1 U12908 ( .IN1(\mem3[127][25] ), .IN2(n1249), .S(n7813), .Q(n13477)
         );
  MUX21X1 U12909 ( .IN1(\mem3[127][24] ), .IN2(n1227), .S(n7813), .Q(n13476)
         );
  AND2X1 U12910 ( .IN1(n7814), .IN2(n7099), .Q(n7813) );
  MUX21X1 U12911 ( .IN1(\mem3[126][31] ), .IN2(n1381), .S(n7815), .Q(n13475)
         );
  MUX21X1 U12912 ( .IN1(\mem3[126][30] ), .IN2(n1359), .S(n7815), .Q(n13474)
         );
  MUX21X1 U12913 ( .IN1(\mem3[126][29] ), .IN2(n1337), .S(n7815), .Q(n13473)
         );
  MUX21X1 U12914 ( .IN1(\mem3[126][28] ), .IN2(n1315), .S(n7815), .Q(n13472)
         );
  MUX21X1 U12915 ( .IN1(\mem3[126][27] ), .IN2(n1293), .S(n7815), .Q(n13471)
         );
  MUX21X1 U12916 ( .IN1(\mem3[126][26] ), .IN2(n1271), .S(n7815), .Q(n13470)
         );
  MUX21X1 U12917 ( .IN1(\mem3[126][25] ), .IN2(n1249), .S(n7815), .Q(n13469)
         );
  MUX21X1 U12918 ( .IN1(\mem3[126][24] ), .IN2(n1227), .S(n7815), .Q(n13468)
         );
  AND2X1 U12919 ( .IN1(n7814), .IN2(n7102), .Q(n7815) );
  MUX21X1 U12920 ( .IN1(\mem3[125][31] ), .IN2(n1381), .S(n7816), .Q(n13467)
         );
  MUX21X1 U12921 ( .IN1(\mem3[125][30] ), .IN2(n1359), .S(n7816), .Q(n13466)
         );
  MUX21X1 U12922 ( .IN1(\mem3[125][29] ), .IN2(n1337), .S(n7816), .Q(n13465)
         );
  MUX21X1 U12923 ( .IN1(\mem3[125][28] ), .IN2(n1315), .S(n7816), .Q(n13464)
         );
  MUX21X1 U12924 ( .IN1(\mem3[125][27] ), .IN2(n1293), .S(n7816), .Q(n13463)
         );
  MUX21X1 U12925 ( .IN1(\mem3[125][26] ), .IN2(n1271), .S(n7816), .Q(n13462)
         );
  MUX21X1 U12926 ( .IN1(\mem3[125][25] ), .IN2(n1249), .S(n7816), .Q(n13461)
         );
  MUX21X1 U12927 ( .IN1(\mem3[125][24] ), .IN2(n1227), .S(n7816), .Q(n13460)
         );
  AND2X1 U12928 ( .IN1(n7814), .IN2(n7104), .Q(n7816) );
  MUX21X1 U12929 ( .IN1(\mem3[124][31] ), .IN2(n1381), .S(n7817), .Q(n13459)
         );
  MUX21X1 U12930 ( .IN1(\mem3[124][30] ), .IN2(n1359), .S(n7817), .Q(n13458)
         );
  MUX21X1 U12931 ( .IN1(\mem3[124][29] ), .IN2(n1337), .S(n7817), .Q(n13457)
         );
  MUX21X1 U12932 ( .IN1(\mem3[124][28] ), .IN2(n1315), .S(n7817), .Q(n13456)
         );
  MUX21X1 U12933 ( .IN1(\mem3[124][27] ), .IN2(n1293), .S(n7817), .Q(n13455)
         );
  MUX21X1 U12934 ( .IN1(\mem3[124][26] ), .IN2(n1271), .S(n7817), .Q(n13454)
         );
  MUX21X1 U12935 ( .IN1(\mem3[124][25] ), .IN2(n1249), .S(n7817), .Q(n13453)
         );
  MUX21X1 U12936 ( .IN1(\mem3[124][24] ), .IN2(n1227), .S(n7817), .Q(n13452)
         );
  AND2X1 U12937 ( .IN1(n7814), .IN2(n7106), .Q(n7817) );
  MUX21X1 U12938 ( .IN1(\mem3[123][31] ), .IN2(n1382), .S(n7818), .Q(n13451)
         );
  MUX21X1 U12939 ( .IN1(\mem3[123][30] ), .IN2(n1360), .S(n7818), .Q(n13450)
         );
  MUX21X1 U12940 ( .IN1(\mem3[123][29] ), .IN2(n1338), .S(n7818), .Q(n13449)
         );
  MUX21X1 U12941 ( .IN1(\mem3[123][28] ), .IN2(n1316), .S(n7818), .Q(n13448)
         );
  MUX21X1 U12942 ( .IN1(\mem3[123][27] ), .IN2(n1294), .S(n7818), .Q(n13447)
         );
  MUX21X1 U12943 ( .IN1(\mem3[123][26] ), .IN2(n1272), .S(n7818), .Q(n13446)
         );
  MUX21X1 U12944 ( .IN1(\mem3[123][25] ), .IN2(n1250), .S(n7818), .Q(n13445)
         );
  MUX21X1 U12945 ( .IN1(\mem3[123][24] ), .IN2(n1228), .S(n7818), .Q(n13444)
         );
  AND2X1 U12946 ( .IN1(n7814), .IN2(n7108), .Q(n7818) );
  MUX21X1 U12947 ( .IN1(\mem3[122][31] ), .IN2(n1382), .S(n7819), .Q(n13443)
         );
  MUX21X1 U12948 ( .IN1(\mem3[122][30] ), .IN2(n1360), .S(n7819), .Q(n13442)
         );
  MUX21X1 U12949 ( .IN1(\mem3[122][29] ), .IN2(n1338), .S(n7819), .Q(n13441)
         );
  MUX21X1 U12950 ( .IN1(\mem3[122][28] ), .IN2(n1316), .S(n7819), .Q(n13440)
         );
  MUX21X1 U12951 ( .IN1(\mem3[122][27] ), .IN2(n1294), .S(n7819), .Q(n13439)
         );
  MUX21X1 U12952 ( .IN1(\mem3[122][26] ), .IN2(n1272), .S(n7819), .Q(n13438)
         );
  MUX21X1 U12953 ( .IN1(\mem3[122][25] ), .IN2(n1250), .S(n7819), .Q(n13437)
         );
  MUX21X1 U12954 ( .IN1(\mem3[122][24] ), .IN2(n1228), .S(n7819), .Q(n13436)
         );
  AND2X1 U12955 ( .IN1(n7814), .IN2(n7110), .Q(n7819) );
  MUX21X1 U12956 ( .IN1(\mem3[121][31] ), .IN2(n1382), .S(n7820), .Q(n13435)
         );
  MUX21X1 U12957 ( .IN1(\mem3[121][30] ), .IN2(n1360), .S(n7820), .Q(n13434)
         );
  MUX21X1 U12958 ( .IN1(\mem3[121][29] ), .IN2(n1338), .S(n7820), .Q(n13433)
         );
  MUX21X1 U12959 ( .IN1(\mem3[121][28] ), .IN2(n1316), .S(n7820), .Q(n13432)
         );
  MUX21X1 U12960 ( .IN1(\mem3[121][27] ), .IN2(n1294), .S(n7820), .Q(n13431)
         );
  MUX21X1 U12961 ( .IN1(\mem3[121][26] ), .IN2(n1272), .S(n7820), .Q(n13430)
         );
  MUX21X1 U12962 ( .IN1(\mem3[121][25] ), .IN2(n1250), .S(n7820), .Q(n13429)
         );
  MUX21X1 U12963 ( .IN1(\mem3[121][24] ), .IN2(n1228), .S(n7820), .Q(n13428)
         );
  AND2X1 U12964 ( .IN1(n7814), .IN2(n7112), .Q(n7820) );
  MUX21X1 U12965 ( .IN1(\mem3[120][31] ), .IN2(n1382), .S(n7821), .Q(n13427)
         );
  MUX21X1 U12966 ( .IN1(\mem3[120][30] ), .IN2(n1360), .S(n7821), .Q(n13426)
         );
  MUX21X1 U12967 ( .IN1(\mem3[120][29] ), .IN2(n1338), .S(n7821), .Q(n13425)
         );
  MUX21X1 U12968 ( .IN1(\mem3[120][28] ), .IN2(n1316), .S(n7821), .Q(n13424)
         );
  MUX21X1 U12969 ( .IN1(\mem3[120][27] ), .IN2(n1294), .S(n7821), .Q(n13423)
         );
  MUX21X1 U12970 ( .IN1(\mem3[120][26] ), .IN2(n1272), .S(n7821), .Q(n13422)
         );
  MUX21X1 U12971 ( .IN1(\mem3[120][25] ), .IN2(n1250), .S(n7821), .Q(n13421)
         );
  MUX21X1 U12972 ( .IN1(\mem3[120][24] ), .IN2(n1228), .S(n7821), .Q(n13420)
         );
  AND2X1 U12973 ( .IN1(n7814), .IN2(n7114), .Q(n7821) );
  MUX21X1 U12974 ( .IN1(\mem3[119][31] ), .IN2(n1382), .S(n7822), .Q(n13419)
         );
  MUX21X1 U12975 ( .IN1(\mem3[119][30] ), .IN2(n1360), .S(n7822), .Q(n13418)
         );
  MUX21X1 U12976 ( .IN1(\mem3[119][29] ), .IN2(n1338), .S(n7822), .Q(n13417)
         );
  MUX21X1 U12977 ( .IN1(\mem3[119][28] ), .IN2(n1316), .S(n7822), .Q(n13416)
         );
  MUX21X1 U12978 ( .IN1(\mem3[119][27] ), .IN2(n1294), .S(n7822), .Q(n13415)
         );
  MUX21X1 U12979 ( .IN1(\mem3[119][26] ), .IN2(n1272), .S(n7822), .Q(n13414)
         );
  MUX21X1 U12980 ( .IN1(\mem3[119][25] ), .IN2(n1250), .S(n7822), .Q(n13413)
         );
  MUX21X1 U12981 ( .IN1(\mem3[119][24] ), .IN2(n1228), .S(n7822), .Q(n13412)
         );
  AND2X1 U12982 ( .IN1(n7814), .IN2(n7116), .Q(n7822) );
  MUX21X1 U12983 ( .IN1(\mem3[118][31] ), .IN2(n1382), .S(n7823), .Q(n13411)
         );
  MUX21X1 U12984 ( .IN1(\mem3[118][30] ), .IN2(n1360), .S(n7823), .Q(n13410)
         );
  MUX21X1 U12985 ( .IN1(\mem3[118][29] ), .IN2(n1338), .S(n7823), .Q(n13409)
         );
  MUX21X1 U12986 ( .IN1(\mem3[118][28] ), .IN2(n1316), .S(n7823), .Q(n13408)
         );
  MUX21X1 U12987 ( .IN1(\mem3[118][27] ), .IN2(n1294), .S(n7823), .Q(n13407)
         );
  MUX21X1 U12988 ( .IN1(\mem3[118][26] ), .IN2(n1272), .S(n7823), .Q(n13406)
         );
  MUX21X1 U12989 ( .IN1(\mem3[118][25] ), .IN2(n1250), .S(n7823), .Q(n13405)
         );
  MUX21X1 U12990 ( .IN1(\mem3[118][24] ), .IN2(n1228), .S(n7823), .Q(n13404)
         );
  AND2X1 U12991 ( .IN1(n7814), .IN2(n7118), .Q(n7823) );
  MUX21X1 U12992 ( .IN1(\mem3[117][31] ), .IN2(n1382), .S(n7824), .Q(n13403)
         );
  MUX21X1 U12993 ( .IN1(\mem3[117][30] ), .IN2(n1360), .S(n7824), .Q(n13402)
         );
  MUX21X1 U12994 ( .IN1(\mem3[117][29] ), .IN2(n1338), .S(n7824), .Q(n13401)
         );
  MUX21X1 U12995 ( .IN1(\mem3[117][28] ), .IN2(n1316), .S(n7824), .Q(n13400)
         );
  MUX21X1 U12996 ( .IN1(\mem3[117][27] ), .IN2(n1294), .S(n7824), .Q(n13399)
         );
  MUX21X1 U12997 ( .IN1(\mem3[117][26] ), .IN2(n1272), .S(n7824), .Q(n13398)
         );
  MUX21X1 U12998 ( .IN1(\mem3[117][25] ), .IN2(n1250), .S(n7824), .Q(n13397)
         );
  MUX21X1 U12999 ( .IN1(\mem3[117][24] ), .IN2(n1228), .S(n7824), .Q(n13396)
         );
  AND2X1 U13000 ( .IN1(n7814), .IN2(n7120), .Q(n7824) );
  MUX21X1 U13001 ( .IN1(\mem3[116][31] ), .IN2(n1382), .S(n7825), .Q(n13395)
         );
  MUX21X1 U13002 ( .IN1(\mem3[116][30] ), .IN2(n1360), .S(n7825), .Q(n13394)
         );
  MUX21X1 U13003 ( .IN1(\mem3[116][29] ), .IN2(n1338), .S(n7825), .Q(n13393)
         );
  MUX21X1 U13004 ( .IN1(\mem3[116][28] ), .IN2(n1316), .S(n7825), .Q(n13392)
         );
  MUX21X1 U13005 ( .IN1(\mem3[116][27] ), .IN2(n1294), .S(n7825), .Q(n13391)
         );
  MUX21X1 U13006 ( .IN1(\mem3[116][26] ), .IN2(n1272), .S(n7825), .Q(n13390)
         );
  MUX21X1 U13007 ( .IN1(\mem3[116][25] ), .IN2(n1250), .S(n7825), .Q(n13389)
         );
  MUX21X1 U13008 ( .IN1(\mem3[116][24] ), .IN2(n1228), .S(n7825), .Q(n13388)
         );
  AND2X1 U13009 ( .IN1(n7814), .IN2(n7122), .Q(n7825) );
  MUX21X1 U13010 ( .IN1(\mem3[115][31] ), .IN2(n1382), .S(n7826), .Q(n13387)
         );
  MUX21X1 U13011 ( .IN1(\mem3[115][30] ), .IN2(n1360), .S(n7826), .Q(n13386)
         );
  MUX21X1 U13012 ( .IN1(\mem3[115][29] ), .IN2(n1338), .S(n7826), .Q(n13385)
         );
  MUX21X1 U13013 ( .IN1(\mem3[115][28] ), .IN2(n1316), .S(n7826), .Q(n13384)
         );
  MUX21X1 U13014 ( .IN1(\mem3[115][27] ), .IN2(n1294), .S(n7826), .Q(n13383)
         );
  MUX21X1 U13015 ( .IN1(\mem3[115][26] ), .IN2(n1272), .S(n7826), .Q(n13382)
         );
  MUX21X1 U13016 ( .IN1(\mem3[115][25] ), .IN2(n1250), .S(n7826), .Q(n13381)
         );
  MUX21X1 U13017 ( .IN1(\mem3[115][24] ), .IN2(n1228), .S(n7826), .Q(n13380)
         );
  AND2X1 U13018 ( .IN1(n7814), .IN2(n7124), .Q(n7826) );
  MUX21X1 U13019 ( .IN1(\mem3[114][31] ), .IN2(n1382), .S(n7827), .Q(n13379)
         );
  MUX21X1 U13020 ( .IN1(\mem3[114][30] ), .IN2(n1360), .S(n7827), .Q(n13378)
         );
  MUX21X1 U13021 ( .IN1(\mem3[114][29] ), .IN2(n1338), .S(n7827), .Q(n13377)
         );
  MUX21X1 U13022 ( .IN1(\mem3[114][28] ), .IN2(n1316), .S(n7827), .Q(n13376)
         );
  MUX21X1 U13023 ( .IN1(\mem3[114][27] ), .IN2(n1294), .S(n7827), .Q(n13375)
         );
  MUX21X1 U13024 ( .IN1(\mem3[114][26] ), .IN2(n1272), .S(n7827), .Q(n13374)
         );
  MUX21X1 U13025 ( .IN1(\mem3[114][25] ), .IN2(n1250), .S(n7827), .Q(n13373)
         );
  MUX21X1 U13026 ( .IN1(\mem3[114][24] ), .IN2(n1228), .S(n7827), .Q(n13372)
         );
  AND2X1 U13027 ( .IN1(n7814), .IN2(n7126), .Q(n7827) );
  MUX21X1 U13028 ( .IN1(\mem3[113][31] ), .IN2(n1382), .S(n7828), .Q(n13371)
         );
  MUX21X1 U13029 ( .IN1(\mem3[113][30] ), .IN2(n1360), .S(n7828), .Q(n13370)
         );
  MUX21X1 U13030 ( .IN1(\mem3[113][29] ), .IN2(n1338), .S(n7828), .Q(n13369)
         );
  MUX21X1 U13031 ( .IN1(\mem3[113][28] ), .IN2(n1316), .S(n7828), .Q(n13368)
         );
  MUX21X1 U13032 ( .IN1(\mem3[113][27] ), .IN2(n1294), .S(n7828), .Q(n13367)
         );
  MUX21X1 U13033 ( .IN1(\mem3[113][26] ), .IN2(n1272), .S(n7828), .Q(n13366)
         );
  MUX21X1 U13034 ( .IN1(\mem3[113][25] ), .IN2(n1250), .S(n7828), .Q(n13365)
         );
  MUX21X1 U13035 ( .IN1(\mem3[113][24] ), .IN2(n1228), .S(n7828), .Q(n13364)
         );
  AND2X1 U13036 ( .IN1(n7814), .IN2(n7128), .Q(n7828) );
  MUX21X1 U13037 ( .IN1(\mem3[112][31] ), .IN2(n1382), .S(n7829), .Q(n13363)
         );
  MUX21X1 U13038 ( .IN1(\mem3[112][30] ), .IN2(n1360), .S(n7829), .Q(n13362)
         );
  MUX21X1 U13039 ( .IN1(\mem3[112][29] ), .IN2(n1338), .S(n7829), .Q(n13361)
         );
  MUX21X1 U13040 ( .IN1(\mem3[112][28] ), .IN2(n1316), .S(n7829), .Q(n13360)
         );
  MUX21X1 U13041 ( .IN1(\mem3[112][27] ), .IN2(n1294), .S(n7829), .Q(n13359)
         );
  MUX21X1 U13042 ( .IN1(\mem3[112][26] ), .IN2(n1272), .S(n7829), .Q(n13358)
         );
  MUX21X1 U13043 ( .IN1(\mem3[112][25] ), .IN2(n1250), .S(n7829), .Q(n13357)
         );
  MUX21X1 U13044 ( .IN1(\mem3[112][24] ), .IN2(n1228), .S(n7829), .Q(n13356)
         );
  AND2X1 U13045 ( .IN1(n7814), .IN2(n7130), .Q(n7829) );
  AND2X1 U13046 ( .IN1(n7693), .IN2(n7276), .Q(n7814) );
  MUX21X1 U13047 ( .IN1(\mem3[111][31] ), .IN2(n1383), .S(n7830), .Q(n13355)
         );
  MUX21X1 U13048 ( .IN1(\mem3[111][30] ), .IN2(n1361), .S(n7830), .Q(n13354)
         );
  MUX21X1 U13049 ( .IN1(\mem3[111][29] ), .IN2(n1339), .S(n7830), .Q(n13353)
         );
  MUX21X1 U13050 ( .IN1(\mem3[111][28] ), .IN2(n1317), .S(n7830), .Q(n13352)
         );
  MUX21X1 U13051 ( .IN1(\mem3[111][27] ), .IN2(n1295), .S(n7830), .Q(n13351)
         );
  MUX21X1 U13052 ( .IN1(\mem3[111][26] ), .IN2(n1273), .S(n7830), .Q(n13350)
         );
  MUX21X1 U13053 ( .IN1(\mem3[111][25] ), .IN2(n1251), .S(n7830), .Q(n13349)
         );
  MUX21X1 U13054 ( .IN1(\mem3[111][24] ), .IN2(n1229), .S(n7830), .Q(n13348)
         );
  AND2X1 U13055 ( .IN1(n7831), .IN2(n7099), .Q(n7830) );
  MUX21X1 U13056 ( .IN1(\mem3[110][31] ), .IN2(n1383), .S(n7832), .Q(n13347)
         );
  MUX21X1 U13057 ( .IN1(\mem3[110][30] ), .IN2(n1361), .S(n7832), .Q(n13346)
         );
  MUX21X1 U13058 ( .IN1(\mem3[110][29] ), .IN2(n1339), .S(n7832), .Q(n13345)
         );
  MUX21X1 U13059 ( .IN1(\mem3[110][28] ), .IN2(n1317), .S(n7832), .Q(n13344)
         );
  MUX21X1 U13060 ( .IN1(\mem3[110][27] ), .IN2(n1295), .S(n7832), .Q(n13343)
         );
  MUX21X1 U13061 ( .IN1(\mem3[110][26] ), .IN2(n1273), .S(n7832), .Q(n13342)
         );
  MUX21X1 U13062 ( .IN1(\mem3[110][25] ), .IN2(n1251), .S(n7832), .Q(n13341)
         );
  MUX21X1 U13063 ( .IN1(\mem3[110][24] ), .IN2(n1229), .S(n7832), .Q(n13340)
         );
  AND2X1 U13064 ( .IN1(n7831), .IN2(n7102), .Q(n7832) );
  MUX21X1 U13065 ( .IN1(\mem3[109][31] ), .IN2(n1383), .S(n7833), .Q(n13339)
         );
  MUX21X1 U13066 ( .IN1(\mem3[109][30] ), .IN2(n1361), .S(n7833), .Q(n13338)
         );
  MUX21X1 U13067 ( .IN1(\mem3[109][29] ), .IN2(n1339), .S(n7833), .Q(n13337)
         );
  MUX21X1 U13068 ( .IN1(\mem3[109][28] ), .IN2(n1317), .S(n7833), .Q(n13336)
         );
  MUX21X1 U13069 ( .IN1(\mem3[109][27] ), .IN2(n1295), .S(n7833), .Q(n13335)
         );
  MUX21X1 U13070 ( .IN1(\mem3[109][26] ), .IN2(n1273), .S(n7833), .Q(n13334)
         );
  MUX21X1 U13071 ( .IN1(\mem3[109][25] ), .IN2(n1251), .S(n7833), .Q(n13333)
         );
  MUX21X1 U13072 ( .IN1(\mem3[109][24] ), .IN2(n1229), .S(n7833), .Q(n13332)
         );
  AND2X1 U13073 ( .IN1(n7831), .IN2(n7104), .Q(n7833) );
  MUX21X1 U13074 ( .IN1(\mem3[108][31] ), .IN2(n1383), .S(n7834), .Q(n13331)
         );
  MUX21X1 U13075 ( .IN1(\mem3[108][30] ), .IN2(n1361), .S(n7834), .Q(n13330)
         );
  MUX21X1 U13076 ( .IN1(\mem3[108][29] ), .IN2(n1339), .S(n7834), .Q(n13329)
         );
  MUX21X1 U13077 ( .IN1(\mem3[108][28] ), .IN2(n1317), .S(n7834), .Q(n13328)
         );
  MUX21X1 U13078 ( .IN1(\mem3[108][27] ), .IN2(n1295), .S(n7834), .Q(n13327)
         );
  MUX21X1 U13079 ( .IN1(\mem3[108][26] ), .IN2(n1273), .S(n7834), .Q(n13326)
         );
  MUX21X1 U13080 ( .IN1(\mem3[108][25] ), .IN2(n1251), .S(n7834), .Q(n13325)
         );
  MUX21X1 U13081 ( .IN1(\mem3[108][24] ), .IN2(n1229), .S(n7834), .Q(n13324)
         );
  AND2X1 U13082 ( .IN1(n7831), .IN2(n7106), .Q(n7834) );
  MUX21X1 U13083 ( .IN1(\mem3[107][31] ), .IN2(n1383), .S(n7835), .Q(n13323)
         );
  MUX21X1 U13084 ( .IN1(\mem3[107][30] ), .IN2(n1361), .S(n7835), .Q(n13322)
         );
  MUX21X1 U13085 ( .IN1(\mem3[107][29] ), .IN2(n1339), .S(n7835), .Q(n13321)
         );
  MUX21X1 U13086 ( .IN1(\mem3[107][28] ), .IN2(n1317), .S(n7835), .Q(n13320)
         );
  MUX21X1 U13087 ( .IN1(\mem3[107][27] ), .IN2(n1295), .S(n7835), .Q(n13319)
         );
  MUX21X1 U13088 ( .IN1(\mem3[107][26] ), .IN2(n1273), .S(n7835), .Q(n13318)
         );
  MUX21X1 U13089 ( .IN1(\mem3[107][25] ), .IN2(n1251), .S(n7835), .Q(n13317)
         );
  MUX21X1 U13090 ( .IN1(\mem3[107][24] ), .IN2(n1229), .S(n7835), .Q(n13316)
         );
  AND2X1 U13091 ( .IN1(n7831), .IN2(n7108), .Q(n7835) );
  MUX21X1 U13092 ( .IN1(\mem3[106][31] ), .IN2(n1383), .S(n7836), .Q(n13315)
         );
  MUX21X1 U13093 ( .IN1(\mem3[106][30] ), .IN2(n1361), .S(n7836), .Q(n13314)
         );
  MUX21X1 U13094 ( .IN1(\mem3[106][29] ), .IN2(n1339), .S(n7836), .Q(n13313)
         );
  MUX21X1 U13095 ( .IN1(\mem3[106][28] ), .IN2(n1317), .S(n7836), .Q(n13312)
         );
  MUX21X1 U13096 ( .IN1(\mem3[106][27] ), .IN2(n1295), .S(n7836), .Q(n13311)
         );
  MUX21X1 U13097 ( .IN1(\mem3[106][26] ), .IN2(n1273), .S(n7836), .Q(n13310)
         );
  MUX21X1 U13098 ( .IN1(\mem3[106][25] ), .IN2(n1251), .S(n7836), .Q(n13309)
         );
  MUX21X1 U13099 ( .IN1(\mem3[106][24] ), .IN2(n1229), .S(n7836), .Q(n13308)
         );
  AND2X1 U13100 ( .IN1(n7831), .IN2(n7110), .Q(n7836) );
  MUX21X1 U13101 ( .IN1(\mem3[105][31] ), .IN2(n1383), .S(n7837), .Q(n13307)
         );
  MUX21X1 U13102 ( .IN1(\mem3[105][30] ), .IN2(n1361), .S(n7837), .Q(n13306)
         );
  MUX21X1 U13103 ( .IN1(\mem3[105][29] ), .IN2(n1339), .S(n7837), .Q(n13305)
         );
  MUX21X1 U13104 ( .IN1(\mem3[105][28] ), .IN2(n1317), .S(n7837), .Q(n13304)
         );
  MUX21X1 U13105 ( .IN1(\mem3[105][27] ), .IN2(n1295), .S(n7837), .Q(n13303)
         );
  MUX21X1 U13106 ( .IN1(\mem3[105][26] ), .IN2(n1273), .S(n7837), .Q(n13302)
         );
  MUX21X1 U13107 ( .IN1(\mem3[105][25] ), .IN2(n1251), .S(n7837), .Q(n13301)
         );
  MUX21X1 U13108 ( .IN1(\mem3[105][24] ), .IN2(n1229), .S(n7837), .Q(n13300)
         );
  AND2X1 U13109 ( .IN1(n7831), .IN2(n7112), .Q(n7837) );
  MUX21X1 U13110 ( .IN1(\mem3[104][31] ), .IN2(n1383), .S(n7838), .Q(n13299)
         );
  MUX21X1 U13111 ( .IN1(\mem3[104][30] ), .IN2(n1361), .S(n7838), .Q(n13298)
         );
  MUX21X1 U13112 ( .IN1(\mem3[104][29] ), .IN2(n1339), .S(n7838), .Q(n13297)
         );
  MUX21X1 U13113 ( .IN1(\mem3[104][28] ), .IN2(n1317), .S(n7838), .Q(n13296)
         );
  MUX21X1 U13114 ( .IN1(\mem3[104][27] ), .IN2(n1295), .S(n7838), .Q(n13295)
         );
  MUX21X1 U13115 ( .IN1(\mem3[104][26] ), .IN2(n1273), .S(n7838), .Q(n13294)
         );
  MUX21X1 U13116 ( .IN1(\mem3[104][25] ), .IN2(n1251), .S(n7838), .Q(n13293)
         );
  MUX21X1 U13117 ( .IN1(\mem3[104][24] ), .IN2(n1229), .S(n7838), .Q(n13292)
         );
  AND2X1 U13118 ( .IN1(n7831), .IN2(n7114), .Q(n7838) );
  MUX21X1 U13119 ( .IN1(\mem3[103][31] ), .IN2(n1383), .S(n7839), .Q(n13291)
         );
  MUX21X1 U13120 ( .IN1(\mem3[103][30] ), .IN2(n1361), .S(n7839), .Q(n13290)
         );
  MUX21X1 U13121 ( .IN1(\mem3[103][29] ), .IN2(n1339), .S(n7839), .Q(n13289)
         );
  MUX21X1 U13122 ( .IN1(\mem3[103][28] ), .IN2(n1317), .S(n7839), .Q(n13288)
         );
  MUX21X1 U13123 ( .IN1(\mem3[103][27] ), .IN2(n1295), .S(n7839), .Q(n13287)
         );
  MUX21X1 U13124 ( .IN1(\mem3[103][26] ), .IN2(n1273), .S(n7839), .Q(n13286)
         );
  MUX21X1 U13125 ( .IN1(\mem3[103][25] ), .IN2(n1251), .S(n7839), .Q(n13285)
         );
  MUX21X1 U13126 ( .IN1(\mem3[103][24] ), .IN2(n1229), .S(n7839), .Q(n13284)
         );
  AND2X1 U13127 ( .IN1(n7831), .IN2(n7116), .Q(n7839) );
  MUX21X1 U13128 ( .IN1(\mem3[102][31] ), .IN2(n1383), .S(n7840), .Q(n13283)
         );
  MUX21X1 U13129 ( .IN1(\mem3[102][30] ), .IN2(n1361), .S(n7840), .Q(n13282)
         );
  MUX21X1 U13130 ( .IN1(\mem3[102][29] ), .IN2(n1339), .S(n7840), .Q(n13281)
         );
  MUX21X1 U13131 ( .IN1(\mem3[102][28] ), .IN2(n1317), .S(n7840), .Q(n13280)
         );
  MUX21X1 U13132 ( .IN1(\mem3[102][27] ), .IN2(n1295), .S(n7840), .Q(n13279)
         );
  MUX21X1 U13133 ( .IN1(\mem3[102][26] ), .IN2(n1273), .S(n7840), .Q(n13278)
         );
  MUX21X1 U13134 ( .IN1(\mem3[102][25] ), .IN2(n1251), .S(n7840), .Q(n13277)
         );
  MUX21X1 U13135 ( .IN1(\mem3[102][24] ), .IN2(n1229), .S(n7840), .Q(n13276)
         );
  AND2X1 U13136 ( .IN1(n7831), .IN2(n7118), .Q(n7840) );
  MUX21X1 U13137 ( .IN1(\mem3[101][31] ), .IN2(n1383), .S(n7841), .Q(n13275)
         );
  MUX21X1 U13138 ( .IN1(\mem3[101][30] ), .IN2(n1361), .S(n7841), .Q(n13274)
         );
  MUX21X1 U13139 ( .IN1(\mem3[101][29] ), .IN2(n1339), .S(n7841), .Q(n13273)
         );
  MUX21X1 U13140 ( .IN1(\mem3[101][28] ), .IN2(n1317), .S(n7841), .Q(n13272)
         );
  MUX21X1 U13141 ( .IN1(\mem3[101][27] ), .IN2(n1295), .S(n7841), .Q(n13271)
         );
  MUX21X1 U13142 ( .IN1(\mem3[101][26] ), .IN2(n1273), .S(n7841), .Q(n13270)
         );
  MUX21X1 U13143 ( .IN1(\mem3[101][25] ), .IN2(n1251), .S(n7841), .Q(n13269)
         );
  MUX21X1 U13144 ( .IN1(\mem3[101][24] ), .IN2(n1229), .S(n7841), .Q(n13268)
         );
  AND2X1 U13145 ( .IN1(n7831), .IN2(n7120), .Q(n7841) );
  MUX21X1 U13146 ( .IN1(\mem3[100][31] ), .IN2(n1383), .S(n7842), .Q(n13267)
         );
  MUX21X1 U13147 ( .IN1(\mem3[100][30] ), .IN2(n1361), .S(n7842), .Q(n13266)
         );
  MUX21X1 U13148 ( .IN1(\mem3[100][29] ), .IN2(n1339), .S(n7842), .Q(n13265)
         );
  MUX21X1 U13149 ( .IN1(\mem3[100][28] ), .IN2(n1317), .S(n7842), .Q(n13264)
         );
  MUX21X1 U13150 ( .IN1(\mem3[100][27] ), .IN2(n1295), .S(n7842), .Q(n13263)
         );
  MUX21X1 U13151 ( .IN1(\mem3[100][26] ), .IN2(n1273), .S(n7842), .Q(n13262)
         );
  MUX21X1 U13152 ( .IN1(\mem3[100][25] ), .IN2(n1251), .S(n7842), .Q(n13261)
         );
  MUX21X1 U13153 ( .IN1(\mem3[100][24] ), .IN2(n1229), .S(n7842), .Q(n13260)
         );
  AND2X1 U13154 ( .IN1(n7831), .IN2(n7122), .Q(n7842) );
  MUX21X1 U13155 ( .IN1(\mem3[99][31] ), .IN2(n1384), .S(n7843), .Q(n13259) );
  MUX21X1 U13156 ( .IN1(\mem3[99][30] ), .IN2(n1362), .S(n7843), .Q(n13258) );
  MUX21X1 U13157 ( .IN1(\mem3[99][29] ), .IN2(n1340), .S(n7843), .Q(n13257) );
  MUX21X1 U13158 ( .IN1(\mem3[99][28] ), .IN2(n1318), .S(n7843), .Q(n13256) );
  MUX21X1 U13159 ( .IN1(\mem3[99][27] ), .IN2(n1296), .S(n7843), .Q(n13255) );
  MUX21X1 U13160 ( .IN1(\mem3[99][26] ), .IN2(n1274), .S(n7843), .Q(n13254) );
  MUX21X1 U13161 ( .IN1(\mem3[99][25] ), .IN2(n1252), .S(n7843), .Q(n13253) );
  MUX21X1 U13162 ( .IN1(\mem3[99][24] ), .IN2(n1230), .S(n7843), .Q(n13252) );
  AND2X1 U13163 ( .IN1(n7831), .IN2(n7124), .Q(n7843) );
  MUX21X1 U13164 ( .IN1(\mem3[98][31] ), .IN2(n1384), .S(n7844), .Q(n13251) );
  MUX21X1 U13165 ( .IN1(\mem3[98][30] ), .IN2(n1362), .S(n7844), .Q(n13250) );
  MUX21X1 U13166 ( .IN1(\mem3[98][29] ), .IN2(n1340), .S(n7844), .Q(n13249) );
  MUX21X1 U13167 ( .IN1(\mem3[98][28] ), .IN2(n1318), .S(n7844), .Q(n13248) );
  MUX21X1 U13168 ( .IN1(\mem3[98][27] ), .IN2(n1296), .S(n7844), .Q(n13247) );
  MUX21X1 U13169 ( .IN1(\mem3[98][26] ), .IN2(n1274), .S(n7844), .Q(n13246) );
  MUX21X1 U13170 ( .IN1(\mem3[98][25] ), .IN2(n1252), .S(n7844), .Q(n13245) );
  MUX21X1 U13171 ( .IN1(\mem3[98][24] ), .IN2(n1230), .S(n7844), .Q(n13244) );
  AND2X1 U13172 ( .IN1(n7831), .IN2(n7126), .Q(n7844) );
  MUX21X1 U13173 ( .IN1(\mem3[97][31] ), .IN2(n1384), .S(n7845), .Q(n13243) );
  MUX21X1 U13174 ( .IN1(\mem3[97][30] ), .IN2(n1362), .S(n7845), .Q(n13242) );
  MUX21X1 U13175 ( .IN1(\mem3[97][29] ), .IN2(n1340), .S(n7845), .Q(n13241) );
  MUX21X1 U13176 ( .IN1(\mem3[97][28] ), .IN2(n1318), .S(n7845), .Q(n13240) );
  MUX21X1 U13177 ( .IN1(\mem3[97][27] ), .IN2(n1296), .S(n7845), .Q(n13239) );
  MUX21X1 U13178 ( .IN1(\mem3[97][26] ), .IN2(n1274), .S(n7845), .Q(n13238) );
  MUX21X1 U13179 ( .IN1(\mem3[97][25] ), .IN2(n1252), .S(n7845), .Q(n13237) );
  MUX21X1 U13180 ( .IN1(\mem3[97][24] ), .IN2(n1230), .S(n7845), .Q(n13236) );
  AND2X1 U13181 ( .IN1(n7831), .IN2(n7128), .Q(n7845) );
  MUX21X1 U13182 ( .IN1(\mem3[96][31] ), .IN2(n1384), .S(n7846), .Q(n13235) );
  MUX21X1 U13183 ( .IN1(\mem3[96][30] ), .IN2(n1362), .S(n7846), .Q(n13234) );
  MUX21X1 U13184 ( .IN1(\mem3[96][29] ), .IN2(n1340), .S(n7846), .Q(n13233) );
  MUX21X1 U13185 ( .IN1(\mem3[96][28] ), .IN2(n1318), .S(n7846), .Q(n13232) );
  MUX21X1 U13186 ( .IN1(\mem3[96][27] ), .IN2(n1296), .S(n7846), .Q(n13231) );
  MUX21X1 U13187 ( .IN1(\mem3[96][26] ), .IN2(n1274), .S(n7846), .Q(n13230) );
  MUX21X1 U13188 ( .IN1(\mem3[96][25] ), .IN2(n1252), .S(n7846), .Q(n13229) );
  MUX21X1 U13189 ( .IN1(\mem3[96][24] ), .IN2(n1230), .S(n7846), .Q(n13228) );
  AND2X1 U13190 ( .IN1(n7831), .IN2(n7130), .Q(n7846) );
  AND2X1 U13191 ( .IN1(n7693), .IN2(n7294), .Q(n7831) );
  MUX21X1 U13192 ( .IN1(\mem3[95][31] ), .IN2(n1384), .S(n7847), .Q(n13227) );
  MUX21X1 U13193 ( .IN1(\mem3[95][30] ), .IN2(n1362), .S(n7847), .Q(n13226) );
  MUX21X1 U13194 ( .IN1(\mem3[95][29] ), .IN2(n1340), .S(n7847), .Q(n13225) );
  MUX21X1 U13195 ( .IN1(\mem3[95][28] ), .IN2(n1318), .S(n7847), .Q(n13224) );
  MUX21X1 U13196 ( .IN1(\mem3[95][27] ), .IN2(n1296), .S(n7847), .Q(n13223) );
  MUX21X1 U13197 ( .IN1(\mem3[95][26] ), .IN2(n1274), .S(n7847), .Q(n13222) );
  MUX21X1 U13198 ( .IN1(\mem3[95][25] ), .IN2(n1252), .S(n7847), .Q(n13221) );
  MUX21X1 U13199 ( .IN1(\mem3[95][24] ), .IN2(n1230), .S(n7847), .Q(n13220) );
  AND2X1 U13200 ( .IN1(n7848), .IN2(n7099), .Q(n7847) );
  MUX21X1 U13201 ( .IN1(\mem3[94][31] ), .IN2(n1384), .S(n7849), .Q(n13219) );
  MUX21X1 U13202 ( .IN1(\mem3[94][30] ), .IN2(n1362), .S(n7849), .Q(n13218) );
  MUX21X1 U13203 ( .IN1(\mem3[94][29] ), .IN2(n1340), .S(n7849), .Q(n13217) );
  MUX21X1 U13204 ( .IN1(\mem3[94][28] ), .IN2(n1318), .S(n7849), .Q(n13216) );
  MUX21X1 U13205 ( .IN1(\mem3[94][27] ), .IN2(n1296), .S(n7849), .Q(n13215) );
  MUX21X1 U13206 ( .IN1(\mem3[94][26] ), .IN2(n1274), .S(n7849), .Q(n13214) );
  MUX21X1 U13207 ( .IN1(\mem3[94][25] ), .IN2(n1252), .S(n7849), .Q(n13213) );
  MUX21X1 U13208 ( .IN1(\mem3[94][24] ), .IN2(n1230), .S(n7849), .Q(n13212) );
  AND2X1 U13209 ( .IN1(n7848), .IN2(n7102), .Q(n7849) );
  MUX21X1 U13210 ( .IN1(\mem3[93][31] ), .IN2(n1384), .S(n7850), .Q(n13211) );
  MUX21X1 U13211 ( .IN1(\mem3[93][30] ), .IN2(n1362), .S(n7850), .Q(n13210) );
  MUX21X1 U13212 ( .IN1(\mem3[93][29] ), .IN2(n1340), .S(n7850), .Q(n13209) );
  MUX21X1 U13213 ( .IN1(\mem3[93][28] ), .IN2(n1318), .S(n7850), .Q(n13208) );
  MUX21X1 U13214 ( .IN1(\mem3[93][27] ), .IN2(n1296), .S(n7850), .Q(n13207) );
  MUX21X1 U13215 ( .IN1(\mem3[93][26] ), .IN2(n1274), .S(n7850), .Q(n13206) );
  MUX21X1 U13216 ( .IN1(\mem3[93][25] ), .IN2(n1252), .S(n7850), .Q(n13205) );
  MUX21X1 U13217 ( .IN1(\mem3[93][24] ), .IN2(n1230), .S(n7850), .Q(n13204) );
  AND2X1 U13218 ( .IN1(n7848), .IN2(n7104), .Q(n7850) );
  MUX21X1 U13219 ( .IN1(\mem3[92][31] ), .IN2(n1384), .S(n7851), .Q(n13203) );
  MUX21X1 U13220 ( .IN1(\mem3[92][30] ), .IN2(n1362), .S(n7851), .Q(n13202) );
  MUX21X1 U13221 ( .IN1(\mem3[92][29] ), .IN2(n1340), .S(n7851), .Q(n13201) );
  MUX21X1 U13222 ( .IN1(\mem3[92][28] ), .IN2(n1318), .S(n7851), .Q(n13200) );
  MUX21X1 U13223 ( .IN1(\mem3[92][27] ), .IN2(n1296), .S(n7851), .Q(n13199) );
  MUX21X1 U13224 ( .IN1(\mem3[92][26] ), .IN2(n1274), .S(n7851), .Q(n13198) );
  MUX21X1 U13225 ( .IN1(\mem3[92][25] ), .IN2(n1252), .S(n7851), .Q(n13197) );
  MUX21X1 U13226 ( .IN1(\mem3[92][24] ), .IN2(n1230), .S(n7851), .Q(n13196) );
  AND2X1 U13227 ( .IN1(n7848), .IN2(n7106), .Q(n7851) );
  MUX21X1 U13228 ( .IN1(\mem3[91][31] ), .IN2(n1384), .S(n7852), .Q(n13195) );
  MUX21X1 U13229 ( .IN1(\mem3[91][30] ), .IN2(n1362), .S(n7852), .Q(n13194) );
  MUX21X1 U13230 ( .IN1(\mem3[91][29] ), .IN2(n1340), .S(n7852), .Q(n13193) );
  MUX21X1 U13231 ( .IN1(\mem3[91][28] ), .IN2(n1318), .S(n7852), .Q(n13192) );
  MUX21X1 U13232 ( .IN1(\mem3[91][27] ), .IN2(n1296), .S(n7852), .Q(n13191) );
  MUX21X1 U13233 ( .IN1(\mem3[91][26] ), .IN2(n1274), .S(n7852), .Q(n13190) );
  MUX21X1 U13234 ( .IN1(\mem3[91][25] ), .IN2(n1252), .S(n7852), .Q(n13189) );
  MUX21X1 U13235 ( .IN1(\mem3[91][24] ), .IN2(n1230), .S(n7852), .Q(n13188) );
  AND2X1 U13236 ( .IN1(n7848), .IN2(n7108), .Q(n7852) );
  MUX21X1 U13237 ( .IN1(\mem3[90][31] ), .IN2(n1384), .S(n7853), .Q(n13187) );
  MUX21X1 U13238 ( .IN1(\mem3[90][30] ), .IN2(n1362), .S(n7853), .Q(n13186) );
  MUX21X1 U13239 ( .IN1(\mem3[90][29] ), .IN2(n1340), .S(n7853), .Q(n13185) );
  MUX21X1 U13240 ( .IN1(\mem3[90][28] ), .IN2(n1318), .S(n7853), .Q(n13184) );
  MUX21X1 U13241 ( .IN1(\mem3[90][27] ), .IN2(n1296), .S(n7853), .Q(n13183) );
  MUX21X1 U13242 ( .IN1(\mem3[90][26] ), .IN2(n1274), .S(n7853), .Q(n13182) );
  MUX21X1 U13243 ( .IN1(\mem3[90][25] ), .IN2(n1252), .S(n7853), .Q(n13181) );
  MUX21X1 U13244 ( .IN1(\mem3[90][24] ), .IN2(n1230), .S(n7853), .Q(n13180) );
  AND2X1 U13245 ( .IN1(n7848), .IN2(n7110), .Q(n7853) );
  MUX21X1 U13246 ( .IN1(\mem3[89][31] ), .IN2(n1384), .S(n7854), .Q(n13179) );
  MUX21X1 U13247 ( .IN1(\mem3[89][30] ), .IN2(n1362), .S(n7854), .Q(n13178) );
  MUX21X1 U13248 ( .IN1(\mem3[89][29] ), .IN2(n1340), .S(n7854), .Q(n13177) );
  MUX21X1 U13249 ( .IN1(\mem3[89][28] ), .IN2(n1318), .S(n7854), .Q(n13176) );
  MUX21X1 U13250 ( .IN1(\mem3[89][27] ), .IN2(n1296), .S(n7854), .Q(n13175) );
  MUX21X1 U13251 ( .IN1(\mem3[89][26] ), .IN2(n1274), .S(n7854), .Q(n13174) );
  MUX21X1 U13252 ( .IN1(\mem3[89][25] ), .IN2(n1252), .S(n7854), .Q(n13173) );
  MUX21X1 U13253 ( .IN1(\mem3[89][24] ), .IN2(n1230), .S(n7854), .Q(n13172) );
  AND2X1 U13254 ( .IN1(n7848), .IN2(n7112), .Q(n7854) );
  MUX21X1 U13255 ( .IN1(\mem3[88][31] ), .IN2(n1384), .S(n7855), .Q(n13171) );
  MUX21X1 U13256 ( .IN1(\mem3[88][30] ), .IN2(n1362), .S(n7855), .Q(n13170) );
  MUX21X1 U13257 ( .IN1(\mem3[88][29] ), .IN2(n1340), .S(n7855), .Q(n13169) );
  MUX21X1 U13258 ( .IN1(\mem3[88][28] ), .IN2(n1318), .S(n7855), .Q(n13168) );
  MUX21X1 U13259 ( .IN1(\mem3[88][27] ), .IN2(n1296), .S(n7855), .Q(n13167) );
  MUX21X1 U13260 ( .IN1(\mem3[88][26] ), .IN2(n1274), .S(n7855), .Q(n13166) );
  MUX21X1 U13261 ( .IN1(\mem3[88][25] ), .IN2(n1252), .S(n7855), .Q(n13165) );
  MUX21X1 U13262 ( .IN1(\mem3[88][24] ), .IN2(n1230), .S(n7855), .Q(n13164) );
  AND2X1 U13263 ( .IN1(n7848), .IN2(n7114), .Q(n7855) );
  MUX21X1 U13264 ( .IN1(\mem3[87][31] ), .IN2(n1385), .S(n7856), .Q(n13163) );
  MUX21X1 U13265 ( .IN1(\mem3[87][30] ), .IN2(n1363), .S(n7856), .Q(n13162) );
  MUX21X1 U13266 ( .IN1(\mem3[87][29] ), .IN2(n1341), .S(n7856), .Q(n13161) );
  MUX21X1 U13267 ( .IN1(\mem3[87][28] ), .IN2(n1319), .S(n7856), .Q(n13160) );
  MUX21X1 U13268 ( .IN1(\mem3[87][27] ), .IN2(n1297), .S(n7856), .Q(n13159) );
  MUX21X1 U13269 ( .IN1(\mem3[87][26] ), .IN2(n1275), .S(n7856), .Q(n13158) );
  MUX21X1 U13270 ( .IN1(\mem3[87][25] ), .IN2(n1253), .S(n7856), .Q(n13157) );
  MUX21X1 U13271 ( .IN1(\mem3[87][24] ), .IN2(n1231), .S(n7856), .Q(n13156) );
  AND2X1 U13272 ( .IN1(n7848), .IN2(n7116), .Q(n7856) );
  MUX21X1 U13273 ( .IN1(\mem3[86][31] ), .IN2(n1385), .S(n7857), .Q(n13155) );
  MUX21X1 U13274 ( .IN1(\mem3[86][30] ), .IN2(n1363), .S(n7857), .Q(n13154) );
  MUX21X1 U13275 ( .IN1(\mem3[86][29] ), .IN2(n1341), .S(n7857), .Q(n13153) );
  MUX21X1 U13276 ( .IN1(\mem3[86][28] ), .IN2(n1319), .S(n7857), .Q(n13152) );
  MUX21X1 U13277 ( .IN1(\mem3[86][27] ), .IN2(n1297), .S(n7857), .Q(n13151) );
  MUX21X1 U13278 ( .IN1(\mem3[86][26] ), .IN2(n1275), .S(n7857), .Q(n13150) );
  MUX21X1 U13279 ( .IN1(\mem3[86][25] ), .IN2(n1253), .S(n7857), .Q(n13149) );
  MUX21X1 U13280 ( .IN1(\mem3[86][24] ), .IN2(n1231), .S(n7857), .Q(n13148) );
  AND2X1 U13281 ( .IN1(n7848), .IN2(n7118), .Q(n7857) );
  MUX21X1 U13282 ( .IN1(\mem3[85][31] ), .IN2(n1385), .S(n7858), .Q(n13147) );
  MUX21X1 U13283 ( .IN1(\mem3[85][30] ), .IN2(n1363), .S(n7858), .Q(n13146) );
  MUX21X1 U13284 ( .IN1(\mem3[85][29] ), .IN2(n1341), .S(n7858), .Q(n13145) );
  MUX21X1 U13285 ( .IN1(\mem3[85][28] ), .IN2(n1319), .S(n7858), .Q(n13144) );
  MUX21X1 U13286 ( .IN1(\mem3[85][27] ), .IN2(n1297), .S(n7858), .Q(n13143) );
  MUX21X1 U13287 ( .IN1(\mem3[85][26] ), .IN2(n1275), .S(n7858), .Q(n13142) );
  MUX21X1 U13288 ( .IN1(\mem3[85][25] ), .IN2(n1253), .S(n7858), .Q(n13141) );
  MUX21X1 U13289 ( .IN1(\mem3[85][24] ), .IN2(n1231), .S(n7858), .Q(n13140) );
  AND2X1 U13290 ( .IN1(n7848), .IN2(n7120), .Q(n7858) );
  MUX21X1 U13291 ( .IN1(\mem3[84][31] ), .IN2(n1385), .S(n7859), .Q(n13139) );
  MUX21X1 U13292 ( .IN1(\mem3[84][30] ), .IN2(n1363), .S(n7859), .Q(n13138) );
  MUX21X1 U13293 ( .IN1(\mem3[84][29] ), .IN2(n1341), .S(n7859), .Q(n13137) );
  MUX21X1 U13294 ( .IN1(\mem3[84][28] ), .IN2(n1319), .S(n7859), .Q(n13136) );
  MUX21X1 U13295 ( .IN1(\mem3[84][27] ), .IN2(n1297), .S(n7859), .Q(n13135) );
  MUX21X1 U13296 ( .IN1(\mem3[84][26] ), .IN2(n1275), .S(n7859), .Q(n13134) );
  MUX21X1 U13297 ( .IN1(\mem3[84][25] ), .IN2(n1253), .S(n7859), .Q(n13133) );
  MUX21X1 U13298 ( .IN1(\mem3[84][24] ), .IN2(n1231), .S(n7859), .Q(n13132) );
  AND2X1 U13299 ( .IN1(n7848), .IN2(n7122), .Q(n7859) );
  MUX21X1 U13300 ( .IN1(\mem3[83][31] ), .IN2(n1385), .S(n7860), .Q(n13131) );
  MUX21X1 U13301 ( .IN1(\mem3[83][30] ), .IN2(n1363), .S(n7860), .Q(n13130) );
  MUX21X1 U13302 ( .IN1(\mem3[83][29] ), .IN2(n1341), .S(n7860), .Q(n13129) );
  MUX21X1 U13303 ( .IN1(\mem3[83][28] ), .IN2(n1319), .S(n7860), .Q(n13128) );
  MUX21X1 U13304 ( .IN1(\mem3[83][27] ), .IN2(n1297), .S(n7860), .Q(n13127) );
  MUX21X1 U13305 ( .IN1(\mem3[83][26] ), .IN2(n1275), .S(n7860), .Q(n13126) );
  MUX21X1 U13306 ( .IN1(\mem3[83][25] ), .IN2(n1253), .S(n7860), .Q(n13125) );
  MUX21X1 U13307 ( .IN1(\mem3[83][24] ), .IN2(n1231), .S(n7860), .Q(n13124) );
  AND2X1 U13308 ( .IN1(n7848), .IN2(n7124), .Q(n7860) );
  MUX21X1 U13309 ( .IN1(\mem3[82][31] ), .IN2(n1385), .S(n7861), .Q(n13123) );
  MUX21X1 U13310 ( .IN1(\mem3[82][30] ), .IN2(n1363), .S(n7861), .Q(n13122) );
  MUX21X1 U13311 ( .IN1(\mem3[82][29] ), .IN2(n1341), .S(n7861), .Q(n13121) );
  MUX21X1 U13312 ( .IN1(\mem3[82][28] ), .IN2(n1319), .S(n7861), .Q(n13120) );
  MUX21X1 U13313 ( .IN1(\mem3[82][27] ), .IN2(n1297), .S(n7861), .Q(n13119) );
  MUX21X1 U13314 ( .IN1(\mem3[82][26] ), .IN2(n1275), .S(n7861), .Q(n13118) );
  MUX21X1 U13315 ( .IN1(\mem3[82][25] ), .IN2(n1253), .S(n7861), .Q(n13117) );
  MUX21X1 U13316 ( .IN1(\mem3[82][24] ), .IN2(n1231), .S(n7861), .Q(n13116) );
  AND2X1 U13317 ( .IN1(n7848), .IN2(n7126), .Q(n7861) );
  MUX21X1 U13318 ( .IN1(\mem3[81][31] ), .IN2(n1385), .S(n7862), .Q(n13115) );
  MUX21X1 U13319 ( .IN1(\mem3[81][30] ), .IN2(n1363), .S(n7862), .Q(n13114) );
  MUX21X1 U13320 ( .IN1(\mem3[81][29] ), .IN2(n1341), .S(n7862), .Q(n13113) );
  MUX21X1 U13321 ( .IN1(\mem3[81][28] ), .IN2(n1319), .S(n7862), .Q(n13112) );
  MUX21X1 U13322 ( .IN1(\mem3[81][27] ), .IN2(n1297), .S(n7862), .Q(n13111) );
  MUX21X1 U13323 ( .IN1(\mem3[81][26] ), .IN2(n1275), .S(n7862), .Q(n13110) );
  MUX21X1 U13324 ( .IN1(\mem3[81][25] ), .IN2(n1253), .S(n7862), .Q(n13109) );
  MUX21X1 U13325 ( .IN1(\mem3[81][24] ), .IN2(n1231), .S(n7862), .Q(n13108) );
  AND2X1 U13326 ( .IN1(n7848), .IN2(n7128), .Q(n7862) );
  MUX21X1 U13327 ( .IN1(\mem3[80][31] ), .IN2(n1385), .S(n7863), .Q(n13107) );
  MUX21X1 U13328 ( .IN1(\mem3[80][30] ), .IN2(n1363), .S(n7863), .Q(n13106) );
  MUX21X1 U13329 ( .IN1(\mem3[80][29] ), .IN2(n1341), .S(n7863), .Q(n13105) );
  MUX21X1 U13330 ( .IN1(\mem3[80][28] ), .IN2(n1319), .S(n7863), .Q(n13104) );
  MUX21X1 U13331 ( .IN1(\mem3[80][27] ), .IN2(n1297), .S(n7863), .Q(n13103) );
  MUX21X1 U13332 ( .IN1(\mem3[80][26] ), .IN2(n1275), .S(n7863), .Q(n13102) );
  MUX21X1 U13333 ( .IN1(\mem3[80][25] ), .IN2(n1253), .S(n7863), .Q(n13101) );
  MUX21X1 U13334 ( .IN1(\mem3[80][24] ), .IN2(n1231), .S(n7863), .Q(n13100) );
  AND2X1 U13335 ( .IN1(n7848), .IN2(n7130), .Q(n7863) );
  AND2X1 U13336 ( .IN1(n7693), .IN2(n7312), .Q(n7848) );
  MUX21X1 U13337 ( .IN1(\mem3[79][31] ), .IN2(n1385), .S(n7864), .Q(n13099) );
  MUX21X1 U13338 ( .IN1(\mem3[79][30] ), .IN2(n1363), .S(n7864), .Q(n13098) );
  MUX21X1 U13339 ( .IN1(\mem3[79][29] ), .IN2(n1341), .S(n7864), .Q(n13097) );
  MUX21X1 U13340 ( .IN1(\mem3[79][28] ), .IN2(n1319), .S(n7864), .Q(n13096) );
  MUX21X1 U13341 ( .IN1(\mem3[79][27] ), .IN2(n1297), .S(n7864), .Q(n13095) );
  MUX21X1 U13342 ( .IN1(\mem3[79][26] ), .IN2(n1275), .S(n7864), .Q(n13094) );
  MUX21X1 U13343 ( .IN1(\mem3[79][25] ), .IN2(n1253), .S(n7864), .Q(n13093) );
  MUX21X1 U13344 ( .IN1(\mem3[79][24] ), .IN2(n1231), .S(n7864), .Q(n13092) );
  AND2X1 U13345 ( .IN1(n7865), .IN2(n7099), .Q(n7864) );
  MUX21X1 U13346 ( .IN1(\mem3[78][31] ), .IN2(n1385), .S(n7866), .Q(n13091) );
  MUX21X1 U13347 ( .IN1(\mem3[78][30] ), .IN2(n1363), .S(n7866), .Q(n13090) );
  MUX21X1 U13348 ( .IN1(\mem3[78][29] ), .IN2(n1341), .S(n7866), .Q(n13089) );
  MUX21X1 U13349 ( .IN1(\mem3[78][28] ), .IN2(n1319), .S(n7866), .Q(n13088) );
  MUX21X1 U13350 ( .IN1(\mem3[78][27] ), .IN2(n1297), .S(n7866), .Q(n13087) );
  MUX21X1 U13351 ( .IN1(\mem3[78][26] ), .IN2(n1275), .S(n7866), .Q(n13086) );
  MUX21X1 U13352 ( .IN1(\mem3[78][25] ), .IN2(n1253), .S(n7866), .Q(n13085) );
  MUX21X1 U13353 ( .IN1(\mem3[78][24] ), .IN2(n1231), .S(n7866), .Q(n13084) );
  AND2X1 U13354 ( .IN1(n7865), .IN2(n7102), .Q(n7866) );
  MUX21X1 U13355 ( .IN1(\mem3[77][31] ), .IN2(n1385), .S(n7867), .Q(n13083) );
  MUX21X1 U13356 ( .IN1(\mem3[77][30] ), .IN2(n1363), .S(n7867), .Q(n13082) );
  MUX21X1 U13357 ( .IN1(\mem3[77][29] ), .IN2(n1341), .S(n7867), .Q(n13081) );
  MUX21X1 U13358 ( .IN1(\mem3[77][28] ), .IN2(n1319), .S(n7867), .Q(n13080) );
  MUX21X1 U13359 ( .IN1(\mem3[77][27] ), .IN2(n1297), .S(n7867), .Q(n13079) );
  MUX21X1 U13360 ( .IN1(\mem3[77][26] ), .IN2(n1275), .S(n7867), .Q(n13078) );
  MUX21X1 U13361 ( .IN1(\mem3[77][25] ), .IN2(n1253), .S(n7867), .Q(n13077) );
  MUX21X1 U13362 ( .IN1(\mem3[77][24] ), .IN2(n1231), .S(n7867), .Q(n13076) );
  AND2X1 U13363 ( .IN1(n7865), .IN2(n7104), .Q(n7867) );
  MUX21X1 U13364 ( .IN1(\mem3[76][31] ), .IN2(n1385), .S(n7868), .Q(n13075) );
  MUX21X1 U13365 ( .IN1(\mem3[76][30] ), .IN2(n1363), .S(n7868), .Q(n13074) );
  MUX21X1 U13366 ( .IN1(\mem3[76][29] ), .IN2(n1341), .S(n7868), .Q(n13073) );
  MUX21X1 U13367 ( .IN1(\mem3[76][28] ), .IN2(n1319), .S(n7868), .Q(n13072) );
  MUX21X1 U13368 ( .IN1(\mem3[76][27] ), .IN2(n1297), .S(n7868), .Q(n13071) );
  MUX21X1 U13369 ( .IN1(\mem3[76][26] ), .IN2(n1275), .S(n7868), .Q(n13070) );
  MUX21X1 U13370 ( .IN1(\mem3[76][25] ), .IN2(n1253), .S(n7868), .Q(n13069) );
  MUX21X1 U13371 ( .IN1(\mem3[76][24] ), .IN2(n1231), .S(n7868), .Q(n13068) );
  AND2X1 U13372 ( .IN1(n7865), .IN2(n7106), .Q(n7868) );
  MUX21X1 U13373 ( .IN1(\mem3[75][31] ), .IN2(n1386), .S(n7869), .Q(n13067) );
  MUX21X1 U13374 ( .IN1(\mem3[75][30] ), .IN2(n1364), .S(n7869), .Q(n13066) );
  MUX21X1 U13375 ( .IN1(\mem3[75][29] ), .IN2(n1342), .S(n7869), .Q(n13065) );
  MUX21X1 U13376 ( .IN1(\mem3[75][28] ), .IN2(n1320), .S(n7869), .Q(n13064) );
  MUX21X1 U13377 ( .IN1(\mem3[75][27] ), .IN2(n1298), .S(n7869), .Q(n13063) );
  MUX21X1 U13378 ( .IN1(\mem3[75][26] ), .IN2(n1276), .S(n7869), .Q(n13062) );
  MUX21X1 U13379 ( .IN1(\mem3[75][25] ), .IN2(n1254), .S(n7869), .Q(n13061) );
  MUX21X1 U13380 ( .IN1(\mem3[75][24] ), .IN2(n1232), .S(n7869), .Q(n13060) );
  AND2X1 U13381 ( .IN1(n7865), .IN2(n7108), .Q(n7869) );
  MUX21X1 U13382 ( .IN1(\mem3[74][31] ), .IN2(n1386), .S(n7870), .Q(n13059) );
  MUX21X1 U13383 ( .IN1(\mem3[74][30] ), .IN2(n1364), .S(n7870), .Q(n13058) );
  MUX21X1 U13384 ( .IN1(\mem3[74][29] ), .IN2(n1342), .S(n7870), .Q(n13057) );
  MUX21X1 U13385 ( .IN1(\mem3[74][28] ), .IN2(n1320), .S(n7870), .Q(n13056) );
  MUX21X1 U13386 ( .IN1(\mem3[74][27] ), .IN2(n1298), .S(n7870), .Q(n13055) );
  MUX21X1 U13387 ( .IN1(\mem3[74][26] ), .IN2(n1276), .S(n7870), .Q(n13054) );
  MUX21X1 U13388 ( .IN1(\mem3[74][25] ), .IN2(n1254), .S(n7870), .Q(n13053) );
  MUX21X1 U13389 ( .IN1(\mem3[74][24] ), .IN2(n1232), .S(n7870), .Q(n13052) );
  AND2X1 U13390 ( .IN1(n7865), .IN2(n7110), .Q(n7870) );
  MUX21X1 U13391 ( .IN1(\mem3[73][31] ), .IN2(n1386), .S(n7871), .Q(n13051) );
  MUX21X1 U13392 ( .IN1(\mem3[73][30] ), .IN2(n1364), .S(n7871), .Q(n13050) );
  MUX21X1 U13393 ( .IN1(\mem3[73][29] ), .IN2(n1342), .S(n7871), .Q(n13049) );
  MUX21X1 U13394 ( .IN1(\mem3[73][28] ), .IN2(n1320), .S(n7871), .Q(n13048) );
  MUX21X1 U13395 ( .IN1(\mem3[73][27] ), .IN2(n1298), .S(n7871), .Q(n13047) );
  MUX21X1 U13396 ( .IN1(\mem3[73][26] ), .IN2(n1276), .S(n7871), .Q(n13046) );
  MUX21X1 U13397 ( .IN1(\mem3[73][25] ), .IN2(n1254), .S(n7871), .Q(n13045) );
  MUX21X1 U13398 ( .IN1(\mem3[73][24] ), .IN2(n1232), .S(n7871), .Q(n13044) );
  AND2X1 U13399 ( .IN1(n7865), .IN2(n7112), .Q(n7871) );
  MUX21X1 U13400 ( .IN1(\mem3[72][31] ), .IN2(n1386), .S(n7872), .Q(n13043) );
  MUX21X1 U13401 ( .IN1(\mem3[72][30] ), .IN2(n1364), .S(n7872), .Q(n13042) );
  MUX21X1 U13402 ( .IN1(\mem3[72][29] ), .IN2(n1342), .S(n7872), .Q(n13041) );
  MUX21X1 U13403 ( .IN1(\mem3[72][28] ), .IN2(n1320), .S(n7872), .Q(n13040) );
  MUX21X1 U13404 ( .IN1(\mem3[72][27] ), .IN2(n1298), .S(n7872), .Q(n13039) );
  MUX21X1 U13405 ( .IN1(\mem3[72][26] ), .IN2(n1276), .S(n7872), .Q(n13038) );
  MUX21X1 U13406 ( .IN1(\mem3[72][25] ), .IN2(n1254), .S(n7872), .Q(n13037) );
  MUX21X1 U13407 ( .IN1(\mem3[72][24] ), .IN2(n1232), .S(n7872), .Q(n13036) );
  AND2X1 U13408 ( .IN1(n7865), .IN2(n7114), .Q(n7872) );
  MUX21X1 U13409 ( .IN1(\mem3[71][31] ), .IN2(n1386), .S(n7873), .Q(n13035) );
  MUX21X1 U13410 ( .IN1(\mem3[71][30] ), .IN2(n1364), .S(n7873), .Q(n13034) );
  MUX21X1 U13411 ( .IN1(\mem3[71][29] ), .IN2(n1342), .S(n7873), .Q(n13033) );
  MUX21X1 U13412 ( .IN1(\mem3[71][28] ), .IN2(n1320), .S(n7873), .Q(n13032) );
  MUX21X1 U13413 ( .IN1(\mem3[71][27] ), .IN2(n1298), .S(n7873), .Q(n13031) );
  MUX21X1 U13414 ( .IN1(\mem3[71][26] ), .IN2(n1276), .S(n7873), .Q(n13030) );
  MUX21X1 U13415 ( .IN1(\mem3[71][25] ), .IN2(n1254), .S(n7873), .Q(n13029) );
  MUX21X1 U13416 ( .IN1(\mem3[71][24] ), .IN2(n1232), .S(n7873), .Q(n13028) );
  AND2X1 U13417 ( .IN1(n7865), .IN2(n7116), .Q(n7873) );
  MUX21X1 U13418 ( .IN1(\mem3[70][31] ), .IN2(n1386), .S(n7874), .Q(n13027) );
  MUX21X1 U13419 ( .IN1(\mem3[70][30] ), .IN2(n1364), .S(n7874), .Q(n13026) );
  MUX21X1 U13420 ( .IN1(\mem3[70][29] ), .IN2(n1342), .S(n7874), .Q(n13025) );
  MUX21X1 U13421 ( .IN1(\mem3[70][28] ), .IN2(n1320), .S(n7874), .Q(n13024) );
  MUX21X1 U13422 ( .IN1(\mem3[70][27] ), .IN2(n1298), .S(n7874), .Q(n13023) );
  MUX21X1 U13423 ( .IN1(\mem3[70][26] ), .IN2(n1276), .S(n7874), .Q(n13022) );
  MUX21X1 U13424 ( .IN1(\mem3[70][25] ), .IN2(n1254), .S(n7874), .Q(n13021) );
  MUX21X1 U13425 ( .IN1(\mem3[70][24] ), .IN2(n1232), .S(n7874), .Q(n13020) );
  AND2X1 U13426 ( .IN1(n7865), .IN2(n7118), .Q(n7874) );
  MUX21X1 U13427 ( .IN1(\mem3[69][31] ), .IN2(n1386), .S(n7875), .Q(n13019) );
  MUX21X1 U13428 ( .IN1(\mem3[69][30] ), .IN2(n1364), .S(n7875), .Q(n13018) );
  MUX21X1 U13429 ( .IN1(\mem3[69][29] ), .IN2(n1342), .S(n7875), .Q(n13017) );
  MUX21X1 U13430 ( .IN1(\mem3[69][28] ), .IN2(n1320), .S(n7875), .Q(n13016) );
  MUX21X1 U13431 ( .IN1(\mem3[69][27] ), .IN2(n1298), .S(n7875), .Q(n13015) );
  MUX21X1 U13432 ( .IN1(\mem3[69][26] ), .IN2(n1276), .S(n7875), .Q(n13014) );
  MUX21X1 U13433 ( .IN1(\mem3[69][25] ), .IN2(n1254), .S(n7875), .Q(n13013) );
  MUX21X1 U13434 ( .IN1(\mem3[69][24] ), .IN2(n1232), .S(n7875), .Q(n13012) );
  AND2X1 U13435 ( .IN1(n7865), .IN2(n7120), .Q(n7875) );
  MUX21X1 U13436 ( .IN1(\mem3[68][31] ), .IN2(n1386), .S(n7876), .Q(n13011) );
  MUX21X1 U13437 ( .IN1(\mem3[68][30] ), .IN2(n1364), .S(n7876), .Q(n13010) );
  MUX21X1 U13438 ( .IN1(\mem3[68][29] ), .IN2(n1342), .S(n7876), .Q(n13009) );
  MUX21X1 U13439 ( .IN1(\mem3[68][28] ), .IN2(n1320), .S(n7876), .Q(n13008) );
  MUX21X1 U13440 ( .IN1(\mem3[68][27] ), .IN2(n1298), .S(n7876), .Q(n13007) );
  MUX21X1 U13441 ( .IN1(\mem3[68][26] ), .IN2(n1276), .S(n7876), .Q(n13006) );
  MUX21X1 U13442 ( .IN1(\mem3[68][25] ), .IN2(n1254), .S(n7876), .Q(n13005) );
  MUX21X1 U13443 ( .IN1(\mem3[68][24] ), .IN2(n1232), .S(n7876), .Q(n13004) );
  AND2X1 U13444 ( .IN1(n7865), .IN2(n7122), .Q(n7876) );
  MUX21X1 U13445 ( .IN1(\mem3[67][31] ), .IN2(n1386), .S(n7877), .Q(n13003) );
  MUX21X1 U13446 ( .IN1(\mem3[67][30] ), .IN2(n1364), .S(n7877), .Q(n13002) );
  MUX21X1 U13447 ( .IN1(\mem3[67][29] ), .IN2(n1342), .S(n7877), .Q(n13001) );
  MUX21X1 U13448 ( .IN1(\mem3[67][28] ), .IN2(n1320), .S(n7877), .Q(n13000) );
  MUX21X1 U13449 ( .IN1(\mem3[67][27] ), .IN2(n1298), .S(n7877), .Q(n12999) );
  MUX21X1 U13450 ( .IN1(\mem3[67][26] ), .IN2(n1276), .S(n7877), .Q(n12998) );
  MUX21X1 U13451 ( .IN1(\mem3[67][25] ), .IN2(n1254), .S(n7877), .Q(n12997) );
  MUX21X1 U13452 ( .IN1(\mem3[67][24] ), .IN2(n1232), .S(n7877), .Q(n12996) );
  AND2X1 U13453 ( .IN1(n7865), .IN2(n7124), .Q(n7877) );
  MUX21X1 U13454 ( .IN1(\mem3[66][31] ), .IN2(n1386), .S(n7878), .Q(n12995) );
  MUX21X1 U13455 ( .IN1(\mem3[66][30] ), .IN2(n1364), .S(n7878), .Q(n12994) );
  MUX21X1 U13456 ( .IN1(\mem3[66][29] ), .IN2(n1342), .S(n7878), .Q(n12993) );
  MUX21X1 U13457 ( .IN1(\mem3[66][28] ), .IN2(n1320), .S(n7878), .Q(n12992) );
  MUX21X1 U13458 ( .IN1(\mem3[66][27] ), .IN2(n1298), .S(n7878), .Q(n12991) );
  MUX21X1 U13459 ( .IN1(\mem3[66][26] ), .IN2(n1276), .S(n7878), .Q(n12990) );
  MUX21X1 U13460 ( .IN1(\mem3[66][25] ), .IN2(n1254), .S(n7878), .Q(n12989) );
  MUX21X1 U13461 ( .IN1(\mem3[66][24] ), .IN2(n1232), .S(n7878), .Q(n12988) );
  AND2X1 U13462 ( .IN1(n7865), .IN2(n7126), .Q(n7878) );
  MUX21X1 U13463 ( .IN1(\mem3[65][31] ), .IN2(n1386), .S(n7879), .Q(n12987) );
  MUX21X1 U13464 ( .IN1(\mem3[65][30] ), .IN2(n1364), .S(n7879), .Q(n12986) );
  MUX21X1 U13465 ( .IN1(\mem3[65][29] ), .IN2(n1342), .S(n7879), .Q(n12985) );
  MUX21X1 U13466 ( .IN1(\mem3[65][28] ), .IN2(n1320), .S(n7879), .Q(n12984) );
  MUX21X1 U13467 ( .IN1(\mem3[65][27] ), .IN2(n1298), .S(n7879), .Q(n12983) );
  MUX21X1 U13468 ( .IN1(\mem3[65][26] ), .IN2(n1276), .S(n7879), .Q(n12982) );
  MUX21X1 U13469 ( .IN1(\mem3[65][25] ), .IN2(n1254), .S(n7879), .Q(n12981) );
  MUX21X1 U13470 ( .IN1(\mem3[65][24] ), .IN2(n1232), .S(n7879), .Q(n12980) );
  AND2X1 U13471 ( .IN1(n7865), .IN2(n7128), .Q(n7879) );
  MUX21X1 U13472 ( .IN1(\mem3[64][31] ), .IN2(n1386), .S(n7880), .Q(n12979) );
  MUX21X1 U13473 ( .IN1(\mem3[64][30] ), .IN2(n1364), .S(n7880), .Q(n12978) );
  MUX21X1 U13474 ( .IN1(\mem3[64][29] ), .IN2(n1342), .S(n7880), .Q(n12977) );
  MUX21X1 U13475 ( .IN1(\mem3[64][28] ), .IN2(n1320), .S(n7880), .Q(n12976) );
  MUX21X1 U13476 ( .IN1(\mem3[64][27] ), .IN2(n1298), .S(n7880), .Q(n12975) );
  MUX21X1 U13477 ( .IN1(\mem3[64][26] ), .IN2(n1276), .S(n7880), .Q(n12974) );
  MUX21X1 U13478 ( .IN1(\mem3[64][25] ), .IN2(n1254), .S(n7880), .Q(n12973) );
  MUX21X1 U13479 ( .IN1(\mem3[64][24] ), .IN2(n1232), .S(n7880), .Q(n12972) );
  AND2X1 U13480 ( .IN1(n7865), .IN2(n7130), .Q(n7880) );
  AND2X1 U13481 ( .IN1(n7693), .IN2(n7330), .Q(n7865) );
  MUX21X1 U13482 ( .IN1(\mem3[63][31] ), .IN2(n1387), .S(n7881), .Q(n12971) );
  MUX21X1 U13483 ( .IN1(\mem3[63][30] ), .IN2(n1365), .S(n7881), .Q(n12970) );
  MUX21X1 U13484 ( .IN1(\mem3[63][29] ), .IN2(n1343), .S(n7881), .Q(n12969) );
  MUX21X1 U13485 ( .IN1(\mem3[63][28] ), .IN2(n1321), .S(n7881), .Q(n12968) );
  MUX21X1 U13486 ( .IN1(\mem3[63][27] ), .IN2(n1299), .S(n7881), .Q(n12967) );
  MUX21X1 U13487 ( .IN1(\mem3[63][26] ), .IN2(n1277), .S(n7881), .Q(n12966) );
  MUX21X1 U13488 ( .IN1(\mem3[63][25] ), .IN2(n1255), .S(n7881), .Q(n12965) );
  MUX21X1 U13489 ( .IN1(\mem3[63][24] ), .IN2(n1233), .S(n7881), .Q(n12964) );
  AND2X1 U13490 ( .IN1(n7882), .IN2(n7099), .Q(n7881) );
  MUX21X1 U13491 ( .IN1(\mem3[62][31] ), .IN2(n1387), .S(n7883), .Q(n12963) );
  MUX21X1 U13492 ( .IN1(\mem3[62][30] ), .IN2(n1365), .S(n7883), .Q(n12962) );
  MUX21X1 U13493 ( .IN1(\mem3[62][29] ), .IN2(n1343), .S(n7883), .Q(n12961) );
  MUX21X1 U13494 ( .IN1(\mem3[62][28] ), .IN2(n1321), .S(n7883), .Q(n12960) );
  MUX21X1 U13495 ( .IN1(\mem3[62][27] ), .IN2(n1299), .S(n7883), .Q(n12959) );
  MUX21X1 U13496 ( .IN1(\mem3[62][26] ), .IN2(n1277), .S(n7883), .Q(n12958) );
  MUX21X1 U13497 ( .IN1(\mem3[62][25] ), .IN2(n1255), .S(n7883), .Q(n12957) );
  MUX21X1 U13498 ( .IN1(\mem3[62][24] ), .IN2(n1233), .S(n7883), .Q(n12956) );
  AND2X1 U13499 ( .IN1(n7882), .IN2(n7102), .Q(n7883) );
  MUX21X1 U13500 ( .IN1(\mem3[61][31] ), .IN2(n1387), .S(n7884), .Q(n12955) );
  MUX21X1 U13501 ( .IN1(\mem3[61][30] ), .IN2(n1365), .S(n7884), .Q(n12954) );
  MUX21X1 U13502 ( .IN1(\mem3[61][29] ), .IN2(n1343), .S(n7884), .Q(n12953) );
  MUX21X1 U13503 ( .IN1(\mem3[61][28] ), .IN2(n1321), .S(n7884), .Q(n12952) );
  MUX21X1 U13504 ( .IN1(\mem3[61][27] ), .IN2(n1299), .S(n7884), .Q(n12951) );
  MUX21X1 U13505 ( .IN1(\mem3[61][26] ), .IN2(n1277), .S(n7884), .Q(n12950) );
  MUX21X1 U13506 ( .IN1(\mem3[61][25] ), .IN2(n1255), .S(n7884), .Q(n12949) );
  MUX21X1 U13507 ( .IN1(\mem3[61][24] ), .IN2(n1233), .S(n7884), .Q(n12948) );
  AND2X1 U13508 ( .IN1(n7882), .IN2(n7104), .Q(n7884) );
  MUX21X1 U13509 ( .IN1(\mem3[60][31] ), .IN2(n1387), .S(n7885), .Q(n12947) );
  MUX21X1 U13510 ( .IN1(\mem3[60][30] ), .IN2(n1365), .S(n7885), .Q(n12946) );
  MUX21X1 U13511 ( .IN1(\mem3[60][29] ), .IN2(n1343), .S(n7885), .Q(n12945) );
  MUX21X1 U13512 ( .IN1(\mem3[60][28] ), .IN2(n1321), .S(n7885), .Q(n12944) );
  MUX21X1 U13513 ( .IN1(\mem3[60][27] ), .IN2(n1299), .S(n7885), .Q(n12943) );
  MUX21X1 U13514 ( .IN1(\mem3[60][26] ), .IN2(n1277), .S(n7885), .Q(n12942) );
  MUX21X1 U13515 ( .IN1(\mem3[60][25] ), .IN2(n1255), .S(n7885), .Q(n12941) );
  MUX21X1 U13516 ( .IN1(\mem3[60][24] ), .IN2(n1233), .S(n7885), .Q(n12940) );
  AND2X1 U13517 ( .IN1(n7882), .IN2(n7106), .Q(n7885) );
  MUX21X1 U13518 ( .IN1(\mem3[59][31] ), .IN2(n1387), .S(n7886), .Q(n12939) );
  MUX21X1 U13519 ( .IN1(\mem3[59][30] ), .IN2(n1365), .S(n7886), .Q(n12938) );
  MUX21X1 U13520 ( .IN1(\mem3[59][29] ), .IN2(n1343), .S(n7886), .Q(n12937) );
  MUX21X1 U13521 ( .IN1(\mem3[59][28] ), .IN2(n1321), .S(n7886), .Q(n12936) );
  MUX21X1 U13522 ( .IN1(\mem3[59][27] ), .IN2(n1299), .S(n7886), .Q(n12935) );
  MUX21X1 U13523 ( .IN1(\mem3[59][26] ), .IN2(n1277), .S(n7886), .Q(n12934) );
  MUX21X1 U13524 ( .IN1(\mem3[59][25] ), .IN2(n1255), .S(n7886), .Q(n12933) );
  MUX21X1 U13525 ( .IN1(\mem3[59][24] ), .IN2(n1233), .S(n7886), .Q(n12932) );
  AND2X1 U13526 ( .IN1(n7882), .IN2(n7108), .Q(n7886) );
  MUX21X1 U13527 ( .IN1(\mem3[58][31] ), .IN2(n1387), .S(n7887), .Q(n12931) );
  MUX21X1 U13528 ( .IN1(\mem3[58][30] ), .IN2(n1365), .S(n7887), .Q(n12930) );
  MUX21X1 U13529 ( .IN1(\mem3[58][29] ), .IN2(n1343), .S(n7887), .Q(n12929) );
  MUX21X1 U13530 ( .IN1(\mem3[58][28] ), .IN2(n1321), .S(n7887), .Q(n12928) );
  MUX21X1 U13531 ( .IN1(\mem3[58][27] ), .IN2(n1299), .S(n7887), .Q(n12927) );
  MUX21X1 U13532 ( .IN1(\mem3[58][26] ), .IN2(n1277), .S(n7887), .Q(n12926) );
  MUX21X1 U13533 ( .IN1(\mem3[58][25] ), .IN2(n1255), .S(n7887), .Q(n12925) );
  MUX21X1 U13534 ( .IN1(\mem3[58][24] ), .IN2(n1233), .S(n7887), .Q(n12924) );
  AND2X1 U13535 ( .IN1(n7882), .IN2(n7110), .Q(n7887) );
  MUX21X1 U13536 ( .IN1(\mem3[57][31] ), .IN2(n1387), .S(n7888), .Q(n12923) );
  MUX21X1 U13537 ( .IN1(\mem3[57][30] ), .IN2(n1365), .S(n7888), .Q(n12922) );
  MUX21X1 U13538 ( .IN1(\mem3[57][29] ), .IN2(n1343), .S(n7888), .Q(n12921) );
  MUX21X1 U13539 ( .IN1(\mem3[57][28] ), .IN2(n1321), .S(n7888), .Q(n12920) );
  MUX21X1 U13540 ( .IN1(\mem3[57][27] ), .IN2(n1299), .S(n7888), .Q(n12919) );
  MUX21X1 U13541 ( .IN1(\mem3[57][26] ), .IN2(n1277), .S(n7888), .Q(n12918) );
  MUX21X1 U13542 ( .IN1(\mem3[57][25] ), .IN2(n1255), .S(n7888), .Q(n12917) );
  MUX21X1 U13543 ( .IN1(\mem3[57][24] ), .IN2(n1233), .S(n7888), .Q(n12916) );
  AND2X1 U13544 ( .IN1(n7882), .IN2(n7112), .Q(n7888) );
  MUX21X1 U13545 ( .IN1(\mem3[56][31] ), .IN2(n1387), .S(n7889), .Q(n12915) );
  MUX21X1 U13546 ( .IN1(\mem3[56][30] ), .IN2(n1365), .S(n7889), .Q(n12914) );
  MUX21X1 U13547 ( .IN1(\mem3[56][29] ), .IN2(n1343), .S(n7889), .Q(n12913) );
  MUX21X1 U13548 ( .IN1(\mem3[56][28] ), .IN2(n1321), .S(n7889), .Q(n12912) );
  MUX21X1 U13549 ( .IN1(\mem3[56][27] ), .IN2(n1299), .S(n7889), .Q(n12911) );
  MUX21X1 U13550 ( .IN1(\mem3[56][26] ), .IN2(n1277), .S(n7889), .Q(n12910) );
  MUX21X1 U13551 ( .IN1(\mem3[56][25] ), .IN2(n1255), .S(n7889), .Q(n12909) );
  MUX21X1 U13552 ( .IN1(\mem3[56][24] ), .IN2(n1233), .S(n7889), .Q(n12908) );
  AND2X1 U13553 ( .IN1(n7882), .IN2(n7114), .Q(n7889) );
  MUX21X1 U13554 ( .IN1(\mem3[55][31] ), .IN2(n1387), .S(n7890), .Q(n12907) );
  MUX21X1 U13555 ( .IN1(\mem3[55][30] ), .IN2(n1365), .S(n7890), .Q(n12906) );
  MUX21X1 U13556 ( .IN1(\mem3[55][29] ), .IN2(n1343), .S(n7890), .Q(n12905) );
  MUX21X1 U13557 ( .IN1(\mem3[55][28] ), .IN2(n1321), .S(n7890), .Q(n12904) );
  MUX21X1 U13558 ( .IN1(\mem3[55][27] ), .IN2(n1299), .S(n7890), .Q(n12903) );
  MUX21X1 U13559 ( .IN1(\mem3[55][26] ), .IN2(n1277), .S(n7890), .Q(n12902) );
  MUX21X1 U13560 ( .IN1(\mem3[55][25] ), .IN2(n1255), .S(n7890), .Q(n12901) );
  MUX21X1 U13561 ( .IN1(\mem3[55][24] ), .IN2(n1233), .S(n7890), .Q(n12900) );
  AND2X1 U13562 ( .IN1(n7882), .IN2(n7116), .Q(n7890) );
  MUX21X1 U13563 ( .IN1(\mem3[54][31] ), .IN2(n1387), .S(n7891), .Q(n12899) );
  MUX21X1 U13564 ( .IN1(\mem3[54][30] ), .IN2(n1365), .S(n7891), .Q(n12898) );
  MUX21X1 U13565 ( .IN1(\mem3[54][29] ), .IN2(n1343), .S(n7891), .Q(n12897) );
  MUX21X1 U13566 ( .IN1(\mem3[54][28] ), .IN2(n1321), .S(n7891), .Q(n12896) );
  MUX21X1 U13567 ( .IN1(\mem3[54][27] ), .IN2(n1299), .S(n7891), .Q(n12895) );
  MUX21X1 U13568 ( .IN1(\mem3[54][26] ), .IN2(n1277), .S(n7891), .Q(n12894) );
  MUX21X1 U13569 ( .IN1(\mem3[54][25] ), .IN2(n1255), .S(n7891), .Q(n12893) );
  MUX21X1 U13570 ( .IN1(\mem3[54][24] ), .IN2(n1233), .S(n7891), .Q(n12892) );
  AND2X1 U13571 ( .IN1(n7882), .IN2(n7118), .Q(n7891) );
  MUX21X1 U13572 ( .IN1(\mem3[53][31] ), .IN2(n1387), .S(n7892), .Q(n12891) );
  MUX21X1 U13573 ( .IN1(\mem3[53][30] ), .IN2(n1365), .S(n7892), .Q(n12890) );
  MUX21X1 U13574 ( .IN1(\mem3[53][29] ), .IN2(n1343), .S(n7892), .Q(n12889) );
  MUX21X1 U13575 ( .IN1(\mem3[53][28] ), .IN2(n1321), .S(n7892), .Q(n12888) );
  MUX21X1 U13576 ( .IN1(\mem3[53][27] ), .IN2(n1299), .S(n7892), .Q(n12887) );
  MUX21X1 U13577 ( .IN1(\mem3[53][26] ), .IN2(n1277), .S(n7892), .Q(n12886) );
  MUX21X1 U13578 ( .IN1(\mem3[53][25] ), .IN2(n1255), .S(n7892), .Q(n12885) );
  MUX21X1 U13579 ( .IN1(\mem3[53][24] ), .IN2(n1233), .S(n7892), .Q(n12884) );
  AND2X1 U13580 ( .IN1(n7882), .IN2(n7120), .Q(n7892) );
  MUX21X1 U13581 ( .IN1(\mem3[52][31] ), .IN2(n1387), .S(n7893), .Q(n12883) );
  MUX21X1 U13582 ( .IN1(\mem3[52][30] ), .IN2(n1365), .S(n7893), .Q(n12882) );
  MUX21X1 U13583 ( .IN1(\mem3[52][29] ), .IN2(n1343), .S(n7893), .Q(n12881) );
  MUX21X1 U13584 ( .IN1(\mem3[52][28] ), .IN2(n1321), .S(n7893), .Q(n12880) );
  MUX21X1 U13585 ( .IN1(\mem3[52][27] ), .IN2(n1299), .S(n7893), .Q(n12879) );
  MUX21X1 U13586 ( .IN1(\mem3[52][26] ), .IN2(n1277), .S(n7893), .Q(n12878) );
  MUX21X1 U13587 ( .IN1(\mem3[52][25] ), .IN2(n1255), .S(n7893), .Q(n12877) );
  MUX21X1 U13588 ( .IN1(\mem3[52][24] ), .IN2(n1233), .S(n7893), .Q(n12876) );
  AND2X1 U13589 ( .IN1(n7882), .IN2(n7122), .Q(n7893) );
  MUX21X1 U13590 ( .IN1(\mem3[51][31] ), .IN2(n1388), .S(n7894), .Q(n12875) );
  MUX21X1 U13591 ( .IN1(\mem3[51][30] ), .IN2(n1366), .S(n7894), .Q(n12874) );
  MUX21X1 U13592 ( .IN1(\mem3[51][29] ), .IN2(n1344), .S(n7894), .Q(n12873) );
  MUX21X1 U13593 ( .IN1(\mem3[51][28] ), .IN2(n1322), .S(n7894), .Q(n12872) );
  MUX21X1 U13594 ( .IN1(\mem3[51][27] ), .IN2(n1300), .S(n7894), .Q(n12871) );
  MUX21X1 U13595 ( .IN1(\mem3[51][26] ), .IN2(n1278), .S(n7894), .Q(n12870) );
  MUX21X1 U13596 ( .IN1(\mem3[51][25] ), .IN2(n1256), .S(n7894), .Q(n12869) );
  MUX21X1 U13597 ( .IN1(\mem3[51][24] ), .IN2(n1234), .S(n7894), .Q(n12868) );
  AND2X1 U13598 ( .IN1(n7882), .IN2(n7124), .Q(n7894) );
  MUX21X1 U13599 ( .IN1(\mem3[50][31] ), .IN2(n1388), .S(n7895), .Q(n12867) );
  MUX21X1 U13600 ( .IN1(\mem3[50][30] ), .IN2(n1366), .S(n7895), .Q(n12866) );
  MUX21X1 U13601 ( .IN1(\mem3[50][29] ), .IN2(n1344), .S(n7895), .Q(n12865) );
  MUX21X1 U13602 ( .IN1(\mem3[50][28] ), .IN2(n1322), .S(n7895), .Q(n12864) );
  MUX21X1 U13603 ( .IN1(\mem3[50][27] ), .IN2(n1300), .S(n7895), .Q(n12863) );
  MUX21X1 U13604 ( .IN1(\mem3[50][26] ), .IN2(n1278), .S(n7895), .Q(n12862) );
  MUX21X1 U13605 ( .IN1(\mem3[50][25] ), .IN2(n1256), .S(n7895), .Q(n12861) );
  MUX21X1 U13606 ( .IN1(\mem3[50][24] ), .IN2(n1234), .S(n7895), .Q(n12860) );
  AND2X1 U13607 ( .IN1(n7882), .IN2(n7126), .Q(n7895) );
  MUX21X1 U13608 ( .IN1(\mem3[49][31] ), .IN2(n1388), .S(n7896), .Q(n12859) );
  MUX21X1 U13609 ( .IN1(\mem3[49][30] ), .IN2(n1366), .S(n7896), .Q(n12858) );
  MUX21X1 U13610 ( .IN1(\mem3[49][29] ), .IN2(n1344), .S(n7896), .Q(n12857) );
  MUX21X1 U13611 ( .IN1(\mem3[49][28] ), .IN2(n1322), .S(n7896), .Q(n12856) );
  MUX21X1 U13612 ( .IN1(\mem3[49][27] ), .IN2(n1300), .S(n7896), .Q(n12855) );
  MUX21X1 U13613 ( .IN1(\mem3[49][26] ), .IN2(n1278), .S(n7896), .Q(n12854) );
  MUX21X1 U13614 ( .IN1(\mem3[49][25] ), .IN2(n1256), .S(n7896), .Q(n12853) );
  MUX21X1 U13615 ( .IN1(\mem3[49][24] ), .IN2(n1234), .S(n7896), .Q(n12852) );
  AND2X1 U13616 ( .IN1(n7882), .IN2(n7128), .Q(n7896) );
  MUX21X1 U13617 ( .IN1(\mem3[48][31] ), .IN2(n1388), .S(n7897), .Q(n12851) );
  MUX21X1 U13618 ( .IN1(\mem3[48][30] ), .IN2(n1366), .S(n7897), .Q(n12850) );
  MUX21X1 U13619 ( .IN1(\mem3[48][29] ), .IN2(n1344), .S(n7897), .Q(n12849) );
  MUX21X1 U13620 ( .IN1(\mem3[48][28] ), .IN2(n1322), .S(n7897), .Q(n12848) );
  MUX21X1 U13621 ( .IN1(\mem3[48][27] ), .IN2(n1300), .S(n7897), .Q(n12847) );
  MUX21X1 U13622 ( .IN1(\mem3[48][26] ), .IN2(n1278), .S(n7897), .Q(n12846) );
  MUX21X1 U13623 ( .IN1(\mem3[48][25] ), .IN2(n1256), .S(n7897), .Q(n12845) );
  MUX21X1 U13624 ( .IN1(\mem3[48][24] ), .IN2(n1234), .S(n7897), .Q(n12844) );
  AND2X1 U13625 ( .IN1(n7882), .IN2(n7130), .Q(n7897) );
  AND2X1 U13626 ( .IN1(n7693), .IN2(n7348), .Q(n7882) );
  MUX21X1 U13627 ( .IN1(\mem3[47][31] ), .IN2(n1388), .S(n7898), .Q(n12843) );
  MUX21X1 U13628 ( .IN1(\mem3[47][30] ), .IN2(n1366), .S(n7898), .Q(n12842) );
  MUX21X1 U13629 ( .IN1(\mem3[47][29] ), .IN2(n1344), .S(n7898), .Q(n12841) );
  MUX21X1 U13630 ( .IN1(\mem3[47][28] ), .IN2(n1322), .S(n7898), .Q(n12840) );
  MUX21X1 U13631 ( .IN1(\mem3[47][27] ), .IN2(n1300), .S(n7898), .Q(n12839) );
  MUX21X1 U13632 ( .IN1(\mem3[47][26] ), .IN2(n1278), .S(n7898), .Q(n12838) );
  MUX21X1 U13633 ( .IN1(\mem3[47][25] ), .IN2(n1256), .S(n7898), .Q(n12837) );
  MUX21X1 U13634 ( .IN1(\mem3[47][24] ), .IN2(n1234), .S(n7898), .Q(n12836) );
  AND2X1 U13635 ( .IN1(n7899), .IN2(n7099), .Q(n7898) );
  MUX21X1 U13636 ( .IN1(\mem3[46][31] ), .IN2(n1388), .S(n7900), .Q(n12835) );
  MUX21X1 U13637 ( .IN1(\mem3[46][30] ), .IN2(n1366), .S(n7900), .Q(n12834) );
  MUX21X1 U13638 ( .IN1(\mem3[46][29] ), .IN2(n1344), .S(n7900), .Q(n12833) );
  MUX21X1 U13639 ( .IN1(\mem3[46][28] ), .IN2(n1322), .S(n7900), .Q(n12832) );
  MUX21X1 U13640 ( .IN1(\mem3[46][27] ), .IN2(n1300), .S(n7900), .Q(n12831) );
  MUX21X1 U13641 ( .IN1(\mem3[46][26] ), .IN2(n1278), .S(n7900), .Q(n12830) );
  MUX21X1 U13642 ( .IN1(\mem3[46][25] ), .IN2(n1256), .S(n7900), .Q(n12829) );
  MUX21X1 U13643 ( .IN1(\mem3[46][24] ), .IN2(n1234), .S(n7900), .Q(n12828) );
  AND2X1 U13644 ( .IN1(n7899), .IN2(n7102), .Q(n7900) );
  MUX21X1 U13645 ( .IN1(\mem3[45][31] ), .IN2(n1388), .S(n7901), .Q(n12827) );
  MUX21X1 U13646 ( .IN1(\mem3[45][30] ), .IN2(n1366), .S(n7901), .Q(n12826) );
  MUX21X1 U13647 ( .IN1(\mem3[45][29] ), .IN2(n1344), .S(n7901), .Q(n12825) );
  MUX21X1 U13648 ( .IN1(\mem3[45][28] ), .IN2(n1322), .S(n7901), .Q(n12824) );
  MUX21X1 U13649 ( .IN1(\mem3[45][27] ), .IN2(n1300), .S(n7901), .Q(n12823) );
  MUX21X1 U13650 ( .IN1(\mem3[45][26] ), .IN2(n1278), .S(n7901), .Q(n12822) );
  MUX21X1 U13651 ( .IN1(\mem3[45][25] ), .IN2(n1256), .S(n7901), .Q(n12821) );
  MUX21X1 U13652 ( .IN1(\mem3[45][24] ), .IN2(n1234), .S(n7901), .Q(n12820) );
  AND2X1 U13653 ( .IN1(n7899), .IN2(n7104), .Q(n7901) );
  MUX21X1 U13654 ( .IN1(\mem3[44][31] ), .IN2(n1388), .S(n7902), .Q(n12819) );
  MUX21X1 U13655 ( .IN1(\mem3[44][30] ), .IN2(n1366), .S(n7902), .Q(n12818) );
  MUX21X1 U13656 ( .IN1(\mem3[44][29] ), .IN2(n1344), .S(n7902), .Q(n12817) );
  MUX21X1 U13657 ( .IN1(\mem3[44][28] ), .IN2(n1322), .S(n7902), .Q(n12816) );
  MUX21X1 U13658 ( .IN1(\mem3[44][27] ), .IN2(n1300), .S(n7902), .Q(n12815) );
  MUX21X1 U13659 ( .IN1(\mem3[44][26] ), .IN2(n1278), .S(n7902), .Q(n12814) );
  MUX21X1 U13660 ( .IN1(\mem3[44][25] ), .IN2(n1256), .S(n7902), .Q(n12813) );
  MUX21X1 U13661 ( .IN1(\mem3[44][24] ), .IN2(n1234), .S(n7902), .Q(n12812) );
  AND2X1 U13662 ( .IN1(n7899), .IN2(n7106), .Q(n7902) );
  MUX21X1 U13663 ( .IN1(\mem3[43][31] ), .IN2(n1388), .S(n7903), .Q(n12811) );
  MUX21X1 U13664 ( .IN1(\mem3[43][30] ), .IN2(n1366), .S(n7903), .Q(n12810) );
  MUX21X1 U13665 ( .IN1(\mem3[43][29] ), .IN2(n1344), .S(n7903), .Q(n12809) );
  MUX21X1 U13666 ( .IN1(\mem3[43][28] ), .IN2(n1322), .S(n7903), .Q(n12808) );
  MUX21X1 U13667 ( .IN1(\mem3[43][27] ), .IN2(n1300), .S(n7903), .Q(n12807) );
  MUX21X1 U13668 ( .IN1(\mem3[43][26] ), .IN2(n1278), .S(n7903), .Q(n12806) );
  MUX21X1 U13669 ( .IN1(\mem3[43][25] ), .IN2(n1256), .S(n7903), .Q(n12805) );
  MUX21X1 U13670 ( .IN1(\mem3[43][24] ), .IN2(n1234), .S(n7903), .Q(n12804) );
  AND2X1 U13671 ( .IN1(n7899), .IN2(n7108), .Q(n7903) );
  MUX21X1 U13672 ( .IN1(\mem3[42][31] ), .IN2(n1388), .S(n7904), .Q(n12803) );
  MUX21X1 U13673 ( .IN1(\mem3[42][30] ), .IN2(n1366), .S(n7904), .Q(n12802) );
  MUX21X1 U13674 ( .IN1(\mem3[42][29] ), .IN2(n1344), .S(n7904), .Q(n12801) );
  MUX21X1 U13675 ( .IN1(\mem3[42][28] ), .IN2(n1322), .S(n7904), .Q(n12800) );
  MUX21X1 U13676 ( .IN1(\mem3[42][27] ), .IN2(n1300), .S(n7904), .Q(n12799) );
  MUX21X1 U13677 ( .IN1(\mem3[42][26] ), .IN2(n1278), .S(n7904), .Q(n12798) );
  MUX21X1 U13678 ( .IN1(\mem3[42][25] ), .IN2(n1256), .S(n7904), .Q(n12797) );
  MUX21X1 U13679 ( .IN1(\mem3[42][24] ), .IN2(n1234), .S(n7904), .Q(n12796) );
  AND2X1 U13680 ( .IN1(n7899), .IN2(n7110), .Q(n7904) );
  MUX21X1 U13681 ( .IN1(\mem3[41][31] ), .IN2(n1388), .S(n7905), .Q(n12795) );
  MUX21X1 U13682 ( .IN1(\mem3[41][30] ), .IN2(n1366), .S(n7905), .Q(n12794) );
  MUX21X1 U13683 ( .IN1(\mem3[41][29] ), .IN2(n1344), .S(n7905), .Q(n12793) );
  MUX21X1 U13684 ( .IN1(\mem3[41][28] ), .IN2(n1322), .S(n7905), .Q(n12792) );
  MUX21X1 U13685 ( .IN1(\mem3[41][27] ), .IN2(n1300), .S(n7905), .Q(n12791) );
  MUX21X1 U13686 ( .IN1(\mem3[41][26] ), .IN2(n1278), .S(n7905), .Q(n12790) );
  MUX21X1 U13687 ( .IN1(\mem3[41][25] ), .IN2(n1256), .S(n7905), .Q(n12789) );
  MUX21X1 U13688 ( .IN1(\mem3[41][24] ), .IN2(n1234), .S(n7905), .Q(n12788) );
  AND2X1 U13689 ( .IN1(n7899), .IN2(n7112), .Q(n7905) );
  MUX21X1 U13690 ( .IN1(\mem3[40][31] ), .IN2(n1388), .S(n7906), .Q(n12787) );
  MUX21X1 U13691 ( .IN1(\mem3[40][30] ), .IN2(n1366), .S(n7906), .Q(n12786) );
  MUX21X1 U13692 ( .IN1(\mem3[40][29] ), .IN2(n1344), .S(n7906), .Q(n12785) );
  MUX21X1 U13693 ( .IN1(\mem3[40][28] ), .IN2(n1322), .S(n7906), .Q(n12784) );
  MUX21X1 U13694 ( .IN1(\mem3[40][27] ), .IN2(n1300), .S(n7906), .Q(n12783) );
  MUX21X1 U13695 ( .IN1(\mem3[40][26] ), .IN2(n1278), .S(n7906), .Q(n12782) );
  MUX21X1 U13696 ( .IN1(\mem3[40][25] ), .IN2(n1256), .S(n7906), .Q(n12781) );
  MUX21X1 U13697 ( .IN1(\mem3[40][24] ), .IN2(n1234), .S(n7906), .Q(n12780) );
  AND2X1 U13698 ( .IN1(n7899), .IN2(n7114), .Q(n7906) );
  MUX21X1 U13699 ( .IN1(\mem3[39][31] ), .IN2(n1389), .S(n7907), .Q(n12779) );
  MUX21X1 U13700 ( .IN1(\mem3[39][30] ), .IN2(n1367), .S(n7907), .Q(n12778) );
  MUX21X1 U13701 ( .IN1(\mem3[39][29] ), .IN2(n1345), .S(n7907), .Q(n12777) );
  MUX21X1 U13702 ( .IN1(\mem3[39][28] ), .IN2(n1323), .S(n7907), .Q(n12776) );
  MUX21X1 U13703 ( .IN1(\mem3[39][27] ), .IN2(n1301), .S(n7907), .Q(n12775) );
  MUX21X1 U13704 ( .IN1(\mem3[39][26] ), .IN2(n1279), .S(n7907), .Q(n12774) );
  MUX21X1 U13705 ( .IN1(\mem3[39][25] ), .IN2(n1257), .S(n7907), .Q(n12773) );
  MUX21X1 U13706 ( .IN1(\mem3[39][24] ), .IN2(n1235), .S(n7907), .Q(n12772) );
  AND2X1 U13707 ( .IN1(n7899), .IN2(n7116), .Q(n7907) );
  MUX21X1 U13708 ( .IN1(\mem3[38][31] ), .IN2(n1389), .S(n7908), .Q(n12771) );
  MUX21X1 U13709 ( .IN1(\mem3[38][30] ), .IN2(n1367), .S(n7908), .Q(n12770) );
  MUX21X1 U13710 ( .IN1(\mem3[38][29] ), .IN2(n1345), .S(n7908), .Q(n12769) );
  MUX21X1 U13711 ( .IN1(\mem3[38][28] ), .IN2(n1323), .S(n7908), .Q(n12768) );
  MUX21X1 U13712 ( .IN1(\mem3[38][27] ), .IN2(n1301), .S(n7908), .Q(n12767) );
  MUX21X1 U13713 ( .IN1(\mem3[38][26] ), .IN2(n1279), .S(n7908), .Q(n12766) );
  MUX21X1 U13714 ( .IN1(\mem3[38][25] ), .IN2(n1257), .S(n7908), .Q(n12765) );
  MUX21X1 U13715 ( .IN1(\mem3[38][24] ), .IN2(n1235), .S(n7908), .Q(n12764) );
  AND2X1 U13716 ( .IN1(n7899), .IN2(n7118), .Q(n7908) );
  MUX21X1 U13717 ( .IN1(\mem3[37][31] ), .IN2(n1389), .S(n7909), .Q(n12763) );
  MUX21X1 U13718 ( .IN1(\mem3[37][30] ), .IN2(n1367), .S(n7909), .Q(n12762) );
  MUX21X1 U13719 ( .IN1(\mem3[37][29] ), .IN2(n1345), .S(n7909), .Q(n12761) );
  MUX21X1 U13720 ( .IN1(\mem3[37][28] ), .IN2(n1323), .S(n7909), .Q(n12760) );
  MUX21X1 U13721 ( .IN1(\mem3[37][27] ), .IN2(n1301), .S(n7909), .Q(n12759) );
  MUX21X1 U13722 ( .IN1(\mem3[37][26] ), .IN2(n1279), .S(n7909), .Q(n12758) );
  MUX21X1 U13723 ( .IN1(\mem3[37][25] ), .IN2(n1257), .S(n7909), .Q(n12757) );
  MUX21X1 U13724 ( .IN1(\mem3[37][24] ), .IN2(n1235), .S(n7909), .Q(n12756) );
  AND2X1 U13725 ( .IN1(n7899), .IN2(n7120), .Q(n7909) );
  MUX21X1 U13726 ( .IN1(\mem3[36][31] ), .IN2(n1389), .S(n7910), .Q(n12755) );
  MUX21X1 U13727 ( .IN1(\mem3[36][30] ), .IN2(n1367), .S(n7910), .Q(n12754) );
  MUX21X1 U13728 ( .IN1(\mem3[36][29] ), .IN2(n1345), .S(n7910), .Q(n12753) );
  MUX21X1 U13729 ( .IN1(\mem3[36][28] ), .IN2(n1323), .S(n7910), .Q(n12752) );
  MUX21X1 U13730 ( .IN1(\mem3[36][27] ), .IN2(n1301), .S(n7910), .Q(n12751) );
  MUX21X1 U13731 ( .IN1(\mem3[36][26] ), .IN2(n1279), .S(n7910), .Q(n12750) );
  MUX21X1 U13732 ( .IN1(\mem3[36][25] ), .IN2(n1257), .S(n7910), .Q(n12749) );
  MUX21X1 U13733 ( .IN1(\mem3[36][24] ), .IN2(n1235), .S(n7910), .Q(n12748) );
  AND2X1 U13734 ( .IN1(n7899), .IN2(n7122), .Q(n7910) );
  MUX21X1 U13735 ( .IN1(\mem3[35][31] ), .IN2(n1389), .S(n7911), .Q(n12747) );
  MUX21X1 U13736 ( .IN1(\mem3[35][30] ), .IN2(n1367), .S(n7911), .Q(n12746) );
  MUX21X1 U13737 ( .IN1(\mem3[35][29] ), .IN2(n1345), .S(n7911), .Q(n12745) );
  MUX21X1 U13738 ( .IN1(\mem3[35][28] ), .IN2(n1323), .S(n7911), .Q(n12744) );
  MUX21X1 U13739 ( .IN1(\mem3[35][27] ), .IN2(n1301), .S(n7911), .Q(n12743) );
  MUX21X1 U13740 ( .IN1(\mem3[35][26] ), .IN2(n1279), .S(n7911), .Q(n12742) );
  MUX21X1 U13741 ( .IN1(\mem3[35][25] ), .IN2(n1257), .S(n7911), .Q(n12741) );
  MUX21X1 U13742 ( .IN1(\mem3[35][24] ), .IN2(n1235), .S(n7911), .Q(n12740) );
  AND2X1 U13743 ( .IN1(n7899), .IN2(n7124), .Q(n7911) );
  MUX21X1 U13744 ( .IN1(\mem3[34][31] ), .IN2(n1389), .S(n7912), .Q(n12739) );
  MUX21X1 U13745 ( .IN1(\mem3[34][30] ), .IN2(n1367), .S(n7912), .Q(n12738) );
  MUX21X1 U13746 ( .IN1(\mem3[34][29] ), .IN2(n1345), .S(n7912), .Q(n12737) );
  MUX21X1 U13747 ( .IN1(\mem3[34][28] ), .IN2(n1323), .S(n7912), .Q(n12736) );
  MUX21X1 U13748 ( .IN1(\mem3[34][27] ), .IN2(n1301), .S(n7912), .Q(n12735) );
  MUX21X1 U13749 ( .IN1(\mem3[34][26] ), .IN2(n1279), .S(n7912), .Q(n12734) );
  MUX21X1 U13750 ( .IN1(\mem3[34][25] ), .IN2(n1257), .S(n7912), .Q(n12733) );
  MUX21X1 U13751 ( .IN1(\mem3[34][24] ), .IN2(n1235), .S(n7912), .Q(n12732) );
  AND2X1 U13752 ( .IN1(n7899), .IN2(n7126), .Q(n7912) );
  MUX21X1 U13753 ( .IN1(\mem3[33][31] ), .IN2(n1389), .S(n7913), .Q(n12731) );
  MUX21X1 U13754 ( .IN1(\mem3[33][30] ), .IN2(n1367), .S(n7913), .Q(n12730) );
  MUX21X1 U13755 ( .IN1(\mem3[33][29] ), .IN2(n1345), .S(n7913), .Q(n12729) );
  MUX21X1 U13756 ( .IN1(\mem3[33][28] ), .IN2(n1323), .S(n7913), .Q(n12728) );
  MUX21X1 U13757 ( .IN1(\mem3[33][27] ), .IN2(n1301), .S(n7913), .Q(n12727) );
  MUX21X1 U13758 ( .IN1(\mem3[33][26] ), .IN2(n1279), .S(n7913), .Q(n12726) );
  MUX21X1 U13759 ( .IN1(\mem3[33][25] ), .IN2(n1257), .S(n7913), .Q(n12725) );
  MUX21X1 U13760 ( .IN1(\mem3[33][24] ), .IN2(n1235), .S(n7913), .Q(n12724) );
  AND2X1 U13761 ( .IN1(n7899), .IN2(n7128), .Q(n7913) );
  MUX21X1 U13762 ( .IN1(\mem3[32][31] ), .IN2(n1389), .S(n7914), .Q(n12723) );
  MUX21X1 U13763 ( .IN1(\mem3[32][30] ), .IN2(n1367), .S(n7914), .Q(n12722) );
  MUX21X1 U13764 ( .IN1(\mem3[32][29] ), .IN2(n1345), .S(n7914), .Q(n12721) );
  MUX21X1 U13765 ( .IN1(\mem3[32][28] ), .IN2(n1323), .S(n7914), .Q(n12720) );
  MUX21X1 U13766 ( .IN1(\mem3[32][27] ), .IN2(n1301), .S(n7914), .Q(n12719) );
  MUX21X1 U13767 ( .IN1(\mem3[32][26] ), .IN2(n1279), .S(n7914), .Q(n12718) );
  MUX21X1 U13768 ( .IN1(\mem3[32][25] ), .IN2(n1257), .S(n7914), .Q(n12717) );
  MUX21X1 U13769 ( .IN1(\mem3[32][24] ), .IN2(n1235), .S(n7914), .Q(n12716) );
  AND2X1 U13770 ( .IN1(n7899), .IN2(n7130), .Q(n7914) );
  AND2X1 U13771 ( .IN1(n7693), .IN2(n7366), .Q(n7899) );
  MUX21X1 U13772 ( .IN1(\mem3[31][31] ), .IN2(n1389), .S(n7915), .Q(n12715) );
  MUX21X1 U13773 ( .IN1(\mem3[31][30] ), .IN2(n1367), .S(n7915), .Q(n12714) );
  MUX21X1 U13774 ( .IN1(\mem3[31][29] ), .IN2(n1345), .S(n7915), .Q(n12713) );
  MUX21X1 U13775 ( .IN1(\mem3[31][28] ), .IN2(n1323), .S(n7915), .Q(n12712) );
  MUX21X1 U13776 ( .IN1(\mem3[31][27] ), .IN2(n1301), .S(n7915), .Q(n12711) );
  MUX21X1 U13777 ( .IN1(\mem3[31][26] ), .IN2(n1279), .S(n7915), .Q(n12710) );
  MUX21X1 U13778 ( .IN1(\mem3[31][25] ), .IN2(n1257), .S(n7915), .Q(n12709) );
  MUX21X1 U13779 ( .IN1(\mem3[31][24] ), .IN2(n1235), .S(n7915), .Q(n12708) );
  AND2X1 U13780 ( .IN1(n7916), .IN2(n7099), .Q(n7915) );
  MUX21X1 U13781 ( .IN1(\mem3[30][31] ), .IN2(n1389), .S(n7917), .Q(n12707) );
  MUX21X1 U13782 ( .IN1(\mem3[30][30] ), .IN2(n1367), .S(n7917), .Q(n12706) );
  MUX21X1 U13783 ( .IN1(\mem3[30][29] ), .IN2(n1345), .S(n7917), .Q(n12705) );
  MUX21X1 U13784 ( .IN1(\mem3[30][28] ), .IN2(n1323), .S(n7917), .Q(n12704) );
  MUX21X1 U13785 ( .IN1(\mem3[30][27] ), .IN2(n1301), .S(n7917), .Q(n12703) );
  MUX21X1 U13786 ( .IN1(\mem3[30][26] ), .IN2(n1279), .S(n7917), .Q(n12702) );
  MUX21X1 U13787 ( .IN1(\mem3[30][25] ), .IN2(n1257), .S(n7917), .Q(n12701) );
  MUX21X1 U13788 ( .IN1(\mem3[30][24] ), .IN2(n1235), .S(n7917), .Q(n12700) );
  AND2X1 U13789 ( .IN1(n7916), .IN2(n7102), .Q(n7917) );
  MUX21X1 U13790 ( .IN1(\mem3[29][31] ), .IN2(n1389), .S(n7918), .Q(n12699) );
  MUX21X1 U13791 ( .IN1(\mem3[29][30] ), .IN2(n1367), .S(n7918), .Q(n12698) );
  MUX21X1 U13792 ( .IN1(\mem3[29][29] ), .IN2(n1345), .S(n7918), .Q(n12697) );
  MUX21X1 U13793 ( .IN1(\mem3[29][28] ), .IN2(n1323), .S(n7918), .Q(n12696) );
  MUX21X1 U13794 ( .IN1(\mem3[29][27] ), .IN2(n1301), .S(n7918), .Q(n12695) );
  MUX21X1 U13795 ( .IN1(\mem3[29][26] ), .IN2(n1279), .S(n7918), .Q(n12694) );
  MUX21X1 U13796 ( .IN1(\mem3[29][25] ), .IN2(n1257), .S(n7918), .Q(n12693) );
  MUX21X1 U13797 ( .IN1(\mem3[29][24] ), .IN2(n1235), .S(n7918), .Q(n12692) );
  AND2X1 U13798 ( .IN1(n7916), .IN2(n7104), .Q(n7918) );
  MUX21X1 U13799 ( .IN1(\mem3[28][31] ), .IN2(n1389), .S(n7919), .Q(n12691) );
  MUX21X1 U13800 ( .IN1(\mem3[28][30] ), .IN2(n1367), .S(n7919), .Q(n12690) );
  MUX21X1 U13801 ( .IN1(\mem3[28][29] ), .IN2(n1345), .S(n7919), .Q(n12689) );
  MUX21X1 U13802 ( .IN1(\mem3[28][28] ), .IN2(n1323), .S(n7919), .Q(n12688) );
  MUX21X1 U13803 ( .IN1(\mem3[28][27] ), .IN2(n1301), .S(n7919), .Q(n12687) );
  MUX21X1 U13804 ( .IN1(\mem3[28][26] ), .IN2(n1279), .S(n7919), .Q(n12686) );
  MUX21X1 U13805 ( .IN1(\mem3[28][25] ), .IN2(n1257), .S(n7919), .Q(n12685) );
  MUX21X1 U13806 ( .IN1(\mem3[28][24] ), .IN2(n1235), .S(n7919), .Q(n12684) );
  AND2X1 U13807 ( .IN1(n7916), .IN2(n7106), .Q(n7919) );
  MUX21X1 U13808 ( .IN1(\mem3[27][31] ), .IN2(n1390), .S(n7920), .Q(n12683) );
  MUX21X1 U13809 ( .IN1(\mem3[27][30] ), .IN2(n1368), .S(n7920), .Q(n12682) );
  MUX21X1 U13810 ( .IN1(\mem3[27][29] ), .IN2(n1346), .S(n7920), .Q(n12681) );
  MUX21X1 U13811 ( .IN1(\mem3[27][28] ), .IN2(n1324), .S(n7920), .Q(n12680) );
  MUX21X1 U13812 ( .IN1(\mem3[27][27] ), .IN2(n1302), .S(n7920), .Q(n12679) );
  MUX21X1 U13813 ( .IN1(\mem3[27][26] ), .IN2(n1280), .S(n7920), .Q(n12678) );
  MUX21X1 U13814 ( .IN1(\mem3[27][25] ), .IN2(n1258), .S(n7920), .Q(n12677) );
  MUX21X1 U13815 ( .IN1(\mem3[27][24] ), .IN2(n1236), .S(n7920), .Q(n12676) );
  AND2X1 U13816 ( .IN1(n7916), .IN2(n7108), .Q(n7920) );
  MUX21X1 U13817 ( .IN1(\mem3[26][31] ), .IN2(n1390), .S(n7921), .Q(n12675) );
  MUX21X1 U13818 ( .IN1(\mem3[26][30] ), .IN2(n1368), .S(n7921), .Q(n12674) );
  MUX21X1 U13819 ( .IN1(\mem3[26][29] ), .IN2(n1346), .S(n7921), .Q(n12673) );
  MUX21X1 U13820 ( .IN1(\mem3[26][28] ), .IN2(n1324), .S(n7921), .Q(n12672) );
  MUX21X1 U13821 ( .IN1(\mem3[26][27] ), .IN2(n1302), .S(n7921), .Q(n12671) );
  MUX21X1 U13822 ( .IN1(\mem3[26][26] ), .IN2(n1280), .S(n7921), .Q(n12670) );
  MUX21X1 U13823 ( .IN1(\mem3[26][25] ), .IN2(n1258), .S(n7921), .Q(n12669) );
  MUX21X1 U13824 ( .IN1(\mem3[26][24] ), .IN2(n1236), .S(n7921), .Q(n12668) );
  AND2X1 U13825 ( .IN1(n7916), .IN2(n7110), .Q(n7921) );
  MUX21X1 U13826 ( .IN1(\mem3[25][31] ), .IN2(n1390), .S(n7922), .Q(n12667) );
  MUX21X1 U13827 ( .IN1(\mem3[25][30] ), .IN2(n1368), .S(n7922), .Q(n12666) );
  MUX21X1 U13828 ( .IN1(\mem3[25][29] ), .IN2(n1346), .S(n7922), .Q(n12665) );
  MUX21X1 U13829 ( .IN1(\mem3[25][28] ), .IN2(n1324), .S(n7922), .Q(n12664) );
  MUX21X1 U13830 ( .IN1(\mem3[25][27] ), .IN2(n1302), .S(n7922), .Q(n12663) );
  MUX21X1 U13831 ( .IN1(\mem3[25][26] ), .IN2(n1280), .S(n7922), .Q(n12662) );
  MUX21X1 U13832 ( .IN1(\mem3[25][25] ), .IN2(n1258), .S(n7922), .Q(n12661) );
  MUX21X1 U13833 ( .IN1(\mem3[25][24] ), .IN2(n1236), .S(n7922), .Q(n12660) );
  AND2X1 U13834 ( .IN1(n7916), .IN2(n7112), .Q(n7922) );
  MUX21X1 U13835 ( .IN1(\mem3[24][31] ), .IN2(n1390), .S(n7923), .Q(n12659) );
  MUX21X1 U13836 ( .IN1(\mem3[24][30] ), .IN2(n1368), .S(n7923), .Q(n12658) );
  MUX21X1 U13837 ( .IN1(\mem3[24][29] ), .IN2(n1346), .S(n7923), .Q(n12657) );
  MUX21X1 U13838 ( .IN1(\mem3[24][28] ), .IN2(n1324), .S(n7923), .Q(n12656) );
  MUX21X1 U13839 ( .IN1(\mem3[24][27] ), .IN2(n1302), .S(n7923), .Q(n12655) );
  MUX21X1 U13840 ( .IN1(\mem3[24][26] ), .IN2(n1280), .S(n7923), .Q(n12654) );
  MUX21X1 U13841 ( .IN1(\mem3[24][25] ), .IN2(n1258), .S(n7923), .Q(n12653) );
  MUX21X1 U13842 ( .IN1(\mem3[24][24] ), .IN2(n1236), .S(n7923), .Q(n12652) );
  AND2X1 U13843 ( .IN1(n7916), .IN2(n7114), .Q(n7923) );
  MUX21X1 U13844 ( .IN1(\mem3[23][31] ), .IN2(n1390), .S(n7924), .Q(n12651) );
  MUX21X1 U13845 ( .IN1(\mem3[23][30] ), .IN2(n1368), .S(n7924), .Q(n12650) );
  MUX21X1 U13846 ( .IN1(\mem3[23][29] ), .IN2(n1346), .S(n7924), .Q(n12649) );
  MUX21X1 U13847 ( .IN1(\mem3[23][28] ), .IN2(n1324), .S(n7924), .Q(n12648) );
  MUX21X1 U13848 ( .IN1(\mem3[23][27] ), .IN2(n1302), .S(n7924), .Q(n12647) );
  MUX21X1 U13849 ( .IN1(\mem3[23][26] ), .IN2(n1280), .S(n7924), .Q(n12646) );
  MUX21X1 U13850 ( .IN1(\mem3[23][25] ), .IN2(n1258), .S(n7924), .Q(n12645) );
  MUX21X1 U13851 ( .IN1(\mem3[23][24] ), .IN2(n1236), .S(n7924), .Q(n12644) );
  AND2X1 U13852 ( .IN1(n7916), .IN2(n7116), .Q(n7924) );
  MUX21X1 U13853 ( .IN1(\mem3[22][31] ), .IN2(n1390), .S(n7925), .Q(n12643) );
  MUX21X1 U13854 ( .IN1(\mem3[22][30] ), .IN2(n1368), .S(n7925), .Q(n12642) );
  MUX21X1 U13855 ( .IN1(\mem3[22][29] ), .IN2(n1346), .S(n7925), .Q(n12641) );
  MUX21X1 U13856 ( .IN1(\mem3[22][28] ), .IN2(n1324), .S(n7925), .Q(n12640) );
  MUX21X1 U13857 ( .IN1(\mem3[22][27] ), .IN2(n1302), .S(n7925), .Q(n12639) );
  MUX21X1 U13858 ( .IN1(\mem3[22][26] ), .IN2(n1280), .S(n7925), .Q(n12638) );
  MUX21X1 U13859 ( .IN1(\mem3[22][25] ), .IN2(n1258), .S(n7925), .Q(n12637) );
  MUX21X1 U13860 ( .IN1(\mem3[22][24] ), .IN2(n1236), .S(n7925), .Q(n12636) );
  AND2X1 U13861 ( .IN1(n7916), .IN2(n7118), .Q(n7925) );
  MUX21X1 U13862 ( .IN1(\mem3[21][31] ), .IN2(n1390), .S(n7926), .Q(n12635) );
  MUX21X1 U13863 ( .IN1(\mem3[21][30] ), .IN2(n1368), .S(n7926), .Q(n12634) );
  MUX21X1 U13864 ( .IN1(\mem3[21][29] ), .IN2(n1346), .S(n7926), .Q(n12633) );
  MUX21X1 U13865 ( .IN1(\mem3[21][28] ), .IN2(n1324), .S(n7926), .Q(n12632) );
  MUX21X1 U13866 ( .IN1(\mem3[21][27] ), .IN2(n1302), .S(n7926), .Q(n12631) );
  MUX21X1 U13867 ( .IN1(\mem3[21][26] ), .IN2(n1280), .S(n7926), .Q(n12630) );
  MUX21X1 U13868 ( .IN1(\mem3[21][25] ), .IN2(n1258), .S(n7926), .Q(n12629) );
  MUX21X1 U13869 ( .IN1(\mem3[21][24] ), .IN2(n1236), .S(n7926), .Q(n12628) );
  AND2X1 U13870 ( .IN1(n7916), .IN2(n7120), .Q(n7926) );
  MUX21X1 U13871 ( .IN1(\mem3[20][31] ), .IN2(n1390), .S(n7927), .Q(n12627) );
  MUX21X1 U13872 ( .IN1(\mem3[20][30] ), .IN2(n1368), .S(n7927), .Q(n12626) );
  MUX21X1 U13873 ( .IN1(\mem3[20][29] ), .IN2(n1346), .S(n7927), .Q(n12625) );
  MUX21X1 U13874 ( .IN1(\mem3[20][28] ), .IN2(n1324), .S(n7927), .Q(n12624) );
  MUX21X1 U13875 ( .IN1(\mem3[20][27] ), .IN2(n1302), .S(n7927), .Q(n12623) );
  MUX21X1 U13876 ( .IN1(\mem3[20][26] ), .IN2(n1280), .S(n7927), .Q(n12622) );
  MUX21X1 U13877 ( .IN1(\mem3[20][25] ), .IN2(n1258), .S(n7927), .Q(n12621) );
  MUX21X1 U13878 ( .IN1(\mem3[20][24] ), .IN2(n1236), .S(n7927), .Q(n12620) );
  AND2X1 U13879 ( .IN1(n7916), .IN2(n7122), .Q(n7927) );
  MUX21X1 U13880 ( .IN1(\mem3[19][31] ), .IN2(n1390), .S(n7928), .Q(n12619) );
  MUX21X1 U13881 ( .IN1(\mem3[19][30] ), .IN2(n1368), .S(n7928), .Q(n12618) );
  MUX21X1 U13882 ( .IN1(\mem3[19][29] ), .IN2(n1346), .S(n7928), .Q(n12617) );
  MUX21X1 U13883 ( .IN1(\mem3[19][28] ), .IN2(n1324), .S(n7928), .Q(n12616) );
  MUX21X1 U13884 ( .IN1(\mem3[19][27] ), .IN2(n1302), .S(n7928), .Q(n12615) );
  MUX21X1 U13885 ( .IN1(\mem3[19][26] ), .IN2(n1280), .S(n7928), .Q(n12614) );
  MUX21X1 U13886 ( .IN1(\mem3[19][25] ), .IN2(n1258), .S(n7928), .Q(n12613) );
  MUX21X1 U13887 ( .IN1(\mem3[19][24] ), .IN2(n1236), .S(n7928), .Q(n12612) );
  AND2X1 U13888 ( .IN1(n7916), .IN2(n7124), .Q(n7928) );
  MUX21X1 U13889 ( .IN1(\mem3[18][31] ), .IN2(n1390), .S(n7929), .Q(n12611) );
  MUX21X1 U13890 ( .IN1(\mem3[18][30] ), .IN2(n1368), .S(n7929), .Q(n12610) );
  MUX21X1 U13891 ( .IN1(\mem3[18][29] ), .IN2(n1346), .S(n7929), .Q(n12609) );
  MUX21X1 U13892 ( .IN1(\mem3[18][28] ), .IN2(n1324), .S(n7929), .Q(n12608) );
  MUX21X1 U13893 ( .IN1(\mem3[18][27] ), .IN2(n1302), .S(n7929), .Q(n12607) );
  MUX21X1 U13894 ( .IN1(\mem3[18][26] ), .IN2(n1280), .S(n7929), .Q(n12606) );
  MUX21X1 U13895 ( .IN1(\mem3[18][25] ), .IN2(n1258), .S(n7929), .Q(n12605) );
  MUX21X1 U13896 ( .IN1(\mem3[18][24] ), .IN2(n1236), .S(n7929), .Q(n12604) );
  AND2X1 U13897 ( .IN1(n7916), .IN2(n7126), .Q(n7929) );
  MUX21X1 U13898 ( .IN1(\mem3[17][31] ), .IN2(n1390), .S(n7930), .Q(n12603) );
  MUX21X1 U13899 ( .IN1(\mem3[17][30] ), .IN2(n1368), .S(n7930), .Q(n12602) );
  MUX21X1 U13900 ( .IN1(\mem3[17][29] ), .IN2(n1346), .S(n7930), .Q(n12601) );
  MUX21X1 U13901 ( .IN1(\mem3[17][28] ), .IN2(n1324), .S(n7930), .Q(n12600) );
  MUX21X1 U13902 ( .IN1(\mem3[17][27] ), .IN2(n1302), .S(n7930), .Q(n12599) );
  MUX21X1 U13903 ( .IN1(\mem3[17][26] ), .IN2(n1280), .S(n7930), .Q(n12598) );
  MUX21X1 U13904 ( .IN1(\mem3[17][25] ), .IN2(n1258), .S(n7930), .Q(n12597) );
  MUX21X1 U13905 ( .IN1(\mem3[17][24] ), .IN2(n1236), .S(n7930), .Q(n12596) );
  AND2X1 U13906 ( .IN1(n7916), .IN2(n7128), .Q(n7930) );
  MUX21X1 U13907 ( .IN1(\mem3[16][31] ), .IN2(n1390), .S(n7931), .Q(n12595) );
  MUX21X1 U13908 ( .IN1(\mem3[16][30] ), .IN2(n1368), .S(n7931), .Q(n12594) );
  MUX21X1 U13909 ( .IN1(\mem3[16][29] ), .IN2(n1346), .S(n7931), .Q(n12593) );
  MUX21X1 U13910 ( .IN1(\mem3[16][28] ), .IN2(n1324), .S(n7931), .Q(n12592) );
  MUX21X1 U13911 ( .IN1(\mem3[16][27] ), .IN2(n1302), .S(n7931), .Q(n12591) );
  MUX21X1 U13912 ( .IN1(\mem3[16][26] ), .IN2(n1280), .S(n7931), .Q(n12590) );
  MUX21X1 U13913 ( .IN1(\mem3[16][25] ), .IN2(n1258), .S(n7931), .Q(n12589) );
  MUX21X1 U13914 ( .IN1(\mem3[16][24] ), .IN2(n1236), .S(n7931), .Q(n12588) );
  AND2X1 U13915 ( .IN1(n7916), .IN2(n7130), .Q(n7931) );
  AND2X1 U13916 ( .IN1(n7693), .IN2(n7384), .Q(n7916) );
  MUX21X1 U13917 ( .IN1(\mem3[15][31] ), .IN2(n1391), .S(n7932), .Q(n12587) );
  MUX21X1 U13918 ( .IN1(\mem3[15][30] ), .IN2(n1369), .S(n7932), .Q(n12586) );
  MUX21X1 U13919 ( .IN1(\mem3[15][29] ), .IN2(n1347), .S(n7932), .Q(n12585) );
  MUX21X1 U13920 ( .IN1(\mem3[15][28] ), .IN2(n1325), .S(n7932), .Q(n12584) );
  MUX21X1 U13921 ( .IN1(\mem3[15][27] ), .IN2(n1303), .S(n7932), .Q(n12583) );
  MUX21X1 U13922 ( .IN1(\mem3[15][26] ), .IN2(n1281), .S(n7932), .Q(n12582) );
  MUX21X1 U13923 ( .IN1(\mem3[15][25] ), .IN2(n1259), .S(n7932), .Q(n12581) );
  MUX21X1 U13924 ( .IN1(\mem3[15][24] ), .IN2(n1237), .S(n7932), .Q(n12580) );
  AND2X1 U13925 ( .IN1(n7933), .IN2(n7099), .Q(n7932) );
  MUX21X1 U13926 ( .IN1(\mem3[14][31] ), .IN2(n1391), .S(n7934), .Q(n12579) );
  MUX21X1 U13927 ( .IN1(\mem3[14][30] ), .IN2(n1369), .S(n7934), .Q(n12578) );
  MUX21X1 U13928 ( .IN1(\mem3[14][29] ), .IN2(n1347), .S(n7934), .Q(n12577) );
  MUX21X1 U13929 ( .IN1(\mem3[14][28] ), .IN2(n1325), .S(n7934), .Q(n12576) );
  MUX21X1 U13930 ( .IN1(\mem3[14][27] ), .IN2(n1303), .S(n7934), .Q(n12575) );
  MUX21X1 U13931 ( .IN1(\mem3[14][26] ), .IN2(n1281), .S(n7934), .Q(n12574) );
  MUX21X1 U13932 ( .IN1(\mem3[14][25] ), .IN2(n1259), .S(n7934), .Q(n12573) );
  MUX21X1 U13933 ( .IN1(\mem3[14][24] ), .IN2(n1237), .S(n7934), .Q(n12572) );
  AND2X1 U13934 ( .IN1(n7933), .IN2(n7102), .Q(n7934) );
  MUX21X1 U13935 ( .IN1(\mem3[13][31] ), .IN2(n1391), .S(n7935), .Q(n12571) );
  MUX21X1 U13936 ( .IN1(\mem3[13][30] ), .IN2(n1369), .S(n7935), .Q(n12570) );
  MUX21X1 U13937 ( .IN1(\mem3[13][29] ), .IN2(n1347), .S(n7935), .Q(n12569) );
  MUX21X1 U13938 ( .IN1(\mem3[13][28] ), .IN2(n1325), .S(n7935), .Q(n12568) );
  MUX21X1 U13939 ( .IN1(\mem3[13][27] ), .IN2(n1303), .S(n7935), .Q(n12567) );
  MUX21X1 U13940 ( .IN1(\mem3[13][26] ), .IN2(n1281), .S(n7935), .Q(n12566) );
  MUX21X1 U13941 ( .IN1(\mem3[13][25] ), .IN2(n1259), .S(n7935), .Q(n12565) );
  MUX21X1 U13942 ( .IN1(\mem3[13][24] ), .IN2(n1237), .S(n7935), .Q(n12564) );
  AND2X1 U13943 ( .IN1(n7933), .IN2(n7104), .Q(n7935) );
  MUX21X1 U13944 ( .IN1(\mem3[12][31] ), .IN2(n1391), .S(n7936), .Q(n12563) );
  MUX21X1 U13945 ( .IN1(\mem3[12][30] ), .IN2(n1369), .S(n7936), .Q(n12562) );
  MUX21X1 U13946 ( .IN1(\mem3[12][29] ), .IN2(n1347), .S(n7936), .Q(n12561) );
  MUX21X1 U13947 ( .IN1(\mem3[12][28] ), .IN2(n1325), .S(n7936), .Q(n12560) );
  MUX21X1 U13948 ( .IN1(\mem3[12][27] ), .IN2(n1303), .S(n7936), .Q(n12559) );
  MUX21X1 U13949 ( .IN1(\mem3[12][26] ), .IN2(n1281), .S(n7936), .Q(n12558) );
  MUX21X1 U13950 ( .IN1(\mem3[12][25] ), .IN2(n1259), .S(n7936), .Q(n12557) );
  MUX21X1 U13951 ( .IN1(\mem3[12][24] ), .IN2(n1237), .S(n7936), .Q(n12556) );
  AND2X1 U13952 ( .IN1(n7933), .IN2(n7106), .Q(n7936) );
  MUX21X1 U13953 ( .IN1(\mem3[11][31] ), .IN2(n1391), .S(n7937), .Q(n12555) );
  MUX21X1 U13954 ( .IN1(\mem3[11][30] ), .IN2(n1369), .S(n7937), .Q(n12554) );
  MUX21X1 U13955 ( .IN1(\mem3[11][29] ), .IN2(n1347), .S(n7937), .Q(n12553) );
  MUX21X1 U13956 ( .IN1(\mem3[11][28] ), .IN2(n1325), .S(n7937), .Q(n12552) );
  MUX21X1 U13957 ( .IN1(\mem3[11][27] ), .IN2(n1303), .S(n7937), .Q(n12551) );
  MUX21X1 U13958 ( .IN1(\mem3[11][26] ), .IN2(n1281), .S(n7937), .Q(n12550) );
  MUX21X1 U13959 ( .IN1(\mem3[11][25] ), .IN2(n1259), .S(n7937), .Q(n12549) );
  MUX21X1 U13960 ( .IN1(\mem3[11][24] ), .IN2(n1237), .S(n7937), .Q(n12548) );
  AND2X1 U13961 ( .IN1(n7933), .IN2(n7108), .Q(n7937) );
  MUX21X1 U13962 ( .IN1(\mem3[10][31] ), .IN2(n1391), .S(n7938), .Q(n12547) );
  MUX21X1 U13963 ( .IN1(\mem3[10][30] ), .IN2(n1369), .S(n7938), .Q(n12546) );
  MUX21X1 U13964 ( .IN1(\mem3[10][29] ), .IN2(n1347), .S(n7938), .Q(n12545) );
  MUX21X1 U13965 ( .IN1(\mem3[10][28] ), .IN2(n1325), .S(n7938), .Q(n12544) );
  MUX21X1 U13966 ( .IN1(\mem3[10][27] ), .IN2(n1303), .S(n7938), .Q(n12543) );
  MUX21X1 U13967 ( .IN1(\mem3[10][26] ), .IN2(n1281), .S(n7938), .Q(n12542) );
  MUX21X1 U13968 ( .IN1(\mem3[10][25] ), .IN2(n1259), .S(n7938), .Q(n12541) );
  MUX21X1 U13969 ( .IN1(\mem3[10][24] ), .IN2(n1237), .S(n7938), .Q(n12540) );
  AND2X1 U13970 ( .IN1(n7933), .IN2(n7110), .Q(n7938) );
  MUX21X1 U13971 ( .IN1(\mem3[9][31] ), .IN2(n1391), .S(n7939), .Q(n12539) );
  MUX21X1 U13972 ( .IN1(\mem3[9][30] ), .IN2(n1369), .S(n7939), .Q(n12538) );
  MUX21X1 U13973 ( .IN1(\mem3[9][29] ), .IN2(n1347), .S(n7939), .Q(n12537) );
  MUX21X1 U13974 ( .IN1(\mem3[9][28] ), .IN2(n1325), .S(n7939), .Q(n12536) );
  MUX21X1 U13975 ( .IN1(\mem3[9][27] ), .IN2(n1303), .S(n7939), .Q(n12535) );
  MUX21X1 U13976 ( .IN1(\mem3[9][26] ), .IN2(n1281), .S(n7939), .Q(n12534) );
  MUX21X1 U13977 ( .IN1(\mem3[9][25] ), .IN2(n1259), .S(n7939), .Q(n12533) );
  MUX21X1 U13978 ( .IN1(\mem3[9][24] ), .IN2(n1237), .S(n7939), .Q(n12532) );
  AND2X1 U13979 ( .IN1(n7933), .IN2(n7112), .Q(n7939) );
  MUX21X1 U13980 ( .IN1(\mem3[8][31] ), .IN2(n1391), .S(n7940), .Q(n12531) );
  MUX21X1 U13981 ( .IN1(\mem3[8][30] ), .IN2(n1369), .S(n7940), .Q(n12530) );
  MUX21X1 U13982 ( .IN1(\mem3[8][29] ), .IN2(n1347), .S(n7940), .Q(n12529) );
  MUX21X1 U13983 ( .IN1(\mem3[8][28] ), .IN2(n1325), .S(n7940), .Q(n12528) );
  MUX21X1 U13984 ( .IN1(\mem3[8][27] ), .IN2(n1303), .S(n7940), .Q(n12527) );
  MUX21X1 U13985 ( .IN1(\mem3[8][26] ), .IN2(n1281), .S(n7940), .Q(n12526) );
  MUX21X1 U13986 ( .IN1(\mem3[8][25] ), .IN2(n1259), .S(n7940), .Q(n12525) );
  MUX21X1 U13987 ( .IN1(\mem3[8][24] ), .IN2(n1237), .S(n7940), .Q(n12524) );
  AND2X1 U13988 ( .IN1(n7933), .IN2(n7114), .Q(n7940) );
  MUX21X1 U13989 ( .IN1(\mem3[7][31] ), .IN2(n1391), .S(n7941), .Q(n12523) );
  MUX21X1 U13990 ( .IN1(\mem3[7][30] ), .IN2(n1369), .S(n7941), .Q(n12522) );
  MUX21X1 U13991 ( .IN1(\mem3[7][29] ), .IN2(n1347), .S(n7941), .Q(n12521) );
  MUX21X1 U13992 ( .IN1(\mem3[7][28] ), .IN2(n1325), .S(n7941), .Q(n12520) );
  MUX21X1 U13993 ( .IN1(\mem3[7][27] ), .IN2(n1303), .S(n7941), .Q(n12519) );
  MUX21X1 U13994 ( .IN1(\mem3[7][26] ), .IN2(n1281), .S(n7941), .Q(n12518) );
  MUX21X1 U13995 ( .IN1(\mem3[7][25] ), .IN2(n1259), .S(n7941), .Q(n12517) );
  MUX21X1 U13996 ( .IN1(\mem3[7][24] ), .IN2(n1237), .S(n7941), .Q(n12516) );
  AND2X1 U13997 ( .IN1(n7933), .IN2(n7116), .Q(n7941) );
  MUX21X1 U13998 ( .IN1(\mem3[6][31] ), .IN2(n1391), .S(n7942), .Q(n12515) );
  MUX21X1 U13999 ( .IN1(\mem3[6][30] ), .IN2(n1369), .S(n7942), .Q(n12514) );
  MUX21X1 U14000 ( .IN1(\mem3[6][29] ), .IN2(n1347), .S(n7942), .Q(n12513) );
  MUX21X1 U14001 ( .IN1(\mem3[6][28] ), .IN2(n1325), .S(n7942), .Q(n12512) );
  MUX21X1 U14002 ( .IN1(\mem3[6][27] ), .IN2(n1303), .S(n7942), .Q(n12511) );
  MUX21X1 U14003 ( .IN1(\mem3[6][26] ), .IN2(n1281), .S(n7942), .Q(n12510) );
  MUX21X1 U14004 ( .IN1(\mem3[6][25] ), .IN2(n1259), .S(n7942), .Q(n12509) );
  MUX21X1 U14005 ( .IN1(\mem3[6][24] ), .IN2(n1237), .S(n7942), .Q(n12508) );
  AND2X1 U14006 ( .IN1(n7933), .IN2(n7118), .Q(n7942) );
  MUX21X1 U14007 ( .IN1(\mem3[5][31] ), .IN2(n1391), .S(n7943), .Q(n12507) );
  MUX21X1 U14008 ( .IN1(\mem3[5][30] ), .IN2(n1369), .S(n7943), .Q(n12506) );
  MUX21X1 U14009 ( .IN1(\mem3[5][29] ), .IN2(n1347), .S(n7943), .Q(n12505) );
  MUX21X1 U14010 ( .IN1(\mem3[5][28] ), .IN2(n1325), .S(n7943), .Q(n12504) );
  MUX21X1 U14011 ( .IN1(\mem3[5][27] ), .IN2(n1303), .S(n7943), .Q(n12503) );
  MUX21X1 U14012 ( .IN1(\mem3[5][26] ), .IN2(n1281), .S(n7943), .Q(n12502) );
  MUX21X1 U14013 ( .IN1(\mem3[5][25] ), .IN2(n1259), .S(n7943), .Q(n12501) );
  MUX21X1 U14014 ( .IN1(\mem3[5][24] ), .IN2(n1237), .S(n7943), .Q(n12500) );
  AND2X1 U14015 ( .IN1(n7933), .IN2(n7120), .Q(n7943) );
  MUX21X1 U14016 ( .IN1(\mem3[4][31] ), .IN2(n1391), .S(n7944), .Q(n12499) );
  MUX21X1 U14017 ( .IN1(\mem3[4][30] ), .IN2(n1369), .S(n7944), .Q(n12498) );
  MUX21X1 U14018 ( .IN1(\mem3[4][29] ), .IN2(n1347), .S(n7944), .Q(n12497) );
  MUX21X1 U14019 ( .IN1(\mem3[4][28] ), .IN2(n1325), .S(n7944), .Q(n12496) );
  MUX21X1 U14020 ( .IN1(\mem3[4][27] ), .IN2(n1303), .S(n7944), .Q(n12495) );
  MUX21X1 U14021 ( .IN1(\mem3[4][26] ), .IN2(n1281), .S(n7944), .Q(n12494) );
  MUX21X1 U14022 ( .IN1(\mem3[4][25] ), .IN2(n1259), .S(n7944), .Q(n12493) );
  MUX21X1 U14023 ( .IN1(\mem3[4][24] ), .IN2(n1237), .S(n7944), .Q(n12492) );
  AND2X1 U14024 ( .IN1(n7933), .IN2(n7122), .Q(n7944) );
  MUX21X1 U14025 ( .IN1(\mem3[3][31] ), .IN2(n1392), .S(n7945), .Q(n12491) );
  MUX21X1 U14026 ( .IN1(\mem3[3][30] ), .IN2(n1370), .S(n7945), .Q(n12490) );
  MUX21X1 U14027 ( .IN1(\mem3[3][29] ), .IN2(n1348), .S(n7945), .Q(n12489) );
  MUX21X1 U14028 ( .IN1(\mem3[3][28] ), .IN2(n1326), .S(n7945), .Q(n12488) );
  MUX21X1 U14029 ( .IN1(\mem3[3][27] ), .IN2(n1304), .S(n7945), .Q(n12487) );
  MUX21X1 U14030 ( .IN1(\mem3[3][26] ), .IN2(n1282), .S(n7945), .Q(n12486) );
  MUX21X1 U14031 ( .IN1(\mem3[3][25] ), .IN2(n1260), .S(n7945), .Q(n12485) );
  MUX21X1 U14032 ( .IN1(\mem3[3][24] ), .IN2(n1238), .S(n7945), .Q(n12484) );
  AND2X1 U14033 ( .IN1(n7933), .IN2(n7124), .Q(n7945) );
  MUX21X1 U14034 ( .IN1(\mem3[2][31] ), .IN2(n1392), .S(n7946), .Q(n12483) );
  MUX21X1 U14035 ( .IN1(\mem3[2][30] ), .IN2(n1370), .S(n7946), .Q(n12482) );
  MUX21X1 U14036 ( .IN1(\mem3[2][29] ), .IN2(n1348), .S(n7946), .Q(n12481) );
  MUX21X1 U14037 ( .IN1(\mem3[2][28] ), .IN2(n1326), .S(n7946), .Q(n12480) );
  MUX21X1 U14038 ( .IN1(\mem3[2][27] ), .IN2(n1304), .S(n7946), .Q(n12479) );
  MUX21X1 U14039 ( .IN1(\mem3[2][26] ), .IN2(n1282), .S(n7946), .Q(n12478) );
  MUX21X1 U14040 ( .IN1(\mem3[2][25] ), .IN2(n1260), .S(n7946), .Q(n12477) );
  MUX21X1 U14041 ( .IN1(\mem3[2][24] ), .IN2(n1238), .S(n7946), .Q(n12476) );
  AND2X1 U14042 ( .IN1(n7933), .IN2(n7126), .Q(n7946) );
  MUX21X1 U14043 ( .IN1(\mem3[1][31] ), .IN2(n1392), .S(n7947), .Q(n12475) );
  MUX21X1 U14044 ( .IN1(\mem3[1][30] ), .IN2(n1370), .S(n7947), .Q(n12474) );
  MUX21X1 U14045 ( .IN1(\mem3[1][29] ), .IN2(n1348), .S(n7947), .Q(n12473) );
  MUX21X1 U14046 ( .IN1(\mem3[1][28] ), .IN2(n1326), .S(n7947), .Q(n12472) );
  MUX21X1 U14047 ( .IN1(\mem3[1][27] ), .IN2(n1304), .S(n7947), .Q(n12471) );
  MUX21X1 U14048 ( .IN1(\mem3[1][26] ), .IN2(n1282), .S(n7947), .Q(n12470) );
  MUX21X1 U14049 ( .IN1(\mem3[1][25] ), .IN2(n1260), .S(n7947), .Q(n12469) );
  MUX21X1 U14050 ( .IN1(\mem3[1][24] ), .IN2(n1238), .S(n7947), .Q(n12468) );
  AND2X1 U14051 ( .IN1(n7933), .IN2(n7128), .Q(n7947) );
  MUX21X1 U14052 ( .IN1(\mem3[0][31] ), .IN2(n1392), .S(n7948), .Q(n12467) );
  MUX21X1 U14053 ( .IN1(\mem3[0][30] ), .IN2(n1370), .S(n7948), .Q(n12466) );
  MUX21X1 U14054 ( .IN1(\mem3[0][29] ), .IN2(n1348), .S(n7948), .Q(n12465) );
  MUX21X1 U14055 ( .IN1(\mem3[0][28] ), .IN2(n1326), .S(n7948), .Q(n12464) );
  MUX21X1 U14056 ( .IN1(\mem3[0][27] ), .IN2(n1304), .S(n7948), .Q(n12463) );
  MUX21X1 U14057 ( .IN1(\mem3[0][26] ), .IN2(n1282), .S(n7948), .Q(n12462) );
  MUX21X1 U14058 ( .IN1(\mem3[0][25] ), .IN2(n1260), .S(n7948), .Q(n12461) );
  MUX21X1 U14059 ( .IN1(\mem3[0][24] ), .IN2(n1238), .S(n7948), .Q(n12460) );
  AND2X1 U14060 ( .IN1(n7933), .IN2(n7130), .Q(n7948) );
  AND2X1 U14061 ( .IN1(n7693), .IN2(n7402), .Q(n7933) );
  AND2X1 U14062 ( .IN1(we[3]), .IN2(ce), .Q(n7693) );
  MUX21X1 U14063 ( .IN1(\mem2[255][23] ), .IN2(n1195), .S(n7949), .Q(n12459)
         );
  MUX21X1 U14064 ( .IN1(\mem2[255][22] ), .IN2(n1173), .S(n7949), .Q(n12458)
         );
  MUX21X1 U14065 ( .IN1(\mem2[255][21] ), .IN2(n1151), .S(n7949), .Q(n12457)
         );
  MUX21X1 U14066 ( .IN1(\mem2[255][20] ), .IN2(n1129), .S(n7949), .Q(n12456)
         );
  MUX21X1 U14067 ( .IN1(\mem2[255][19] ), .IN2(n1107), .S(n7949), .Q(n12455)
         );
  MUX21X1 U14068 ( .IN1(\mem2[255][18] ), .IN2(n1085), .S(n7949), .Q(n12454)
         );
  MUX21X1 U14069 ( .IN1(\mem2[255][17] ), .IN2(n1063), .S(n7949), .Q(n12453)
         );
  MUX21X1 U14070 ( .IN1(\mem2[255][16] ), .IN2(n1041), .S(n7949), .Q(n12452)
         );
  AND2X1 U14071 ( .IN1(n7950), .IN2(n7099), .Q(n7949) );
  MUX21X1 U14072 ( .IN1(\mem2[254][23] ), .IN2(n1195), .S(n7951), .Q(n12451)
         );
  MUX21X1 U14073 ( .IN1(\mem2[254][22] ), .IN2(n1173), .S(n7951), .Q(n12450)
         );
  MUX21X1 U14074 ( .IN1(\mem2[254][21] ), .IN2(n1151), .S(n7951), .Q(n12449)
         );
  MUX21X1 U14075 ( .IN1(\mem2[254][20] ), .IN2(n1129), .S(n7951), .Q(n12448)
         );
  MUX21X1 U14076 ( .IN1(\mem2[254][19] ), .IN2(n1107), .S(n7951), .Q(n12447)
         );
  MUX21X1 U14077 ( .IN1(\mem2[254][18] ), .IN2(n1085), .S(n7951), .Q(n12446)
         );
  MUX21X1 U14078 ( .IN1(\mem2[254][17] ), .IN2(n1063), .S(n7951), .Q(n12445)
         );
  MUX21X1 U14079 ( .IN1(\mem2[254][16] ), .IN2(n1041), .S(n7951), .Q(n12444)
         );
  AND2X1 U14080 ( .IN1(n7950), .IN2(n7102), .Q(n7951) );
  MUX21X1 U14081 ( .IN1(\mem2[253][23] ), .IN2(n1195), .S(n7952), .Q(n12443)
         );
  MUX21X1 U14082 ( .IN1(\mem2[253][22] ), .IN2(n1173), .S(n7952), .Q(n12442)
         );
  MUX21X1 U14083 ( .IN1(\mem2[253][21] ), .IN2(n1151), .S(n7952), .Q(n12441)
         );
  MUX21X1 U14084 ( .IN1(\mem2[253][20] ), .IN2(n1129), .S(n7952), .Q(n12440)
         );
  MUX21X1 U14085 ( .IN1(\mem2[253][19] ), .IN2(n1107), .S(n7952), .Q(n12439)
         );
  MUX21X1 U14086 ( .IN1(\mem2[253][18] ), .IN2(n1085), .S(n7952), .Q(n12438)
         );
  MUX21X1 U14087 ( .IN1(\mem2[253][17] ), .IN2(n1063), .S(n7952), .Q(n12437)
         );
  MUX21X1 U14088 ( .IN1(\mem2[253][16] ), .IN2(n1041), .S(n7952), .Q(n12436)
         );
  AND2X1 U14089 ( .IN1(n7950), .IN2(n7104), .Q(n7952) );
  MUX21X1 U14090 ( .IN1(\mem2[252][23] ), .IN2(n1195), .S(n7953), .Q(n12435)
         );
  MUX21X1 U14091 ( .IN1(\mem2[252][22] ), .IN2(n1173), .S(n7953), .Q(n12434)
         );
  MUX21X1 U14092 ( .IN1(\mem2[252][21] ), .IN2(n1151), .S(n7953), .Q(n12433)
         );
  MUX21X1 U14093 ( .IN1(\mem2[252][20] ), .IN2(n1129), .S(n7953), .Q(n12432)
         );
  MUX21X1 U14094 ( .IN1(\mem2[252][19] ), .IN2(n1107), .S(n7953), .Q(n12431)
         );
  MUX21X1 U14095 ( .IN1(\mem2[252][18] ), .IN2(n1085), .S(n7953), .Q(n12430)
         );
  MUX21X1 U14096 ( .IN1(\mem2[252][17] ), .IN2(n1063), .S(n7953), .Q(n12429)
         );
  MUX21X1 U14097 ( .IN1(\mem2[252][16] ), .IN2(n1041), .S(n7953), .Q(n12428)
         );
  AND2X1 U14098 ( .IN1(n7950), .IN2(n7106), .Q(n7953) );
  MUX21X1 U14099 ( .IN1(\mem2[251][23] ), .IN2(n1195), .S(n7954), .Q(n12427)
         );
  MUX21X1 U14100 ( .IN1(\mem2[251][22] ), .IN2(n1173), .S(n7954), .Q(n12426)
         );
  MUX21X1 U14101 ( .IN1(\mem2[251][21] ), .IN2(n1151), .S(n7954), .Q(n12425)
         );
  MUX21X1 U14102 ( .IN1(\mem2[251][20] ), .IN2(n1129), .S(n7954), .Q(n12424)
         );
  MUX21X1 U14103 ( .IN1(\mem2[251][19] ), .IN2(n1107), .S(n7954), .Q(n12423)
         );
  MUX21X1 U14104 ( .IN1(\mem2[251][18] ), .IN2(n1085), .S(n7954), .Q(n12422)
         );
  MUX21X1 U14105 ( .IN1(\mem2[251][17] ), .IN2(n1063), .S(n7954), .Q(n12421)
         );
  MUX21X1 U14106 ( .IN1(\mem2[251][16] ), .IN2(n1041), .S(n7954), .Q(n12420)
         );
  AND2X1 U14107 ( .IN1(n7950), .IN2(n7108), .Q(n7954) );
  MUX21X1 U14108 ( .IN1(\mem2[250][23] ), .IN2(n1195), .S(n7955), .Q(n12419)
         );
  MUX21X1 U14109 ( .IN1(\mem2[250][22] ), .IN2(n1173), .S(n7955), .Q(n12418)
         );
  MUX21X1 U14110 ( .IN1(\mem2[250][21] ), .IN2(n1151), .S(n7955), .Q(n12417)
         );
  MUX21X1 U14111 ( .IN1(\mem2[250][20] ), .IN2(n1129), .S(n7955), .Q(n12416)
         );
  MUX21X1 U14112 ( .IN1(\mem2[250][19] ), .IN2(n1107), .S(n7955), .Q(n12415)
         );
  MUX21X1 U14113 ( .IN1(\mem2[250][18] ), .IN2(n1085), .S(n7955), .Q(n12414)
         );
  MUX21X1 U14114 ( .IN1(\mem2[250][17] ), .IN2(n1063), .S(n7955), .Q(n12413)
         );
  MUX21X1 U14115 ( .IN1(\mem2[250][16] ), .IN2(n1041), .S(n7955), .Q(n12412)
         );
  AND2X1 U14116 ( .IN1(n7950), .IN2(n7110), .Q(n7955) );
  MUX21X1 U14117 ( .IN1(\mem2[249][23] ), .IN2(n1195), .S(n7956), .Q(n12411)
         );
  MUX21X1 U14118 ( .IN1(\mem2[249][22] ), .IN2(n1173), .S(n7956), .Q(n12410)
         );
  MUX21X1 U14119 ( .IN1(\mem2[249][21] ), .IN2(n1151), .S(n7956), .Q(n12409)
         );
  MUX21X1 U14120 ( .IN1(\mem2[249][20] ), .IN2(n1129), .S(n7956), .Q(n12408)
         );
  MUX21X1 U14121 ( .IN1(\mem2[249][19] ), .IN2(n1107), .S(n7956), .Q(n12407)
         );
  MUX21X1 U14122 ( .IN1(\mem2[249][18] ), .IN2(n1085), .S(n7956), .Q(n12406)
         );
  MUX21X1 U14123 ( .IN1(\mem2[249][17] ), .IN2(n1063), .S(n7956), .Q(n12405)
         );
  MUX21X1 U14124 ( .IN1(\mem2[249][16] ), .IN2(n1041), .S(n7956), .Q(n12404)
         );
  AND2X1 U14125 ( .IN1(n7950), .IN2(n7112), .Q(n7956) );
  MUX21X1 U14126 ( .IN1(\mem2[248][23] ), .IN2(n1195), .S(n7957), .Q(n12403)
         );
  MUX21X1 U14127 ( .IN1(\mem2[248][22] ), .IN2(n1173), .S(n7957), .Q(n12402)
         );
  MUX21X1 U14128 ( .IN1(\mem2[248][21] ), .IN2(n1151), .S(n7957), .Q(n12401)
         );
  MUX21X1 U14129 ( .IN1(\mem2[248][20] ), .IN2(n1129), .S(n7957), .Q(n12400)
         );
  MUX21X1 U14130 ( .IN1(\mem2[248][19] ), .IN2(n1107), .S(n7957), .Q(n12399)
         );
  MUX21X1 U14131 ( .IN1(\mem2[248][18] ), .IN2(n1085), .S(n7957), .Q(n12398)
         );
  MUX21X1 U14132 ( .IN1(\mem2[248][17] ), .IN2(n1063), .S(n7957), .Q(n12397)
         );
  MUX21X1 U14133 ( .IN1(\mem2[248][16] ), .IN2(n1041), .S(n7957), .Q(n12396)
         );
  AND2X1 U14134 ( .IN1(n7950), .IN2(n7114), .Q(n7957) );
  MUX21X1 U14135 ( .IN1(\mem2[247][23] ), .IN2(n1195), .S(n7958), .Q(n12395)
         );
  MUX21X1 U14136 ( .IN1(\mem2[247][22] ), .IN2(n1173), .S(n7958), .Q(n12394)
         );
  MUX21X1 U14137 ( .IN1(\mem2[247][21] ), .IN2(n1151), .S(n7958), .Q(n12393)
         );
  MUX21X1 U14138 ( .IN1(\mem2[247][20] ), .IN2(n1129), .S(n7958), .Q(n12392)
         );
  MUX21X1 U14139 ( .IN1(\mem2[247][19] ), .IN2(n1107), .S(n7958), .Q(n12391)
         );
  MUX21X1 U14140 ( .IN1(\mem2[247][18] ), .IN2(n1085), .S(n7958), .Q(n12390)
         );
  MUX21X1 U14141 ( .IN1(\mem2[247][17] ), .IN2(n1063), .S(n7958), .Q(n12389)
         );
  MUX21X1 U14142 ( .IN1(\mem2[247][16] ), .IN2(n1041), .S(n7958), .Q(n12388)
         );
  AND2X1 U14143 ( .IN1(n7950), .IN2(n7116), .Q(n7958) );
  MUX21X1 U14144 ( .IN1(\mem2[246][23] ), .IN2(n1195), .S(n7959), .Q(n12387)
         );
  MUX21X1 U14145 ( .IN1(\mem2[246][22] ), .IN2(n1173), .S(n7959), .Q(n12386)
         );
  MUX21X1 U14146 ( .IN1(\mem2[246][21] ), .IN2(n1151), .S(n7959), .Q(n12385)
         );
  MUX21X1 U14147 ( .IN1(\mem2[246][20] ), .IN2(n1129), .S(n7959), .Q(n12384)
         );
  MUX21X1 U14148 ( .IN1(\mem2[246][19] ), .IN2(n1107), .S(n7959), .Q(n12383)
         );
  MUX21X1 U14149 ( .IN1(\mem2[246][18] ), .IN2(n1085), .S(n7959), .Q(n12382)
         );
  MUX21X1 U14150 ( .IN1(\mem2[246][17] ), .IN2(n1063), .S(n7959), .Q(n12381)
         );
  MUX21X1 U14151 ( .IN1(\mem2[246][16] ), .IN2(n1041), .S(n7959), .Q(n12380)
         );
  AND2X1 U14152 ( .IN1(n7950), .IN2(n7118), .Q(n7959) );
  MUX21X1 U14153 ( .IN1(\mem2[245][23] ), .IN2(n1195), .S(n7960), .Q(n12379)
         );
  MUX21X1 U14154 ( .IN1(\mem2[245][22] ), .IN2(n1173), .S(n7960), .Q(n12378)
         );
  MUX21X1 U14155 ( .IN1(\mem2[245][21] ), .IN2(n1151), .S(n7960), .Q(n12377)
         );
  MUX21X1 U14156 ( .IN1(\mem2[245][20] ), .IN2(n1129), .S(n7960), .Q(n12376)
         );
  MUX21X1 U14157 ( .IN1(\mem2[245][19] ), .IN2(n1107), .S(n7960), .Q(n12375)
         );
  MUX21X1 U14158 ( .IN1(\mem2[245][18] ), .IN2(n1085), .S(n7960), .Q(n12374)
         );
  MUX21X1 U14159 ( .IN1(\mem2[245][17] ), .IN2(n1063), .S(n7960), .Q(n12373)
         );
  MUX21X1 U14160 ( .IN1(\mem2[245][16] ), .IN2(n1041), .S(n7960), .Q(n12372)
         );
  AND2X1 U14161 ( .IN1(n7950), .IN2(n7120), .Q(n7960) );
  MUX21X1 U14162 ( .IN1(\mem2[244][23] ), .IN2(n1195), .S(n7961), .Q(n12371)
         );
  MUX21X1 U14163 ( .IN1(\mem2[244][22] ), .IN2(n1173), .S(n7961), .Q(n12370)
         );
  MUX21X1 U14164 ( .IN1(\mem2[244][21] ), .IN2(n1151), .S(n7961), .Q(n12369)
         );
  MUX21X1 U14165 ( .IN1(\mem2[244][20] ), .IN2(n1129), .S(n7961), .Q(n12368)
         );
  MUX21X1 U14166 ( .IN1(\mem2[244][19] ), .IN2(n1107), .S(n7961), .Q(n12367)
         );
  MUX21X1 U14167 ( .IN1(\mem2[244][18] ), .IN2(n1085), .S(n7961), .Q(n12366)
         );
  MUX21X1 U14168 ( .IN1(\mem2[244][17] ), .IN2(n1063), .S(n7961), .Q(n12365)
         );
  MUX21X1 U14169 ( .IN1(\mem2[244][16] ), .IN2(n1041), .S(n7961), .Q(n12364)
         );
  AND2X1 U14170 ( .IN1(n7950), .IN2(n7122), .Q(n7961) );
  MUX21X1 U14171 ( .IN1(\mem2[243][23] ), .IN2(n1196), .S(n7962), .Q(n12363)
         );
  MUX21X1 U14172 ( .IN1(\mem2[243][22] ), .IN2(n1174), .S(n7962), .Q(n12362)
         );
  MUX21X1 U14173 ( .IN1(\mem2[243][21] ), .IN2(n1152), .S(n7962), .Q(n12361)
         );
  MUX21X1 U14174 ( .IN1(\mem2[243][20] ), .IN2(n1130), .S(n7962), .Q(n12360)
         );
  MUX21X1 U14175 ( .IN1(\mem2[243][19] ), .IN2(n1108), .S(n7962), .Q(n12359)
         );
  MUX21X1 U14176 ( .IN1(\mem2[243][18] ), .IN2(n1086), .S(n7962), .Q(n12358)
         );
  MUX21X1 U14177 ( .IN1(\mem2[243][17] ), .IN2(n1064), .S(n7962), .Q(n12357)
         );
  MUX21X1 U14178 ( .IN1(\mem2[243][16] ), .IN2(n1042), .S(n7962), .Q(n12356)
         );
  AND2X1 U14179 ( .IN1(n7950), .IN2(n7124), .Q(n7962) );
  MUX21X1 U14180 ( .IN1(\mem2[242][23] ), .IN2(n1196), .S(n7963), .Q(n12355)
         );
  MUX21X1 U14181 ( .IN1(\mem2[242][22] ), .IN2(n1174), .S(n7963), .Q(n12354)
         );
  MUX21X1 U14182 ( .IN1(\mem2[242][21] ), .IN2(n1152), .S(n7963), .Q(n12353)
         );
  MUX21X1 U14183 ( .IN1(\mem2[242][20] ), .IN2(n1130), .S(n7963), .Q(n12352)
         );
  MUX21X1 U14184 ( .IN1(\mem2[242][19] ), .IN2(n1108), .S(n7963), .Q(n12351)
         );
  MUX21X1 U14185 ( .IN1(\mem2[242][18] ), .IN2(n1086), .S(n7963), .Q(n12350)
         );
  MUX21X1 U14186 ( .IN1(\mem2[242][17] ), .IN2(n1064), .S(n7963), .Q(n12349)
         );
  MUX21X1 U14187 ( .IN1(\mem2[242][16] ), .IN2(n1042), .S(n7963), .Q(n12348)
         );
  AND2X1 U14188 ( .IN1(n7950), .IN2(n7126), .Q(n7963) );
  MUX21X1 U14189 ( .IN1(\mem2[241][23] ), .IN2(n1196), .S(n7964), .Q(n12347)
         );
  MUX21X1 U14190 ( .IN1(\mem2[241][22] ), .IN2(n1174), .S(n7964), .Q(n12346)
         );
  MUX21X1 U14191 ( .IN1(\mem2[241][21] ), .IN2(n1152), .S(n7964), .Q(n12345)
         );
  MUX21X1 U14192 ( .IN1(\mem2[241][20] ), .IN2(n1130), .S(n7964), .Q(n12344)
         );
  MUX21X1 U14193 ( .IN1(\mem2[241][19] ), .IN2(n1108), .S(n7964), .Q(n12343)
         );
  MUX21X1 U14194 ( .IN1(\mem2[241][18] ), .IN2(n1086), .S(n7964), .Q(n12342)
         );
  MUX21X1 U14195 ( .IN1(\mem2[241][17] ), .IN2(n1064), .S(n7964), .Q(n12341)
         );
  MUX21X1 U14196 ( .IN1(\mem2[241][16] ), .IN2(n1042), .S(n7964), .Q(n12340)
         );
  AND2X1 U14197 ( .IN1(n7950), .IN2(n7128), .Q(n7964) );
  MUX21X1 U14198 ( .IN1(\mem2[240][23] ), .IN2(n1196), .S(n7965), .Q(n12339)
         );
  MUX21X1 U14199 ( .IN1(\mem2[240][22] ), .IN2(n1174), .S(n7965), .Q(n12338)
         );
  MUX21X1 U14200 ( .IN1(\mem2[240][21] ), .IN2(n1152), .S(n7965), .Q(n12337)
         );
  MUX21X1 U14201 ( .IN1(\mem2[240][20] ), .IN2(n1130), .S(n7965), .Q(n12336)
         );
  MUX21X1 U14202 ( .IN1(\mem2[240][19] ), .IN2(n1108), .S(n7965), .Q(n12335)
         );
  MUX21X1 U14203 ( .IN1(\mem2[240][18] ), .IN2(n1086), .S(n7965), .Q(n12334)
         );
  MUX21X1 U14204 ( .IN1(\mem2[240][17] ), .IN2(n1064), .S(n7965), .Q(n12333)
         );
  MUX21X1 U14205 ( .IN1(\mem2[240][16] ), .IN2(n1042), .S(n7965), .Q(n12332)
         );
  AND2X1 U14206 ( .IN1(n7950), .IN2(n7130), .Q(n7965) );
  AND2X1 U14207 ( .IN1(n7966), .IN2(n7131), .Q(n7950) );
  AND2X1 U14208 ( .IN1(n7967), .IN2(n7968), .Q(n7131) );
  MUX21X1 U14209 ( .IN1(\mem2[239][23] ), .IN2(n1196), .S(n7969), .Q(n12331)
         );
  MUX21X1 U14210 ( .IN1(\mem2[239][22] ), .IN2(n1174), .S(n7969), .Q(n12330)
         );
  MUX21X1 U14211 ( .IN1(\mem2[239][21] ), .IN2(n1152), .S(n7969), .Q(n12329)
         );
  MUX21X1 U14212 ( .IN1(\mem2[239][20] ), .IN2(n1130), .S(n7969), .Q(n12328)
         );
  MUX21X1 U14213 ( .IN1(\mem2[239][19] ), .IN2(n1108), .S(n7969), .Q(n12327)
         );
  MUX21X1 U14214 ( .IN1(\mem2[239][18] ), .IN2(n1086), .S(n7969), .Q(n12326)
         );
  MUX21X1 U14215 ( .IN1(\mem2[239][17] ), .IN2(n1064), .S(n7969), .Q(n12325)
         );
  MUX21X1 U14216 ( .IN1(\mem2[239][16] ), .IN2(n1042), .S(n7969), .Q(n12324)
         );
  AND2X1 U14217 ( .IN1(n7970), .IN2(n7099), .Q(n7969) );
  MUX21X1 U14218 ( .IN1(\mem2[238][23] ), .IN2(n1196), .S(n7971), .Q(n12323)
         );
  MUX21X1 U14219 ( .IN1(\mem2[238][22] ), .IN2(n1174), .S(n7971), .Q(n12322)
         );
  MUX21X1 U14220 ( .IN1(\mem2[238][21] ), .IN2(n1152), .S(n7971), .Q(n12321)
         );
  MUX21X1 U14221 ( .IN1(\mem2[238][20] ), .IN2(n1130), .S(n7971), .Q(n12320)
         );
  MUX21X1 U14222 ( .IN1(\mem2[238][19] ), .IN2(n1108), .S(n7971), .Q(n12319)
         );
  MUX21X1 U14223 ( .IN1(\mem2[238][18] ), .IN2(n1086), .S(n7971), .Q(n12318)
         );
  MUX21X1 U14224 ( .IN1(\mem2[238][17] ), .IN2(n1064), .S(n7971), .Q(n12317)
         );
  MUX21X1 U14225 ( .IN1(\mem2[238][16] ), .IN2(n1042), .S(n7971), .Q(n12316)
         );
  AND2X1 U14226 ( .IN1(n7970), .IN2(n7102), .Q(n7971) );
  MUX21X1 U14227 ( .IN1(\mem2[237][23] ), .IN2(n1196), .S(n7972), .Q(n12315)
         );
  MUX21X1 U14228 ( .IN1(\mem2[237][22] ), .IN2(n1174), .S(n7972), .Q(n12314)
         );
  MUX21X1 U14229 ( .IN1(\mem2[237][21] ), .IN2(n1152), .S(n7972), .Q(n12313)
         );
  MUX21X1 U14230 ( .IN1(\mem2[237][20] ), .IN2(n1130), .S(n7972), .Q(n12312)
         );
  MUX21X1 U14231 ( .IN1(\mem2[237][19] ), .IN2(n1108), .S(n7972), .Q(n12311)
         );
  MUX21X1 U14232 ( .IN1(\mem2[237][18] ), .IN2(n1086), .S(n7972), .Q(n12310)
         );
  MUX21X1 U14233 ( .IN1(\mem2[237][17] ), .IN2(n1064), .S(n7972), .Q(n12309)
         );
  MUX21X1 U14234 ( .IN1(\mem2[237][16] ), .IN2(n1042), .S(n7972), .Q(n12308)
         );
  AND2X1 U14235 ( .IN1(n7970), .IN2(n7104), .Q(n7972) );
  MUX21X1 U14236 ( .IN1(\mem2[236][23] ), .IN2(n1196), .S(n7973), .Q(n12307)
         );
  MUX21X1 U14237 ( .IN1(\mem2[236][22] ), .IN2(n1174), .S(n7973), .Q(n12306)
         );
  MUX21X1 U14238 ( .IN1(\mem2[236][21] ), .IN2(n1152), .S(n7973), .Q(n12305)
         );
  MUX21X1 U14239 ( .IN1(\mem2[236][20] ), .IN2(n1130), .S(n7973), .Q(n12304)
         );
  MUX21X1 U14240 ( .IN1(\mem2[236][19] ), .IN2(n1108), .S(n7973), .Q(n12303)
         );
  MUX21X1 U14241 ( .IN1(\mem2[236][18] ), .IN2(n1086), .S(n7973), .Q(n12302)
         );
  MUX21X1 U14242 ( .IN1(\mem2[236][17] ), .IN2(n1064), .S(n7973), .Q(n12301)
         );
  MUX21X1 U14243 ( .IN1(\mem2[236][16] ), .IN2(n1042), .S(n7973), .Q(n12300)
         );
  AND2X1 U14244 ( .IN1(n7970), .IN2(n7106), .Q(n7973) );
  MUX21X1 U14245 ( .IN1(\mem2[235][23] ), .IN2(n1196), .S(n7974), .Q(n12299)
         );
  MUX21X1 U14246 ( .IN1(\mem2[235][22] ), .IN2(n1174), .S(n7974), .Q(n12298)
         );
  MUX21X1 U14247 ( .IN1(\mem2[235][21] ), .IN2(n1152), .S(n7974), .Q(n12297)
         );
  MUX21X1 U14248 ( .IN1(\mem2[235][20] ), .IN2(n1130), .S(n7974), .Q(n12296)
         );
  MUX21X1 U14249 ( .IN1(\mem2[235][19] ), .IN2(n1108), .S(n7974), .Q(n12295)
         );
  MUX21X1 U14250 ( .IN1(\mem2[235][18] ), .IN2(n1086), .S(n7974), .Q(n12294)
         );
  MUX21X1 U14251 ( .IN1(\mem2[235][17] ), .IN2(n1064), .S(n7974), .Q(n12293)
         );
  MUX21X1 U14252 ( .IN1(\mem2[235][16] ), .IN2(n1042), .S(n7974), .Q(n12292)
         );
  AND2X1 U14253 ( .IN1(n7970), .IN2(n7108), .Q(n7974) );
  MUX21X1 U14254 ( .IN1(\mem2[234][23] ), .IN2(n1196), .S(n7975), .Q(n12291)
         );
  MUX21X1 U14255 ( .IN1(\mem2[234][22] ), .IN2(n1174), .S(n7975), .Q(n12290)
         );
  MUX21X1 U14256 ( .IN1(\mem2[234][21] ), .IN2(n1152), .S(n7975), .Q(n12289)
         );
  MUX21X1 U14257 ( .IN1(\mem2[234][20] ), .IN2(n1130), .S(n7975), .Q(n12288)
         );
  MUX21X1 U14258 ( .IN1(\mem2[234][19] ), .IN2(n1108), .S(n7975), .Q(n12287)
         );
  MUX21X1 U14259 ( .IN1(\mem2[234][18] ), .IN2(n1086), .S(n7975), .Q(n12286)
         );
  MUX21X1 U14260 ( .IN1(\mem2[234][17] ), .IN2(n1064), .S(n7975), .Q(n12285)
         );
  MUX21X1 U14261 ( .IN1(\mem2[234][16] ), .IN2(n1042), .S(n7975), .Q(n12284)
         );
  AND2X1 U14262 ( .IN1(n7970), .IN2(n7110), .Q(n7975) );
  MUX21X1 U14263 ( .IN1(\mem2[233][23] ), .IN2(n1196), .S(n7976), .Q(n12283)
         );
  MUX21X1 U14264 ( .IN1(\mem2[233][22] ), .IN2(n1174), .S(n7976), .Q(n12282)
         );
  MUX21X1 U14265 ( .IN1(\mem2[233][21] ), .IN2(n1152), .S(n7976), .Q(n12281)
         );
  MUX21X1 U14266 ( .IN1(\mem2[233][20] ), .IN2(n1130), .S(n7976), .Q(n12280)
         );
  MUX21X1 U14267 ( .IN1(\mem2[233][19] ), .IN2(n1108), .S(n7976), .Q(n12279)
         );
  MUX21X1 U14268 ( .IN1(\mem2[233][18] ), .IN2(n1086), .S(n7976), .Q(n12278)
         );
  MUX21X1 U14269 ( .IN1(\mem2[233][17] ), .IN2(n1064), .S(n7976), .Q(n12277)
         );
  MUX21X1 U14270 ( .IN1(\mem2[233][16] ), .IN2(n1042), .S(n7976), .Q(n12276)
         );
  AND2X1 U14271 ( .IN1(n7970), .IN2(n7112), .Q(n7976) );
  MUX21X1 U14272 ( .IN1(\mem2[232][23] ), .IN2(n1196), .S(n7977), .Q(n12275)
         );
  MUX21X1 U14273 ( .IN1(\mem2[232][22] ), .IN2(n1174), .S(n7977), .Q(n12274)
         );
  MUX21X1 U14274 ( .IN1(\mem2[232][21] ), .IN2(n1152), .S(n7977), .Q(n12273)
         );
  MUX21X1 U14275 ( .IN1(\mem2[232][20] ), .IN2(n1130), .S(n7977), .Q(n12272)
         );
  MUX21X1 U14276 ( .IN1(\mem2[232][19] ), .IN2(n1108), .S(n7977), .Q(n12271)
         );
  MUX21X1 U14277 ( .IN1(\mem2[232][18] ), .IN2(n1086), .S(n7977), .Q(n12270)
         );
  MUX21X1 U14278 ( .IN1(\mem2[232][17] ), .IN2(n1064), .S(n7977), .Q(n12269)
         );
  MUX21X1 U14279 ( .IN1(\mem2[232][16] ), .IN2(n1042), .S(n7977), .Q(n12268)
         );
  AND2X1 U14280 ( .IN1(n7970), .IN2(n7114), .Q(n7977) );
  MUX21X1 U14281 ( .IN1(\mem2[231][23] ), .IN2(n1197), .S(n7978), .Q(n12267)
         );
  MUX21X1 U14282 ( .IN1(\mem2[231][22] ), .IN2(n1175), .S(n7978), .Q(n12266)
         );
  MUX21X1 U14283 ( .IN1(\mem2[231][21] ), .IN2(n1153), .S(n7978), .Q(n12265)
         );
  MUX21X1 U14284 ( .IN1(\mem2[231][20] ), .IN2(n1131), .S(n7978), .Q(n12264)
         );
  MUX21X1 U14285 ( .IN1(\mem2[231][19] ), .IN2(n1109), .S(n7978), .Q(n12263)
         );
  MUX21X1 U14286 ( .IN1(\mem2[231][18] ), .IN2(n1087), .S(n7978), .Q(n12262)
         );
  MUX21X1 U14287 ( .IN1(\mem2[231][17] ), .IN2(n1065), .S(n7978), .Q(n12261)
         );
  MUX21X1 U14288 ( .IN1(\mem2[231][16] ), .IN2(n1043), .S(n7978), .Q(n12260)
         );
  AND2X1 U14289 ( .IN1(n7970), .IN2(n7116), .Q(n7978) );
  MUX21X1 U14290 ( .IN1(\mem2[230][23] ), .IN2(n1197), .S(n7979), .Q(n12259)
         );
  MUX21X1 U14291 ( .IN1(\mem2[230][22] ), .IN2(n1175), .S(n7979), .Q(n12258)
         );
  MUX21X1 U14292 ( .IN1(\mem2[230][21] ), .IN2(n1153), .S(n7979), .Q(n12257)
         );
  MUX21X1 U14293 ( .IN1(\mem2[230][20] ), .IN2(n1131), .S(n7979), .Q(n12256)
         );
  MUX21X1 U14294 ( .IN1(\mem2[230][19] ), .IN2(n1109), .S(n7979), .Q(n12255)
         );
  MUX21X1 U14295 ( .IN1(\mem2[230][18] ), .IN2(n1087), .S(n7979), .Q(n12254)
         );
  MUX21X1 U14296 ( .IN1(\mem2[230][17] ), .IN2(n1065), .S(n7979), .Q(n12253)
         );
  MUX21X1 U14297 ( .IN1(\mem2[230][16] ), .IN2(n1043), .S(n7979), .Q(n12252)
         );
  AND2X1 U14298 ( .IN1(n7970), .IN2(n7118), .Q(n7979) );
  MUX21X1 U14299 ( .IN1(\mem2[229][23] ), .IN2(n1197), .S(n7980), .Q(n12251)
         );
  MUX21X1 U14300 ( .IN1(\mem2[229][22] ), .IN2(n1175), .S(n7980), .Q(n12250)
         );
  MUX21X1 U14301 ( .IN1(\mem2[229][21] ), .IN2(n1153), .S(n7980), .Q(n12249)
         );
  MUX21X1 U14302 ( .IN1(\mem2[229][20] ), .IN2(n1131), .S(n7980), .Q(n12248)
         );
  MUX21X1 U14303 ( .IN1(\mem2[229][19] ), .IN2(n1109), .S(n7980), .Q(n12247)
         );
  MUX21X1 U14304 ( .IN1(\mem2[229][18] ), .IN2(n1087), .S(n7980), .Q(n12246)
         );
  MUX21X1 U14305 ( .IN1(\mem2[229][17] ), .IN2(n1065), .S(n7980), .Q(n12245)
         );
  MUX21X1 U14306 ( .IN1(\mem2[229][16] ), .IN2(n1043), .S(n7980), .Q(n12244)
         );
  AND2X1 U14307 ( .IN1(n7970), .IN2(n7120), .Q(n7980) );
  MUX21X1 U14308 ( .IN1(\mem2[228][23] ), .IN2(n1197), .S(n7981), .Q(n12243)
         );
  MUX21X1 U14309 ( .IN1(\mem2[228][22] ), .IN2(n1175), .S(n7981), .Q(n12242)
         );
  MUX21X1 U14310 ( .IN1(\mem2[228][21] ), .IN2(n1153), .S(n7981), .Q(n12241)
         );
  MUX21X1 U14311 ( .IN1(\mem2[228][20] ), .IN2(n1131), .S(n7981), .Q(n12240)
         );
  MUX21X1 U14312 ( .IN1(\mem2[228][19] ), .IN2(n1109), .S(n7981), .Q(n12239)
         );
  MUX21X1 U14313 ( .IN1(\mem2[228][18] ), .IN2(n1087), .S(n7981), .Q(n12238)
         );
  MUX21X1 U14314 ( .IN1(\mem2[228][17] ), .IN2(n1065), .S(n7981), .Q(n12237)
         );
  MUX21X1 U14315 ( .IN1(\mem2[228][16] ), .IN2(n1043), .S(n7981), .Q(n12236)
         );
  AND2X1 U14316 ( .IN1(n7970), .IN2(n7122), .Q(n7981) );
  MUX21X1 U14317 ( .IN1(\mem2[227][23] ), .IN2(n1197), .S(n7982), .Q(n12235)
         );
  MUX21X1 U14318 ( .IN1(\mem2[227][22] ), .IN2(n1175), .S(n7982), .Q(n12234)
         );
  MUX21X1 U14319 ( .IN1(\mem2[227][21] ), .IN2(n1153), .S(n7982), .Q(n12233)
         );
  MUX21X1 U14320 ( .IN1(\mem2[227][20] ), .IN2(n1131), .S(n7982), .Q(n12232)
         );
  MUX21X1 U14321 ( .IN1(\mem2[227][19] ), .IN2(n1109), .S(n7982), .Q(n12231)
         );
  MUX21X1 U14322 ( .IN1(\mem2[227][18] ), .IN2(n1087), .S(n7982), .Q(n12230)
         );
  MUX21X1 U14323 ( .IN1(\mem2[227][17] ), .IN2(n1065), .S(n7982), .Q(n12229)
         );
  MUX21X1 U14324 ( .IN1(\mem2[227][16] ), .IN2(n1043), .S(n7982), .Q(n12228)
         );
  AND2X1 U14325 ( .IN1(n7970), .IN2(n7124), .Q(n7982) );
  MUX21X1 U14326 ( .IN1(\mem2[226][23] ), .IN2(n1197), .S(n7983), .Q(n12227)
         );
  MUX21X1 U14327 ( .IN1(\mem2[226][22] ), .IN2(n1175), .S(n7983), .Q(n12226)
         );
  MUX21X1 U14328 ( .IN1(\mem2[226][21] ), .IN2(n1153), .S(n7983), .Q(n12225)
         );
  MUX21X1 U14329 ( .IN1(\mem2[226][20] ), .IN2(n1131), .S(n7983), .Q(n12224)
         );
  MUX21X1 U14330 ( .IN1(\mem2[226][19] ), .IN2(n1109), .S(n7983), .Q(n12223)
         );
  MUX21X1 U14331 ( .IN1(\mem2[226][18] ), .IN2(n1087), .S(n7983), .Q(n12222)
         );
  MUX21X1 U14332 ( .IN1(\mem2[226][17] ), .IN2(n1065), .S(n7983), .Q(n12221)
         );
  MUX21X1 U14333 ( .IN1(\mem2[226][16] ), .IN2(n1043), .S(n7983), .Q(n12220)
         );
  AND2X1 U14334 ( .IN1(n7970), .IN2(n7126), .Q(n7983) );
  MUX21X1 U14335 ( .IN1(\mem2[225][23] ), .IN2(n1197), .S(n7984), .Q(n12219)
         );
  MUX21X1 U14336 ( .IN1(\mem2[225][22] ), .IN2(n1175), .S(n7984), .Q(n12218)
         );
  MUX21X1 U14337 ( .IN1(\mem2[225][21] ), .IN2(n1153), .S(n7984), .Q(n12217)
         );
  MUX21X1 U14338 ( .IN1(\mem2[225][20] ), .IN2(n1131), .S(n7984), .Q(n12216)
         );
  MUX21X1 U14339 ( .IN1(\mem2[225][19] ), .IN2(n1109), .S(n7984), .Q(n12215)
         );
  MUX21X1 U14340 ( .IN1(\mem2[225][18] ), .IN2(n1087), .S(n7984), .Q(n12214)
         );
  MUX21X1 U14341 ( .IN1(\mem2[225][17] ), .IN2(n1065), .S(n7984), .Q(n12213)
         );
  MUX21X1 U14342 ( .IN1(\mem2[225][16] ), .IN2(n1043), .S(n7984), .Q(n12212)
         );
  AND2X1 U14343 ( .IN1(n7970), .IN2(n7128), .Q(n7984) );
  MUX21X1 U14344 ( .IN1(\mem2[224][23] ), .IN2(n1197), .S(n7985), .Q(n12211)
         );
  MUX21X1 U14345 ( .IN1(\mem2[224][22] ), .IN2(n1175), .S(n7985), .Q(n12210)
         );
  MUX21X1 U14346 ( .IN1(\mem2[224][21] ), .IN2(n1153), .S(n7985), .Q(n12209)
         );
  MUX21X1 U14347 ( .IN1(\mem2[224][20] ), .IN2(n1131), .S(n7985), .Q(n12208)
         );
  MUX21X1 U14348 ( .IN1(\mem2[224][19] ), .IN2(n1109), .S(n7985), .Q(n12207)
         );
  MUX21X1 U14349 ( .IN1(\mem2[224][18] ), .IN2(n1087), .S(n7985), .Q(n12206)
         );
  MUX21X1 U14350 ( .IN1(\mem2[224][17] ), .IN2(n1065), .S(n7985), .Q(n12205)
         );
  MUX21X1 U14351 ( .IN1(\mem2[224][16] ), .IN2(n1043), .S(n7985), .Q(n12204)
         );
  AND2X1 U14352 ( .IN1(n7970), .IN2(n7130), .Q(n7985) );
  AND2X1 U14353 ( .IN1(n7966), .IN2(n7150), .Q(n7970) );
  AND2X1 U14354 ( .IN1(n7986), .IN2(n7967), .Q(n7150) );
  MUX21X1 U14355 ( .IN1(\mem2[223][23] ), .IN2(n1197), .S(n7987), .Q(n12203)
         );
  MUX21X1 U14356 ( .IN1(\mem2[223][22] ), .IN2(n1175), .S(n7987), .Q(n12202)
         );
  MUX21X1 U14357 ( .IN1(\mem2[223][21] ), .IN2(n1153), .S(n7987), .Q(n12201)
         );
  MUX21X1 U14358 ( .IN1(\mem2[223][20] ), .IN2(n1131), .S(n7987), .Q(n12200)
         );
  MUX21X1 U14359 ( .IN1(\mem2[223][19] ), .IN2(n1109), .S(n7987), .Q(n12199)
         );
  MUX21X1 U14360 ( .IN1(\mem2[223][18] ), .IN2(n1087), .S(n7987), .Q(n12198)
         );
  MUX21X1 U14361 ( .IN1(\mem2[223][17] ), .IN2(n1065), .S(n7987), .Q(n12197)
         );
  MUX21X1 U14362 ( .IN1(\mem2[223][16] ), .IN2(n1043), .S(n7987), .Q(n12196)
         );
  AND2X1 U14363 ( .IN1(n7988), .IN2(n7099), .Q(n7987) );
  MUX21X1 U14364 ( .IN1(\mem2[222][23] ), .IN2(n1197), .S(n7989), .Q(n12195)
         );
  MUX21X1 U14365 ( .IN1(\mem2[222][22] ), .IN2(n1175), .S(n7989), .Q(n12194)
         );
  MUX21X1 U14366 ( .IN1(\mem2[222][21] ), .IN2(n1153), .S(n7989), .Q(n12193)
         );
  MUX21X1 U14367 ( .IN1(\mem2[222][20] ), .IN2(n1131), .S(n7989), .Q(n12192)
         );
  MUX21X1 U14368 ( .IN1(\mem2[222][19] ), .IN2(n1109), .S(n7989), .Q(n12191)
         );
  MUX21X1 U14369 ( .IN1(\mem2[222][18] ), .IN2(n1087), .S(n7989), .Q(n12190)
         );
  MUX21X1 U14370 ( .IN1(\mem2[222][17] ), .IN2(n1065), .S(n7989), .Q(n12189)
         );
  MUX21X1 U14371 ( .IN1(\mem2[222][16] ), .IN2(n1043), .S(n7989), .Q(n12188)
         );
  AND2X1 U14372 ( .IN1(n7988), .IN2(n7102), .Q(n7989) );
  MUX21X1 U14373 ( .IN1(\mem2[221][23] ), .IN2(n1197), .S(n7990), .Q(n12187)
         );
  MUX21X1 U14374 ( .IN1(\mem2[221][22] ), .IN2(n1175), .S(n7990), .Q(n12186)
         );
  MUX21X1 U14375 ( .IN1(\mem2[221][21] ), .IN2(n1153), .S(n7990), .Q(n12185)
         );
  MUX21X1 U14376 ( .IN1(\mem2[221][20] ), .IN2(n1131), .S(n7990), .Q(n12184)
         );
  MUX21X1 U14377 ( .IN1(\mem2[221][19] ), .IN2(n1109), .S(n7990), .Q(n12183)
         );
  MUX21X1 U14378 ( .IN1(\mem2[221][18] ), .IN2(n1087), .S(n7990), .Q(n12182)
         );
  MUX21X1 U14379 ( .IN1(\mem2[221][17] ), .IN2(n1065), .S(n7990), .Q(n12181)
         );
  MUX21X1 U14380 ( .IN1(\mem2[221][16] ), .IN2(n1043), .S(n7990), .Q(n12180)
         );
  AND2X1 U14381 ( .IN1(n7988), .IN2(n7104), .Q(n7990) );
  MUX21X1 U14382 ( .IN1(\mem2[220][23] ), .IN2(n1197), .S(n7991), .Q(n12179)
         );
  MUX21X1 U14383 ( .IN1(\mem2[220][22] ), .IN2(n1175), .S(n7991), .Q(n12178)
         );
  MUX21X1 U14384 ( .IN1(\mem2[220][21] ), .IN2(n1153), .S(n7991), .Q(n12177)
         );
  MUX21X1 U14385 ( .IN1(\mem2[220][20] ), .IN2(n1131), .S(n7991), .Q(n12176)
         );
  MUX21X1 U14386 ( .IN1(\mem2[220][19] ), .IN2(n1109), .S(n7991), .Q(n12175)
         );
  MUX21X1 U14387 ( .IN1(\mem2[220][18] ), .IN2(n1087), .S(n7991), .Q(n12174)
         );
  MUX21X1 U14388 ( .IN1(\mem2[220][17] ), .IN2(n1065), .S(n7991), .Q(n12173)
         );
  MUX21X1 U14389 ( .IN1(\mem2[220][16] ), .IN2(n1043), .S(n7991), .Q(n12172)
         );
  AND2X1 U14390 ( .IN1(n7988), .IN2(n7106), .Q(n7991) );
  MUX21X1 U14391 ( .IN1(\mem2[219][23] ), .IN2(n1198), .S(n7992), .Q(n12171)
         );
  MUX21X1 U14392 ( .IN1(\mem2[219][22] ), .IN2(n1176), .S(n7992), .Q(n12170)
         );
  MUX21X1 U14393 ( .IN1(\mem2[219][21] ), .IN2(n1154), .S(n7992), .Q(n12169)
         );
  MUX21X1 U14394 ( .IN1(\mem2[219][20] ), .IN2(n1132), .S(n7992), .Q(n12168)
         );
  MUX21X1 U14395 ( .IN1(\mem2[219][19] ), .IN2(n1110), .S(n7992), .Q(n12167)
         );
  MUX21X1 U14396 ( .IN1(\mem2[219][18] ), .IN2(n1088), .S(n7992), .Q(n12166)
         );
  MUX21X1 U14397 ( .IN1(\mem2[219][17] ), .IN2(n1066), .S(n7992), .Q(n12165)
         );
  MUX21X1 U14398 ( .IN1(\mem2[219][16] ), .IN2(n1044), .S(n7992), .Q(n12164)
         );
  AND2X1 U14399 ( .IN1(n7988), .IN2(n7108), .Q(n7992) );
  MUX21X1 U14400 ( .IN1(\mem2[218][23] ), .IN2(n1198), .S(n7993), .Q(n12163)
         );
  MUX21X1 U14401 ( .IN1(\mem2[218][22] ), .IN2(n1176), .S(n7993), .Q(n12162)
         );
  MUX21X1 U14402 ( .IN1(\mem2[218][21] ), .IN2(n1154), .S(n7993), .Q(n12161)
         );
  MUX21X1 U14403 ( .IN1(\mem2[218][20] ), .IN2(n1132), .S(n7993), .Q(n12160)
         );
  MUX21X1 U14404 ( .IN1(\mem2[218][19] ), .IN2(n1110), .S(n7993), .Q(n12159)
         );
  MUX21X1 U14405 ( .IN1(\mem2[218][18] ), .IN2(n1088), .S(n7993), .Q(n12158)
         );
  MUX21X1 U14406 ( .IN1(\mem2[218][17] ), .IN2(n1066), .S(n7993), .Q(n12157)
         );
  MUX21X1 U14407 ( .IN1(\mem2[218][16] ), .IN2(n1044), .S(n7993), .Q(n12156)
         );
  AND2X1 U14408 ( .IN1(n7988), .IN2(n7110), .Q(n7993) );
  MUX21X1 U14409 ( .IN1(\mem2[217][23] ), .IN2(n1198), .S(n7994), .Q(n12155)
         );
  MUX21X1 U14410 ( .IN1(\mem2[217][22] ), .IN2(n1176), .S(n7994), .Q(n12154)
         );
  MUX21X1 U14411 ( .IN1(\mem2[217][21] ), .IN2(n1154), .S(n7994), .Q(n12153)
         );
  MUX21X1 U14412 ( .IN1(\mem2[217][20] ), .IN2(n1132), .S(n7994), .Q(n12152)
         );
  MUX21X1 U14413 ( .IN1(\mem2[217][19] ), .IN2(n1110), .S(n7994), .Q(n12151)
         );
  MUX21X1 U14414 ( .IN1(\mem2[217][18] ), .IN2(n1088), .S(n7994), .Q(n12150)
         );
  MUX21X1 U14415 ( .IN1(\mem2[217][17] ), .IN2(n1066), .S(n7994), .Q(n12149)
         );
  MUX21X1 U14416 ( .IN1(\mem2[217][16] ), .IN2(n1044), .S(n7994), .Q(n12148)
         );
  AND2X1 U14417 ( .IN1(n7988), .IN2(n7112), .Q(n7994) );
  MUX21X1 U14418 ( .IN1(\mem2[216][23] ), .IN2(n1198), .S(n7995), .Q(n12147)
         );
  MUX21X1 U14419 ( .IN1(\mem2[216][22] ), .IN2(n1176), .S(n7995), .Q(n12146)
         );
  MUX21X1 U14420 ( .IN1(\mem2[216][21] ), .IN2(n1154), .S(n7995), .Q(n12145)
         );
  MUX21X1 U14421 ( .IN1(\mem2[216][20] ), .IN2(n1132), .S(n7995), .Q(n12144)
         );
  MUX21X1 U14422 ( .IN1(\mem2[216][19] ), .IN2(n1110), .S(n7995), .Q(n12143)
         );
  MUX21X1 U14423 ( .IN1(\mem2[216][18] ), .IN2(n1088), .S(n7995), .Q(n12142)
         );
  MUX21X1 U14424 ( .IN1(\mem2[216][17] ), .IN2(n1066), .S(n7995), .Q(n12141)
         );
  MUX21X1 U14425 ( .IN1(\mem2[216][16] ), .IN2(n1044), .S(n7995), .Q(n12140)
         );
  AND2X1 U14426 ( .IN1(n7988), .IN2(n7114), .Q(n7995) );
  MUX21X1 U14427 ( .IN1(\mem2[215][23] ), .IN2(n1198), .S(n7996), .Q(n12139)
         );
  MUX21X1 U14428 ( .IN1(\mem2[215][22] ), .IN2(n1176), .S(n7996), .Q(n12138)
         );
  MUX21X1 U14429 ( .IN1(\mem2[215][21] ), .IN2(n1154), .S(n7996), .Q(n12137)
         );
  MUX21X1 U14430 ( .IN1(\mem2[215][20] ), .IN2(n1132), .S(n7996), .Q(n12136)
         );
  MUX21X1 U14431 ( .IN1(\mem2[215][19] ), .IN2(n1110), .S(n7996), .Q(n12135)
         );
  MUX21X1 U14432 ( .IN1(\mem2[215][18] ), .IN2(n1088), .S(n7996), .Q(n12134)
         );
  MUX21X1 U14433 ( .IN1(\mem2[215][17] ), .IN2(n1066), .S(n7996), .Q(n12133)
         );
  MUX21X1 U14434 ( .IN1(\mem2[215][16] ), .IN2(n1044), .S(n7996), .Q(n12132)
         );
  AND2X1 U14435 ( .IN1(n7988), .IN2(n7116), .Q(n7996) );
  MUX21X1 U14436 ( .IN1(\mem2[214][23] ), .IN2(n1198), .S(n7997), .Q(n12131)
         );
  MUX21X1 U14437 ( .IN1(\mem2[214][22] ), .IN2(n1176), .S(n7997), .Q(n12130)
         );
  MUX21X1 U14438 ( .IN1(\mem2[214][21] ), .IN2(n1154), .S(n7997), .Q(n12129)
         );
  MUX21X1 U14439 ( .IN1(\mem2[214][20] ), .IN2(n1132), .S(n7997), .Q(n12128)
         );
  MUX21X1 U14440 ( .IN1(\mem2[214][19] ), .IN2(n1110), .S(n7997), .Q(n12127)
         );
  MUX21X1 U14441 ( .IN1(\mem2[214][18] ), .IN2(n1088), .S(n7997), .Q(n12126)
         );
  MUX21X1 U14442 ( .IN1(\mem2[214][17] ), .IN2(n1066), .S(n7997), .Q(n12125)
         );
  MUX21X1 U14443 ( .IN1(\mem2[214][16] ), .IN2(n1044), .S(n7997), .Q(n12124)
         );
  AND2X1 U14444 ( .IN1(n7988), .IN2(n7118), .Q(n7997) );
  MUX21X1 U14445 ( .IN1(\mem2[213][23] ), .IN2(n1198), .S(n7998), .Q(n12123)
         );
  MUX21X1 U14446 ( .IN1(\mem2[213][22] ), .IN2(n1176), .S(n7998), .Q(n12122)
         );
  MUX21X1 U14447 ( .IN1(\mem2[213][21] ), .IN2(n1154), .S(n7998), .Q(n12121)
         );
  MUX21X1 U14448 ( .IN1(\mem2[213][20] ), .IN2(n1132), .S(n7998), .Q(n12120)
         );
  MUX21X1 U14449 ( .IN1(\mem2[213][19] ), .IN2(n1110), .S(n7998), .Q(n12119)
         );
  MUX21X1 U14450 ( .IN1(\mem2[213][18] ), .IN2(n1088), .S(n7998), .Q(n12118)
         );
  MUX21X1 U14451 ( .IN1(\mem2[213][17] ), .IN2(n1066), .S(n7998), .Q(n12117)
         );
  MUX21X1 U14452 ( .IN1(\mem2[213][16] ), .IN2(n1044), .S(n7998), .Q(n12116)
         );
  AND2X1 U14453 ( .IN1(n7988), .IN2(n7120), .Q(n7998) );
  MUX21X1 U14454 ( .IN1(\mem2[212][23] ), .IN2(n1198), .S(n7999), .Q(n12115)
         );
  MUX21X1 U14455 ( .IN1(\mem2[212][22] ), .IN2(n1176), .S(n7999), .Q(n12114)
         );
  MUX21X1 U14456 ( .IN1(\mem2[212][21] ), .IN2(n1154), .S(n7999), .Q(n12113)
         );
  MUX21X1 U14457 ( .IN1(\mem2[212][20] ), .IN2(n1132), .S(n7999), .Q(n12112)
         );
  MUX21X1 U14458 ( .IN1(\mem2[212][19] ), .IN2(n1110), .S(n7999), .Q(n12111)
         );
  MUX21X1 U14459 ( .IN1(\mem2[212][18] ), .IN2(n1088), .S(n7999), .Q(n12110)
         );
  MUX21X1 U14460 ( .IN1(\mem2[212][17] ), .IN2(n1066), .S(n7999), .Q(n12109)
         );
  MUX21X1 U14461 ( .IN1(\mem2[212][16] ), .IN2(n1044), .S(n7999), .Q(n12108)
         );
  AND2X1 U14462 ( .IN1(n7988), .IN2(n7122), .Q(n7999) );
  MUX21X1 U14463 ( .IN1(\mem2[211][23] ), .IN2(n1198), .S(n8000), .Q(n12107)
         );
  MUX21X1 U14464 ( .IN1(\mem2[211][22] ), .IN2(n1176), .S(n8000), .Q(n12106)
         );
  MUX21X1 U14465 ( .IN1(\mem2[211][21] ), .IN2(n1154), .S(n8000), .Q(n12105)
         );
  MUX21X1 U14466 ( .IN1(\mem2[211][20] ), .IN2(n1132), .S(n8000), .Q(n12104)
         );
  MUX21X1 U14467 ( .IN1(\mem2[211][19] ), .IN2(n1110), .S(n8000), .Q(n12103)
         );
  MUX21X1 U14468 ( .IN1(\mem2[211][18] ), .IN2(n1088), .S(n8000), .Q(n12102)
         );
  MUX21X1 U14469 ( .IN1(\mem2[211][17] ), .IN2(n1066), .S(n8000), .Q(n12101)
         );
  MUX21X1 U14470 ( .IN1(\mem2[211][16] ), .IN2(n1044), .S(n8000), .Q(n12100)
         );
  AND2X1 U14471 ( .IN1(n7988), .IN2(n7124), .Q(n8000) );
  MUX21X1 U14472 ( .IN1(\mem2[210][23] ), .IN2(n1198), .S(n8001), .Q(n12099)
         );
  MUX21X1 U14473 ( .IN1(\mem2[210][22] ), .IN2(n1176), .S(n8001), .Q(n12098)
         );
  MUX21X1 U14474 ( .IN1(\mem2[210][21] ), .IN2(n1154), .S(n8001), .Q(n12097)
         );
  MUX21X1 U14475 ( .IN1(\mem2[210][20] ), .IN2(n1132), .S(n8001), .Q(n12096)
         );
  MUX21X1 U14476 ( .IN1(\mem2[210][19] ), .IN2(n1110), .S(n8001), .Q(n12095)
         );
  MUX21X1 U14477 ( .IN1(\mem2[210][18] ), .IN2(n1088), .S(n8001), .Q(n12094)
         );
  MUX21X1 U14478 ( .IN1(\mem2[210][17] ), .IN2(n1066), .S(n8001), .Q(n12093)
         );
  MUX21X1 U14479 ( .IN1(\mem2[210][16] ), .IN2(n1044), .S(n8001), .Q(n12092)
         );
  AND2X1 U14480 ( .IN1(n7988), .IN2(n7126), .Q(n8001) );
  MUX21X1 U14481 ( .IN1(\mem2[209][23] ), .IN2(n1198), .S(n8002), .Q(n12091)
         );
  MUX21X1 U14482 ( .IN1(\mem2[209][22] ), .IN2(n1176), .S(n8002), .Q(n12090)
         );
  MUX21X1 U14483 ( .IN1(\mem2[209][21] ), .IN2(n1154), .S(n8002), .Q(n12089)
         );
  MUX21X1 U14484 ( .IN1(\mem2[209][20] ), .IN2(n1132), .S(n8002), .Q(n12088)
         );
  MUX21X1 U14485 ( .IN1(\mem2[209][19] ), .IN2(n1110), .S(n8002), .Q(n12087)
         );
  MUX21X1 U14486 ( .IN1(\mem2[209][18] ), .IN2(n1088), .S(n8002), .Q(n12086)
         );
  MUX21X1 U14487 ( .IN1(\mem2[209][17] ), .IN2(n1066), .S(n8002), .Q(n12085)
         );
  MUX21X1 U14488 ( .IN1(\mem2[209][16] ), .IN2(n1044), .S(n8002), .Q(n12084)
         );
  AND2X1 U14489 ( .IN1(n7988), .IN2(n7128), .Q(n8002) );
  MUX21X1 U14490 ( .IN1(\mem2[208][23] ), .IN2(n1198), .S(n8003), .Q(n12083)
         );
  MUX21X1 U14491 ( .IN1(\mem2[208][22] ), .IN2(n1176), .S(n8003), .Q(n12082)
         );
  MUX21X1 U14492 ( .IN1(\mem2[208][21] ), .IN2(n1154), .S(n8003), .Q(n12081)
         );
  MUX21X1 U14493 ( .IN1(\mem2[208][20] ), .IN2(n1132), .S(n8003), .Q(n12080)
         );
  MUX21X1 U14494 ( .IN1(\mem2[208][19] ), .IN2(n1110), .S(n8003), .Q(n12079)
         );
  MUX21X1 U14495 ( .IN1(\mem2[208][18] ), .IN2(n1088), .S(n8003), .Q(n12078)
         );
  MUX21X1 U14496 ( .IN1(\mem2[208][17] ), .IN2(n1066), .S(n8003), .Q(n12077)
         );
  MUX21X1 U14497 ( .IN1(\mem2[208][16] ), .IN2(n1044), .S(n8003), .Q(n12076)
         );
  AND2X1 U14498 ( .IN1(n7988), .IN2(n7130), .Q(n8003) );
  AND2X1 U14499 ( .IN1(n7966), .IN2(n7168), .Q(n7988) );
  AND2X1 U14500 ( .IN1(n8004), .IN2(n7967), .Q(n7168) );
  MUX21X1 U14501 ( .IN1(\mem2[207][23] ), .IN2(n1199), .S(n8005), .Q(n12075)
         );
  MUX21X1 U14502 ( .IN1(\mem2[207][22] ), .IN2(n1177), .S(n8005), .Q(n12074)
         );
  MUX21X1 U14503 ( .IN1(\mem2[207][21] ), .IN2(n1155), .S(n8005), .Q(n12073)
         );
  MUX21X1 U14504 ( .IN1(\mem2[207][20] ), .IN2(n1133), .S(n8005), .Q(n12072)
         );
  MUX21X1 U14505 ( .IN1(\mem2[207][19] ), .IN2(n1111), .S(n8005), .Q(n12071)
         );
  MUX21X1 U14506 ( .IN1(\mem2[207][18] ), .IN2(n1089), .S(n8005), .Q(n12070)
         );
  MUX21X1 U14507 ( .IN1(\mem2[207][17] ), .IN2(n1067), .S(n8005), .Q(n12069)
         );
  MUX21X1 U14508 ( .IN1(\mem2[207][16] ), .IN2(n1045), .S(n8005), .Q(n12068)
         );
  AND2X1 U14509 ( .IN1(n8006), .IN2(n7099), .Q(n8005) );
  MUX21X1 U14510 ( .IN1(\mem2[206][23] ), .IN2(n1199), .S(n8007), .Q(n12067)
         );
  MUX21X1 U14511 ( .IN1(\mem2[206][22] ), .IN2(n1177), .S(n8007), .Q(n12066)
         );
  MUX21X1 U14512 ( .IN1(\mem2[206][21] ), .IN2(n1155), .S(n8007), .Q(n12065)
         );
  MUX21X1 U14513 ( .IN1(\mem2[206][20] ), .IN2(n1133), .S(n8007), .Q(n12064)
         );
  MUX21X1 U14514 ( .IN1(\mem2[206][19] ), .IN2(n1111), .S(n8007), .Q(n12063)
         );
  MUX21X1 U14515 ( .IN1(\mem2[206][18] ), .IN2(n1089), .S(n8007), .Q(n12062)
         );
  MUX21X1 U14516 ( .IN1(\mem2[206][17] ), .IN2(n1067), .S(n8007), .Q(n12061)
         );
  MUX21X1 U14517 ( .IN1(\mem2[206][16] ), .IN2(n1045), .S(n8007), .Q(n12060)
         );
  AND2X1 U14518 ( .IN1(n8006), .IN2(n7102), .Q(n8007) );
  MUX21X1 U14519 ( .IN1(\mem2[205][23] ), .IN2(n1199), .S(n8008), .Q(n12059)
         );
  MUX21X1 U14520 ( .IN1(\mem2[205][22] ), .IN2(n1177), .S(n8008), .Q(n12058)
         );
  MUX21X1 U14521 ( .IN1(\mem2[205][21] ), .IN2(n1155), .S(n8008), .Q(n12057)
         );
  MUX21X1 U14522 ( .IN1(\mem2[205][20] ), .IN2(n1133), .S(n8008), .Q(n12056)
         );
  MUX21X1 U14523 ( .IN1(\mem2[205][19] ), .IN2(n1111), .S(n8008), .Q(n12055)
         );
  MUX21X1 U14524 ( .IN1(\mem2[205][18] ), .IN2(n1089), .S(n8008), .Q(n12054)
         );
  MUX21X1 U14525 ( .IN1(\mem2[205][17] ), .IN2(n1067), .S(n8008), .Q(n12053)
         );
  MUX21X1 U14526 ( .IN1(\mem2[205][16] ), .IN2(n1045), .S(n8008), .Q(n12052)
         );
  AND2X1 U14527 ( .IN1(n8006), .IN2(n7104), .Q(n8008) );
  MUX21X1 U14528 ( .IN1(\mem2[204][23] ), .IN2(n1199), .S(n8009), .Q(n12051)
         );
  MUX21X1 U14529 ( .IN1(\mem2[204][22] ), .IN2(n1177), .S(n8009), .Q(n12050)
         );
  MUX21X1 U14530 ( .IN1(\mem2[204][21] ), .IN2(n1155), .S(n8009), .Q(n12049)
         );
  MUX21X1 U14531 ( .IN1(\mem2[204][20] ), .IN2(n1133), .S(n8009), .Q(n12048)
         );
  MUX21X1 U14532 ( .IN1(\mem2[204][19] ), .IN2(n1111), .S(n8009), .Q(n12047)
         );
  MUX21X1 U14533 ( .IN1(\mem2[204][18] ), .IN2(n1089), .S(n8009), .Q(n12046)
         );
  MUX21X1 U14534 ( .IN1(\mem2[204][17] ), .IN2(n1067), .S(n8009), .Q(n12045)
         );
  MUX21X1 U14535 ( .IN1(\mem2[204][16] ), .IN2(n1045), .S(n8009), .Q(n12044)
         );
  AND2X1 U14536 ( .IN1(n8006), .IN2(n7106), .Q(n8009) );
  MUX21X1 U14537 ( .IN1(\mem2[203][23] ), .IN2(n1199), .S(n8010), .Q(n12043)
         );
  MUX21X1 U14538 ( .IN1(\mem2[203][22] ), .IN2(n1177), .S(n8010), .Q(n12042)
         );
  MUX21X1 U14539 ( .IN1(\mem2[203][21] ), .IN2(n1155), .S(n8010), .Q(n12041)
         );
  MUX21X1 U14540 ( .IN1(\mem2[203][20] ), .IN2(n1133), .S(n8010), .Q(n12040)
         );
  MUX21X1 U14541 ( .IN1(\mem2[203][19] ), .IN2(n1111), .S(n8010), .Q(n12039)
         );
  MUX21X1 U14542 ( .IN1(\mem2[203][18] ), .IN2(n1089), .S(n8010), .Q(n12038)
         );
  MUX21X1 U14543 ( .IN1(\mem2[203][17] ), .IN2(n1067), .S(n8010), .Q(n12037)
         );
  MUX21X1 U14544 ( .IN1(\mem2[203][16] ), .IN2(n1045), .S(n8010), .Q(n12036)
         );
  AND2X1 U14545 ( .IN1(n8006), .IN2(n7108), .Q(n8010) );
  MUX21X1 U14546 ( .IN1(\mem2[202][23] ), .IN2(n1199), .S(n8011), .Q(n12035)
         );
  MUX21X1 U14547 ( .IN1(\mem2[202][22] ), .IN2(n1177), .S(n8011), .Q(n12034)
         );
  MUX21X1 U14548 ( .IN1(\mem2[202][21] ), .IN2(n1155), .S(n8011), .Q(n12033)
         );
  MUX21X1 U14549 ( .IN1(\mem2[202][20] ), .IN2(n1133), .S(n8011), .Q(n12032)
         );
  MUX21X1 U14550 ( .IN1(\mem2[202][19] ), .IN2(n1111), .S(n8011), .Q(n12031)
         );
  MUX21X1 U14551 ( .IN1(\mem2[202][18] ), .IN2(n1089), .S(n8011), .Q(n12030)
         );
  MUX21X1 U14552 ( .IN1(\mem2[202][17] ), .IN2(n1067), .S(n8011), .Q(n12029)
         );
  MUX21X1 U14553 ( .IN1(\mem2[202][16] ), .IN2(n1045), .S(n8011), .Q(n12028)
         );
  AND2X1 U14554 ( .IN1(n8006), .IN2(n7110), .Q(n8011) );
  MUX21X1 U14555 ( .IN1(\mem2[201][23] ), .IN2(n1199), .S(n8012), .Q(n12027)
         );
  MUX21X1 U14556 ( .IN1(\mem2[201][22] ), .IN2(n1177), .S(n8012), .Q(n12026)
         );
  MUX21X1 U14557 ( .IN1(\mem2[201][21] ), .IN2(n1155), .S(n8012), .Q(n12025)
         );
  MUX21X1 U14558 ( .IN1(\mem2[201][20] ), .IN2(n1133), .S(n8012), .Q(n12024)
         );
  MUX21X1 U14559 ( .IN1(\mem2[201][19] ), .IN2(n1111), .S(n8012), .Q(n12023)
         );
  MUX21X1 U14560 ( .IN1(\mem2[201][18] ), .IN2(n1089), .S(n8012), .Q(n12022)
         );
  MUX21X1 U14561 ( .IN1(\mem2[201][17] ), .IN2(n1067), .S(n8012), .Q(n12021)
         );
  MUX21X1 U14562 ( .IN1(\mem2[201][16] ), .IN2(n1045), .S(n8012), .Q(n12020)
         );
  AND2X1 U14563 ( .IN1(n8006), .IN2(n7112), .Q(n8012) );
  MUX21X1 U14564 ( .IN1(\mem2[200][23] ), .IN2(n1199), .S(n8013), .Q(n12019)
         );
  MUX21X1 U14565 ( .IN1(\mem2[200][22] ), .IN2(n1177), .S(n8013), .Q(n12018)
         );
  MUX21X1 U14566 ( .IN1(\mem2[200][21] ), .IN2(n1155), .S(n8013), .Q(n12017)
         );
  MUX21X1 U14567 ( .IN1(\mem2[200][20] ), .IN2(n1133), .S(n8013), .Q(n12016)
         );
  MUX21X1 U14568 ( .IN1(\mem2[200][19] ), .IN2(n1111), .S(n8013), .Q(n12015)
         );
  MUX21X1 U14569 ( .IN1(\mem2[200][18] ), .IN2(n1089), .S(n8013), .Q(n12014)
         );
  MUX21X1 U14570 ( .IN1(\mem2[200][17] ), .IN2(n1067), .S(n8013), .Q(n12013)
         );
  MUX21X1 U14571 ( .IN1(\mem2[200][16] ), .IN2(n1045), .S(n8013), .Q(n12012)
         );
  AND2X1 U14572 ( .IN1(n8006), .IN2(n7114), .Q(n8013) );
  MUX21X1 U14573 ( .IN1(\mem2[199][23] ), .IN2(n1199), .S(n8014), .Q(n12011)
         );
  MUX21X1 U14574 ( .IN1(\mem2[199][22] ), .IN2(n1177), .S(n8014), .Q(n12010)
         );
  MUX21X1 U14575 ( .IN1(\mem2[199][21] ), .IN2(n1155), .S(n8014), .Q(n12009)
         );
  MUX21X1 U14576 ( .IN1(\mem2[199][20] ), .IN2(n1133), .S(n8014), .Q(n12008)
         );
  MUX21X1 U14577 ( .IN1(\mem2[199][19] ), .IN2(n1111), .S(n8014), .Q(n12007)
         );
  MUX21X1 U14578 ( .IN1(\mem2[199][18] ), .IN2(n1089), .S(n8014), .Q(n12006)
         );
  MUX21X1 U14579 ( .IN1(\mem2[199][17] ), .IN2(n1067), .S(n8014), .Q(n12005)
         );
  MUX21X1 U14580 ( .IN1(\mem2[199][16] ), .IN2(n1045), .S(n8014), .Q(n12004)
         );
  AND2X1 U14581 ( .IN1(n8006), .IN2(n7116), .Q(n8014) );
  MUX21X1 U14582 ( .IN1(\mem2[198][23] ), .IN2(n1199), .S(n8015), .Q(n12003)
         );
  MUX21X1 U14583 ( .IN1(\mem2[198][22] ), .IN2(n1177), .S(n8015), .Q(n12002)
         );
  MUX21X1 U14584 ( .IN1(\mem2[198][21] ), .IN2(n1155), .S(n8015), .Q(n12001)
         );
  MUX21X1 U14585 ( .IN1(\mem2[198][20] ), .IN2(n1133), .S(n8015), .Q(n12000)
         );
  MUX21X1 U14586 ( .IN1(\mem2[198][19] ), .IN2(n1111), .S(n8015), .Q(n11999)
         );
  MUX21X1 U14587 ( .IN1(\mem2[198][18] ), .IN2(n1089), .S(n8015), .Q(n11998)
         );
  MUX21X1 U14588 ( .IN1(\mem2[198][17] ), .IN2(n1067), .S(n8015), .Q(n11997)
         );
  MUX21X1 U14589 ( .IN1(\mem2[198][16] ), .IN2(n1045), .S(n8015), .Q(n11996)
         );
  AND2X1 U14590 ( .IN1(n8006), .IN2(n7118), .Q(n8015) );
  MUX21X1 U14591 ( .IN1(\mem2[197][23] ), .IN2(n1199), .S(n8016), .Q(n11995)
         );
  MUX21X1 U14592 ( .IN1(\mem2[197][22] ), .IN2(n1177), .S(n8016), .Q(n11994)
         );
  MUX21X1 U14593 ( .IN1(\mem2[197][21] ), .IN2(n1155), .S(n8016), .Q(n11993)
         );
  MUX21X1 U14594 ( .IN1(\mem2[197][20] ), .IN2(n1133), .S(n8016), .Q(n11992)
         );
  MUX21X1 U14595 ( .IN1(\mem2[197][19] ), .IN2(n1111), .S(n8016), .Q(n11991)
         );
  MUX21X1 U14596 ( .IN1(\mem2[197][18] ), .IN2(n1089), .S(n8016), .Q(n11990)
         );
  MUX21X1 U14597 ( .IN1(\mem2[197][17] ), .IN2(n1067), .S(n8016), .Q(n11989)
         );
  MUX21X1 U14598 ( .IN1(\mem2[197][16] ), .IN2(n1045), .S(n8016), .Q(n11988)
         );
  AND2X1 U14599 ( .IN1(n8006), .IN2(n7120), .Q(n8016) );
  MUX21X1 U14600 ( .IN1(\mem2[196][23] ), .IN2(n1199), .S(n8017), .Q(n11987)
         );
  MUX21X1 U14601 ( .IN1(\mem2[196][22] ), .IN2(n1177), .S(n8017), .Q(n11986)
         );
  MUX21X1 U14602 ( .IN1(\mem2[196][21] ), .IN2(n1155), .S(n8017), .Q(n11985)
         );
  MUX21X1 U14603 ( .IN1(\mem2[196][20] ), .IN2(n1133), .S(n8017), .Q(n11984)
         );
  MUX21X1 U14604 ( .IN1(\mem2[196][19] ), .IN2(n1111), .S(n8017), .Q(n11983)
         );
  MUX21X1 U14605 ( .IN1(\mem2[196][18] ), .IN2(n1089), .S(n8017), .Q(n11982)
         );
  MUX21X1 U14606 ( .IN1(\mem2[196][17] ), .IN2(n1067), .S(n8017), .Q(n11981)
         );
  MUX21X1 U14607 ( .IN1(\mem2[196][16] ), .IN2(n1045), .S(n8017), .Q(n11980)
         );
  AND2X1 U14608 ( .IN1(n8006), .IN2(n7122), .Q(n8017) );
  MUX21X1 U14609 ( .IN1(\mem2[195][23] ), .IN2(n1200), .S(n8018), .Q(n11979)
         );
  MUX21X1 U14610 ( .IN1(\mem2[195][22] ), .IN2(n1178), .S(n8018), .Q(n11978)
         );
  MUX21X1 U14611 ( .IN1(\mem2[195][21] ), .IN2(n1156), .S(n8018), .Q(n11977)
         );
  MUX21X1 U14612 ( .IN1(\mem2[195][20] ), .IN2(n1134), .S(n8018), .Q(n11976)
         );
  MUX21X1 U14613 ( .IN1(\mem2[195][19] ), .IN2(n1112), .S(n8018), .Q(n11975)
         );
  MUX21X1 U14614 ( .IN1(\mem2[195][18] ), .IN2(n1090), .S(n8018), .Q(n11974)
         );
  MUX21X1 U14615 ( .IN1(\mem2[195][17] ), .IN2(n1068), .S(n8018), .Q(n11973)
         );
  MUX21X1 U14616 ( .IN1(\mem2[195][16] ), .IN2(n1046), .S(n8018), .Q(n11972)
         );
  AND2X1 U14617 ( .IN1(n8006), .IN2(n7124), .Q(n8018) );
  MUX21X1 U14618 ( .IN1(\mem2[194][23] ), .IN2(n1200), .S(n8019), .Q(n11971)
         );
  MUX21X1 U14619 ( .IN1(\mem2[194][22] ), .IN2(n1178), .S(n8019), .Q(n11970)
         );
  MUX21X1 U14620 ( .IN1(\mem2[194][21] ), .IN2(n1156), .S(n8019), .Q(n11969)
         );
  MUX21X1 U14621 ( .IN1(\mem2[194][20] ), .IN2(n1134), .S(n8019), .Q(n11968)
         );
  MUX21X1 U14622 ( .IN1(\mem2[194][19] ), .IN2(n1112), .S(n8019), .Q(n11967)
         );
  MUX21X1 U14623 ( .IN1(\mem2[194][18] ), .IN2(n1090), .S(n8019), .Q(n11966)
         );
  MUX21X1 U14624 ( .IN1(\mem2[194][17] ), .IN2(n1068), .S(n8019), .Q(n11965)
         );
  MUX21X1 U14625 ( .IN1(\mem2[194][16] ), .IN2(n1046), .S(n8019), .Q(n11964)
         );
  AND2X1 U14626 ( .IN1(n8006), .IN2(n7126), .Q(n8019) );
  MUX21X1 U14627 ( .IN1(\mem2[193][23] ), .IN2(n1200), .S(n8020), .Q(n11963)
         );
  MUX21X1 U14628 ( .IN1(\mem2[193][22] ), .IN2(n1178), .S(n8020), .Q(n11962)
         );
  MUX21X1 U14629 ( .IN1(\mem2[193][21] ), .IN2(n1156), .S(n8020), .Q(n11961)
         );
  MUX21X1 U14630 ( .IN1(\mem2[193][20] ), .IN2(n1134), .S(n8020), .Q(n11960)
         );
  MUX21X1 U14631 ( .IN1(\mem2[193][19] ), .IN2(n1112), .S(n8020), .Q(n11959)
         );
  MUX21X1 U14632 ( .IN1(\mem2[193][18] ), .IN2(n1090), .S(n8020), .Q(n11958)
         );
  MUX21X1 U14633 ( .IN1(\mem2[193][17] ), .IN2(n1068), .S(n8020), .Q(n11957)
         );
  MUX21X1 U14634 ( .IN1(\mem2[193][16] ), .IN2(n1046), .S(n8020), .Q(n11956)
         );
  AND2X1 U14635 ( .IN1(n8006), .IN2(n7128), .Q(n8020) );
  MUX21X1 U14636 ( .IN1(\mem2[192][23] ), .IN2(n1200), .S(n8021), .Q(n11955)
         );
  MUX21X1 U14637 ( .IN1(\mem2[192][22] ), .IN2(n1178), .S(n8021), .Q(n11954)
         );
  MUX21X1 U14638 ( .IN1(\mem2[192][21] ), .IN2(n1156), .S(n8021), .Q(n11953)
         );
  MUX21X1 U14639 ( .IN1(\mem2[192][20] ), .IN2(n1134), .S(n8021), .Q(n11952)
         );
  MUX21X1 U14640 ( .IN1(\mem2[192][19] ), .IN2(n1112), .S(n8021), .Q(n11951)
         );
  MUX21X1 U14641 ( .IN1(\mem2[192][18] ), .IN2(n1090), .S(n8021), .Q(n11950)
         );
  MUX21X1 U14642 ( .IN1(\mem2[192][17] ), .IN2(n1068), .S(n8021), .Q(n11949)
         );
  MUX21X1 U14643 ( .IN1(\mem2[192][16] ), .IN2(n1046), .S(n8021), .Q(n11948)
         );
  AND2X1 U14644 ( .IN1(n8006), .IN2(n7130), .Q(n8021) );
  AND2X1 U14645 ( .IN1(n7966), .IN2(n7186), .Q(n8006) );
  AND2X1 U14646 ( .IN1(n8022), .IN2(n7967), .Q(n7186) );
  NOR2X0 U14647 ( .IN1(n8023), .IN2(n8024), .QN(n7967) );
  MUX21X1 U14648 ( .IN1(\mem2[191][23] ), .IN2(n1200), .S(n8025), .Q(n11947)
         );
  MUX21X1 U14649 ( .IN1(\mem2[191][22] ), .IN2(n1178), .S(n8025), .Q(n11946)
         );
  MUX21X1 U14650 ( .IN1(\mem2[191][21] ), .IN2(n1156), .S(n8025), .Q(n11945)
         );
  MUX21X1 U14651 ( .IN1(\mem2[191][20] ), .IN2(n1134), .S(n8025), .Q(n11944)
         );
  MUX21X1 U14652 ( .IN1(\mem2[191][19] ), .IN2(n1112), .S(n8025), .Q(n11943)
         );
  MUX21X1 U14653 ( .IN1(\mem2[191][18] ), .IN2(n1090), .S(n8025), .Q(n11942)
         );
  MUX21X1 U14654 ( .IN1(\mem2[191][17] ), .IN2(n1068), .S(n8025), .Q(n11941)
         );
  MUX21X1 U14655 ( .IN1(\mem2[191][16] ), .IN2(n1046), .S(n8025), .Q(n11940)
         );
  AND2X1 U14656 ( .IN1(n8026), .IN2(n7099), .Q(n8025) );
  MUX21X1 U14657 ( .IN1(\mem2[190][23] ), .IN2(n1200), .S(n8027), .Q(n11939)
         );
  MUX21X1 U14658 ( .IN1(\mem2[190][22] ), .IN2(n1178), .S(n8027), .Q(n11938)
         );
  MUX21X1 U14659 ( .IN1(\mem2[190][21] ), .IN2(n1156), .S(n8027), .Q(n11937)
         );
  MUX21X1 U14660 ( .IN1(\mem2[190][20] ), .IN2(n1134), .S(n8027), .Q(n11936)
         );
  MUX21X1 U14661 ( .IN1(\mem2[190][19] ), .IN2(n1112), .S(n8027), .Q(n11935)
         );
  MUX21X1 U14662 ( .IN1(\mem2[190][18] ), .IN2(n1090), .S(n8027), .Q(n11934)
         );
  MUX21X1 U14663 ( .IN1(\mem2[190][17] ), .IN2(n1068), .S(n8027), .Q(n11933)
         );
  MUX21X1 U14664 ( .IN1(\mem2[190][16] ), .IN2(n1046), .S(n8027), .Q(n11932)
         );
  AND2X1 U14665 ( .IN1(n8026), .IN2(n7102), .Q(n8027) );
  MUX21X1 U14666 ( .IN1(\mem2[189][23] ), .IN2(n1200), .S(n8028), .Q(n11931)
         );
  MUX21X1 U14667 ( .IN1(\mem2[189][22] ), .IN2(n1178), .S(n8028), .Q(n11930)
         );
  MUX21X1 U14668 ( .IN1(\mem2[189][21] ), .IN2(n1156), .S(n8028), .Q(n11929)
         );
  MUX21X1 U14669 ( .IN1(\mem2[189][20] ), .IN2(n1134), .S(n8028), .Q(n11928)
         );
  MUX21X1 U14670 ( .IN1(\mem2[189][19] ), .IN2(n1112), .S(n8028), .Q(n11927)
         );
  MUX21X1 U14671 ( .IN1(\mem2[189][18] ), .IN2(n1090), .S(n8028), .Q(n11926)
         );
  MUX21X1 U14672 ( .IN1(\mem2[189][17] ), .IN2(n1068), .S(n8028), .Q(n11925)
         );
  MUX21X1 U14673 ( .IN1(\mem2[189][16] ), .IN2(n1046), .S(n8028), .Q(n11924)
         );
  AND2X1 U14674 ( .IN1(n8026), .IN2(n7104), .Q(n8028) );
  MUX21X1 U14675 ( .IN1(\mem2[188][23] ), .IN2(n1200), .S(n8029), .Q(n11923)
         );
  MUX21X1 U14676 ( .IN1(\mem2[188][22] ), .IN2(n1178), .S(n8029), .Q(n11922)
         );
  MUX21X1 U14677 ( .IN1(\mem2[188][21] ), .IN2(n1156), .S(n8029), .Q(n11921)
         );
  MUX21X1 U14678 ( .IN1(\mem2[188][20] ), .IN2(n1134), .S(n8029), .Q(n11920)
         );
  MUX21X1 U14679 ( .IN1(\mem2[188][19] ), .IN2(n1112), .S(n8029), .Q(n11919)
         );
  MUX21X1 U14680 ( .IN1(\mem2[188][18] ), .IN2(n1090), .S(n8029), .Q(n11918)
         );
  MUX21X1 U14681 ( .IN1(\mem2[188][17] ), .IN2(n1068), .S(n8029), .Q(n11917)
         );
  MUX21X1 U14682 ( .IN1(\mem2[188][16] ), .IN2(n1046), .S(n8029), .Q(n11916)
         );
  AND2X1 U14683 ( .IN1(n8026), .IN2(n7106), .Q(n8029) );
  MUX21X1 U14684 ( .IN1(\mem2[187][23] ), .IN2(n1200), .S(n8030), .Q(n11915)
         );
  MUX21X1 U14685 ( .IN1(\mem2[187][22] ), .IN2(n1178), .S(n8030), .Q(n11914)
         );
  MUX21X1 U14686 ( .IN1(\mem2[187][21] ), .IN2(n1156), .S(n8030), .Q(n11913)
         );
  MUX21X1 U14687 ( .IN1(\mem2[187][20] ), .IN2(n1134), .S(n8030), .Q(n11912)
         );
  MUX21X1 U14688 ( .IN1(\mem2[187][19] ), .IN2(n1112), .S(n8030), .Q(n11911)
         );
  MUX21X1 U14689 ( .IN1(\mem2[187][18] ), .IN2(n1090), .S(n8030), .Q(n11910)
         );
  MUX21X1 U14690 ( .IN1(\mem2[187][17] ), .IN2(n1068), .S(n8030), .Q(n11909)
         );
  MUX21X1 U14691 ( .IN1(\mem2[187][16] ), .IN2(n1046), .S(n8030), .Q(n11908)
         );
  AND2X1 U14692 ( .IN1(n8026), .IN2(n7108), .Q(n8030) );
  MUX21X1 U14693 ( .IN1(\mem2[186][23] ), .IN2(n1200), .S(n8031), .Q(n11907)
         );
  MUX21X1 U14694 ( .IN1(\mem2[186][22] ), .IN2(n1178), .S(n8031), .Q(n11906)
         );
  MUX21X1 U14695 ( .IN1(\mem2[186][21] ), .IN2(n1156), .S(n8031), .Q(n11905)
         );
  MUX21X1 U14696 ( .IN1(\mem2[186][20] ), .IN2(n1134), .S(n8031), .Q(n11904)
         );
  MUX21X1 U14697 ( .IN1(\mem2[186][19] ), .IN2(n1112), .S(n8031), .Q(n11903)
         );
  MUX21X1 U14698 ( .IN1(\mem2[186][18] ), .IN2(n1090), .S(n8031), .Q(n11902)
         );
  MUX21X1 U14699 ( .IN1(\mem2[186][17] ), .IN2(n1068), .S(n8031), .Q(n11901)
         );
  MUX21X1 U14700 ( .IN1(\mem2[186][16] ), .IN2(n1046), .S(n8031), .Q(n11900)
         );
  AND2X1 U14701 ( .IN1(n8026), .IN2(n7110), .Q(n8031) );
  MUX21X1 U14702 ( .IN1(\mem2[185][23] ), .IN2(n1200), .S(n8032), .Q(n11899)
         );
  MUX21X1 U14703 ( .IN1(\mem2[185][22] ), .IN2(n1178), .S(n8032), .Q(n11898)
         );
  MUX21X1 U14704 ( .IN1(\mem2[185][21] ), .IN2(n1156), .S(n8032), .Q(n11897)
         );
  MUX21X1 U14705 ( .IN1(\mem2[185][20] ), .IN2(n1134), .S(n8032), .Q(n11896)
         );
  MUX21X1 U14706 ( .IN1(\mem2[185][19] ), .IN2(n1112), .S(n8032), .Q(n11895)
         );
  MUX21X1 U14707 ( .IN1(\mem2[185][18] ), .IN2(n1090), .S(n8032), .Q(n11894)
         );
  MUX21X1 U14708 ( .IN1(\mem2[185][17] ), .IN2(n1068), .S(n8032), .Q(n11893)
         );
  MUX21X1 U14709 ( .IN1(\mem2[185][16] ), .IN2(n1046), .S(n8032), .Q(n11892)
         );
  AND2X1 U14710 ( .IN1(n8026), .IN2(n7112), .Q(n8032) );
  MUX21X1 U14711 ( .IN1(\mem2[184][23] ), .IN2(n1200), .S(n8033), .Q(n11891)
         );
  MUX21X1 U14712 ( .IN1(\mem2[184][22] ), .IN2(n1178), .S(n8033), .Q(n11890)
         );
  MUX21X1 U14713 ( .IN1(\mem2[184][21] ), .IN2(n1156), .S(n8033), .Q(n11889)
         );
  MUX21X1 U14714 ( .IN1(\mem2[184][20] ), .IN2(n1134), .S(n8033), .Q(n11888)
         );
  MUX21X1 U14715 ( .IN1(\mem2[184][19] ), .IN2(n1112), .S(n8033), .Q(n11887)
         );
  MUX21X1 U14716 ( .IN1(\mem2[184][18] ), .IN2(n1090), .S(n8033), .Q(n11886)
         );
  MUX21X1 U14717 ( .IN1(\mem2[184][17] ), .IN2(n1068), .S(n8033), .Q(n11885)
         );
  MUX21X1 U14718 ( .IN1(\mem2[184][16] ), .IN2(n1046), .S(n8033), .Q(n11884)
         );
  AND2X1 U14719 ( .IN1(n8026), .IN2(n7114), .Q(n8033) );
  MUX21X1 U14720 ( .IN1(\mem2[183][23] ), .IN2(n1201), .S(n8034), .Q(n11883)
         );
  MUX21X1 U14721 ( .IN1(\mem2[183][22] ), .IN2(n1179), .S(n8034), .Q(n11882)
         );
  MUX21X1 U14722 ( .IN1(\mem2[183][21] ), .IN2(n1157), .S(n8034), .Q(n11881)
         );
  MUX21X1 U14723 ( .IN1(\mem2[183][20] ), .IN2(n1135), .S(n8034), .Q(n11880)
         );
  MUX21X1 U14724 ( .IN1(\mem2[183][19] ), .IN2(n1113), .S(n8034), .Q(n11879)
         );
  MUX21X1 U14725 ( .IN1(\mem2[183][18] ), .IN2(n1091), .S(n8034), .Q(n11878)
         );
  MUX21X1 U14726 ( .IN1(\mem2[183][17] ), .IN2(n1069), .S(n8034), .Q(n11877)
         );
  MUX21X1 U14727 ( .IN1(\mem2[183][16] ), .IN2(n1047), .S(n8034), .Q(n11876)
         );
  AND2X1 U14728 ( .IN1(n8026), .IN2(n7116), .Q(n8034) );
  MUX21X1 U14729 ( .IN1(\mem2[182][23] ), .IN2(n1201), .S(n8035), .Q(n11875)
         );
  MUX21X1 U14730 ( .IN1(\mem2[182][22] ), .IN2(n1179), .S(n8035), .Q(n11874)
         );
  MUX21X1 U14731 ( .IN1(\mem2[182][21] ), .IN2(n1157), .S(n8035), .Q(n11873)
         );
  MUX21X1 U14732 ( .IN1(\mem2[182][20] ), .IN2(n1135), .S(n8035), .Q(n11872)
         );
  MUX21X1 U14733 ( .IN1(\mem2[182][19] ), .IN2(n1113), .S(n8035), .Q(n11871)
         );
  MUX21X1 U14734 ( .IN1(\mem2[182][18] ), .IN2(n1091), .S(n8035), .Q(n11870)
         );
  MUX21X1 U14735 ( .IN1(\mem2[182][17] ), .IN2(n1069), .S(n8035), .Q(n11869)
         );
  MUX21X1 U14736 ( .IN1(\mem2[182][16] ), .IN2(n1047), .S(n8035), .Q(n11868)
         );
  AND2X1 U14737 ( .IN1(n8026), .IN2(n7118), .Q(n8035) );
  MUX21X1 U14738 ( .IN1(\mem2[181][23] ), .IN2(n1201), .S(n8036), .Q(n11867)
         );
  MUX21X1 U14739 ( .IN1(\mem2[181][22] ), .IN2(n1179), .S(n8036), .Q(n11866)
         );
  MUX21X1 U14740 ( .IN1(\mem2[181][21] ), .IN2(n1157), .S(n8036), .Q(n11865)
         );
  MUX21X1 U14741 ( .IN1(\mem2[181][20] ), .IN2(n1135), .S(n8036), .Q(n11864)
         );
  MUX21X1 U14742 ( .IN1(\mem2[181][19] ), .IN2(n1113), .S(n8036), .Q(n11863)
         );
  MUX21X1 U14743 ( .IN1(\mem2[181][18] ), .IN2(n1091), .S(n8036), .Q(n11862)
         );
  MUX21X1 U14744 ( .IN1(\mem2[181][17] ), .IN2(n1069), .S(n8036), .Q(n11861)
         );
  MUX21X1 U14745 ( .IN1(\mem2[181][16] ), .IN2(n1047), .S(n8036), .Q(n11860)
         );
  AND2X1 U14746 ( .IN1(n8026), .IN2(n7120), .Q(n8036) );
  MUX21X1 U14747 ( .IN1(\mem2[180][23] ), .IN2(n1201), .S(n8037), .Q(n11859)
         );
  MUX21X1 U14748 ( .IN1(\mem2[180][22] ), .IN2(n1179), .S(n8037), .Q(n11858)
         );
  MUX21X1 U14749 ( .IN1(\mem2[180][21] ), .IN2(n1157), .S(n8037), .Q(n11857)
         );
  MUX21X1 U14750 ( .IN1(\mem2[180][20] ), .IN2(n1135), .S(n8037), .Q(n11856)
         );
  MUX21X1 U14751 ( .IN1(\mem2[180][19] ), .IN2(n1113), .S(n8037), .Q(n11855)
         );
  MUX21X1 U14752 ( .IN1(\mem2[180][18] ), .IN2(n1091), .S(n8037), .Q(n11854)
         );
  MUX21X1 U14753 ( .IN1(\mem2[180][17] ), .IN2(n1069), .S(n8037), .Q(n11853)
         );
  MUX21X1 U14754 ( .IN1(\mem2[180][16] ), .IN2(n1047), .S(n8037), .Q(n11852)
         );
  AND2X1 U14755 ( .IN1(n8026), .IN2(n7122), .Q(n8037) );
  MUX21X1 U14756 ( .IN1(\mem2[179][23] ), .IN2(n1201), .S(n8038), .Q(n11851)
         );
  MUX21X1 U14757 ( .IN1(\mem2[179][22] ), .IN2(n1179), .S(n8038), .Q(n11850)
         );
  MUX21X1 U14758 ( .IN1(\mem2[179][21] ), .IN2(n1157), .S(n8038), .Q(n11849)
         );
  MUX21X1 U14759 ( .IN1(\mem2[179][20] ), .IN2(n1135), .S(n8038), .Q(n11848)
         );
  MUX21X1 U14760 ( .IN1(\mem2[179][19] ), .IN2(n1113), .S(n8038), .Q(n11847)
         );
  MUX21X1 U14761 ( .IN1(\mem2[179][18] ), .IN2(n1091), .S(n8038), .Q(n11846)
         );
  MUX21X1 U14762 ( .IN1(\mem2[179][17] ), .IN2(n1069), .S(n8038), .Q(n11845)
         );
  MUX21X1 U14763 ( .IN1(\mem2[179][16] ), .IN2(n1047), .S(n8038), .Q(n11844)
         );
  AND2X1 U14764 ( .IN1(n8026), .IN2(n7124), .Q(n8038) );
  MUX21X1 U14765 ( .IN1(\mem2[178][23] ), .IN2(n1201), .S(n8039), .Q(n11843)
         );
  MUX21X1 U14766 ( .IN1(\mem2[178][22] ), .IN2(n1179), .S(n8039), .Q(n11842)
         );
  MUX21X1 U14767 ( .IN1(\mem2[178][21] ), .IN2(n1157), .S(n8039), .Q(n11841)
         );
  MUX21X1 U14768 ( .IN1(\mem2[178][20] ), .IN2(n1135), .S(n8039), .Q(n11840)
         );
  MUX21X1 U14769 ( .IN1(\mem2[178][19] ), .IN2(n1113), .S(n8039), .Q(n11839)
         );
  MUX21X1 U14770 ( .IN1(\mem2[178][18] ), .IN2(n1091), .S(n8039), .Q(n11838)
         );
  MUX21X1 U14771 ( .IN1(\mem2[178][17] ), .IN2(n1069), .S(n8039), .Q(n11837)
         );
  MUX21X1 U14772 ( .IN1(\mem2[178][16] ), .IN2(n1047), .S(n8039), .Q(n11836)
         );
  AND2X1 U14773 ( .IN1(n8026), .IN2(n7126), .Q(n8039) );
  MUX21X1 U14774 ( .IN1(\mem2[177][23] ), .IN2(n1201), .S(n8040), .Q(n11835)
         );
  MUX21X1 U14775 ( .IN1(\mem2[177][22] ), .IN2(n1179), .S(n8040), .Q(n11834)
         );
  MUX21X1 U14776 ( .IN1(\mem2[177][21] ), .IN2(n1157), .S(n8040), .Q(n11833)
         );
  MUX21X1 U14777 ( .IN1(\mem2[177][20] ), .IN2(n1135), .S(n8040), .Q(n11832)
         );
  MUX21X1 U14778 ( .IN1(\mem2[177][19] ), .IN2(n1113), .S(n8040), .Q(n11831)
         );
  MUX21X1 U14779 ( .IN1(\mem2[177][18] ), .IN2(n1091), .S(n8040), .Q(n11830)
         );
  MUX21X1 U14780 ( .IN1(\mem2[177][17] ), .IN2(n1069), .S(n8040), .Q(n11829)
         );
  MUX21X1 U14781 ( .IN1(\mem2[177][16] ), .IN2(n1047), .S(n8040), .Q(n11828)
         );
  AND2X1 U14782 ( .IN1(n8026), .IN2(n7128), .Q(n8040) );
  MUX21X1 U14783 ( .IN1(\mem2[176][23] ), .IN2(n1201), .S(n8041), .Q(n11827)
         );
  MUX21X1 U14784 ( .IN1(\mem2[176][22] ), .IN2(n1179), .S(n8041), .Q(n11826)
         );
  MUX21X1 U14785 ( .IN1(\mem2[176][21] ), .IN2(n1157), .S(n8041), .Q(n11825)
         );
  MUX21X1 U14786 ( .IN1(\mem2[176][20] ), .IN2(n1135), .S(n8041), .Q(n11824)
         );
  MUX21X1 U14787 ( .IN1(\mem2[176][19] ), .IN2(n1113), .S(n8041), .Q(n11823)
         );
  MUX21X1 U14788 ( .IN1(\mem2[176][18] ), .IN2(n1091), .S(n8041), .Q(n11822)
         );
  MUX21X1 U14789 ( .IN1(\mem2[176][17] ), .IN2(n1069), .S(n8041), .Q(n11821)
         );
  MUX21X1 U14790 ( .IN1(\mem2[176][16] ), .IN2(n1047), .S(n8041), .Q(n11820)
         );
  AND2X1 U14791 ( .IN1(n8026), .IN2(n7130), .Q(n8041) );
  AND2X1 U14792 ( .IN1(n7966), .IN2(n7204), .Q(n8026) );
  AND2X1 U14793 ( .IN1(n8042), .IN2(n7968), .Q(n7204) );
  MUX21X1 U14794 ( .IN1(\mem2[175][23] ), .IN2(n1201), .S(n8043), .Q(n11819)
         );
  MUX21X1 U14795 ( .IN1(\mem2[175][22] ), .IN2(n1179), .S(n8043), .Q(n11818)
         );
  MUX21X1 U14796 ( .IN1(\mem2[175][21] ), .IN2(n1157), .S(n8043), .Q(n11817)
         );
  MUX21X1 U14797 ( .IN1(\mem2[175][20] ), .IN2(n1135), .S(n8043), .Q(n11816)
         );
  MUX21X1 U14798 ( .IN1(\mem2[175][19] ), .IN2(n1113), .S(n8043), .Q(n11815)
         );
  MUX21X1 U14799 ( .IN1(\mem2[175][18] ), .IN2(n1091), .S(n8043), .Q(n11814)
         );
  MUX21X1 U14800 ( .IN1(\mem2[175][17] ), .IN2(n1069), .S(n8043), .Q(n11813)
         );
  MUX21X1 U14801 ( .IN1(\mem2[175][16] ), .IN2(n1047), .S(n8043), .Q(n11812)
         );
  AND2X1 U14802 ( .IN1(n8044), .IN2(n7099), .Q(n8043) );
  MUX21X1 U14803 ( .IN1(\mem2[174][23] ), .IN2(n1201), .S(n8045), .Q(n11811)
         );
  MUX21X1 U14804 ( .IN1(\mem2[174][22] ), .IN2(n1179), .S(n8045), .Q(n11810)
         );
  MUX21X1 U14805 ( .IN1(\mem2[174][21] ), .IN2(n1157), .S(n8045), .Q(n11809)
         );
  MUX21X1 U14806 ( .IN1(\mem2[174][20] ), .IN2(n1135), .S(n8045), .Q(n11808)
         );
  MUX21X1 U14807 ( .IN1(\mem2[174][19] ), .IN2(n1113), .S(n8045), .Q(n11807)
         );
  MUX21X1 U14808 ( .IN1(\mem2[174][18] ), .IN2(n1091), .S(n8045), .Q(n11806)
         );
  MUX21X1 U14809 ( .IN1(\mem2[174][17] ), .IN2(n1069), .S(n8045), .Q(n11805)
         );
  MUX21X1 U14810 ( .IN1(\mem2[174][16] ), .IN2(n1047), .S(n8045), .Q(n11804)
         );
  AND2X1 U14811 ( .IN1(n8044), .IN2(n7102), .Q(n8045) );
  MUX21X1 U14812 ( .IN1(\mem2[173][23] ), .IN2(n1201), .S(n8046), .Q(n11803)
         );
  MUX21X1 U14813 ( .IN1(\mem2[173][22] ), .IN2(n1179), .S(n8046), .Q(n11802)
         );
  MUX21X1 U14814 ( .IN1(\mem2[173][21] ), .IN2(n1157), .S(n8046), .Q(n11801)
         );
  MUX21X1 U14815 ( .IN1(\mem2[173][20] ), .IN2(n1135), .S(n8046), .Q(n11800)
         );
  MUX21X1 U14816 ( .IN1(\mem2[173][19] ), .IN2(n1113), .S(n8046), .Q(n11799)
         );
  MUX21X1 U14817 ( .IN1(\mem2[173][18] ), .IN2(n1091), .S(n8046), .Q(n11798)
         );
  MUX21X1 U14818 ( .IN1(\mem2[173][17] ), .IN2(n1069), .S(n8046), .Q(n11797)
         );
  MUX21X1 U14819 ( .IN1(\mem2[173][16] ), .IN2(n1047), .S(n8046), .Q(n11796)
         );
  AND2X1 U14820 ( .IN1(n8044), .IN2(n7104), .Q(n8046) );
  MUX21X1 U14821 ( .IN1(\mem2[172][23] ), .IN2(n1201), .S(n8047), .Q(n11795)
         );
  MUX21X1 U14822 ( .IN1(\mem2[172][22] ), .IN2(n1179), .S(n8047), .Q(n11794)
         );
  MUX21X1 U14823 ( .IN1(\mem2[172][21] ), .IN2(n1157), .S(n8047), .Q(n11793)
         );
  MUX21X1 U14824 ( .IN1(\mem2[172][20] ), .IN2(n1135), .S(n8047), .Q(n11792)
         );
  MUX21X1 U14825 ( .IN1(\mem2[172][19] ), .IN2(n1113), .S(n8047), .Q(n11791)
         );
  MUX21X1 U14826 ( .IN1(\mem2[172][18] ), .IN2(n1091), .S(n8047), .Q(n11790)
         );
  MUX21X1 U14827 ( .IN1(\mem2[172][17] ), .IN2(n1069), .S(n8047), .Q(n11789)
         );
  MUX21X1 U14828 ( .IN1(\mem2[172][16] ), .IN2(n1047), .S(n8047), .Q(n11788)
         );
  AND2X1 U14829 ( .IN1(n8044), .IN2(n7106), .Q(n8047) );
  MUX21X1 U14830 ( .IN1(\mem2[171][23] ), .IN2(n1202), .S(n8048), .Q(n11787)
         );
  MUX21X1 U14831 ( .IN1(\mem2[171][22] ), .IN2(n1180), .S(n8048), .Q(n11786)
         );
  MUX21X1 U14832 ( .IN1(\mem2[171][21] ), .IN2(n1158), .S(n8048), .Q(n11785)
         );
  MUX21X1 U14833 ( .IN1(\mem2[171][20] ), .IN2(n1136), .S(n8048), .Q(n11784)
         );
  MUX21X1 U14834 ( .IN1(\mem2[171][19] ), .IN2(n1114), .S(n8048), .Q(n11783)
         );
  MUX21X1 U14835 ( .IN1(\mem2[171][18] ), .IN2(n1092), .S(n8048), .Q(n11782)
         );
  MUX21X1 U14836 ( .IN1(\mem2[171][17] ), .IN2(n1070), .S(n8048), .Q(n11781)
         );
  MUX21X1 U14837 ( .IN1(\mem2[171][16] ), .IN2(n1048), .S(n8048), .Q(n11780)
         );
  AND2X1 U14838 ( .IN1(n8044), .IN2(n7108), .Q(n8048) );
  MUX21X1 U14839 ( .IN1(\mem2[170][23] ), .IN2(n1202), .S(n8049), .Q(n11779)
         );
  MUX21X1 U14840 ( .IN1(\mem2[170][22] ), .IN2(n1180), .S(n8049), .Q(n11778)
         );
  MUX21X1 U14841 ( .IN1(\mem2[170][21] ), .IN2(n1158), .S(n8049), .Q(n11777)
         );
  MUX21X1 U14842 ( .IN1(\mem2[170][20] ), .IN2(n1136), .S(n8049), .Q(n11776)
         );
  MUX21X1 U14843 ( .IN1(\mem2[170][19] ), .IN2(n1114), .S(n8049), .Q(n11775)
         );
  MUX21X1 U14844 ( .IN1(\mem2[170][18] ), .IN2(n1092), .S(n8049), .Q(n11774)
         );
  MUX21X1 U14845 ( .IN1(\mem2[170][17] ), .IN2(n1070), .S(n8049), .Q(n11773)
         );
  MUX21X1 U14846 ( .IN1(\mem2[170][16] ), .IN2(n1048), .S(n8049), .Q(n11772)
         );
  AND2X1 U14847 ( .IN1(n8044), .IN2(n7110), .Q(n8049) );
  MUX21X1 U14848 ( .IN1(\mem2[169][23] ), .IN2(n1202), .S(n8050), .Q(n11771)
         );
  MUX21X1 U14849 ( .IN1(\mem2[169][22] ), .IN2(n1180), .S(n8050), .Q(n11770)
         );
  MUX21X1 U14850 ( .IN1(\mem2[169][21] ), .IN2(n1158), .S(n8050), .Q(n11769)
         );
  MUX21X1 U14851 ( .IN1(\mem2[169][20] ), .IN2(n1136), .S(n8050), .Q(n11768)
         );
  MUX21X1 U14852 ( .IN1(\mem2[169][19] ), .IN2(n1114), .S(n8050), .Q(n11767)
         );
  MUX21X1 U14853 ( .IN1(\mem2[169][18] ), .IN2(n1092), .S(n8050), .Q(n11766)
         );
  MUX21X1 U14854 ( .IN1(\mem2[169][17] ), .IN2(n1070), .S(n8050), .Q(n11765)
         );
  MUX21X1 U14855 ( .IN1(\mem2[169][16] ), .IN2(n1048), .S(n8050), .Q(n11764)
         );
  AND2X1 U14856 ( .IN1(n8044), .IN2(n7112), .Q(n8050) );
  MUX21X1 U14857 ( .IN1(\mem2[168][23] ), .IN2(n1202), .S(n8051), .Q(n11763)
         );
  MUX21X1 U14858 ( .IN1(\mem2[168][22] ), .IN2(n1180), .S(n8051), .Q(n11762)
         );
  MUX21X1 U14859 ( .IN1(\mem2[168][21] ), .IN2(n1158), .S(n8051), .Q(n11761)
         );
  MUX21X1 U14860 ( .IN1(\mem2[168][20] ), .IN2(n1136), .S(n8051), .Q(n11760)
         );
  MUX21X1 U14861 ( .IN1(\mem2[168][19] ), .IN2(n1114), .S(n8051), .Q(n11759)
         );
  MUX21X1 U14862 ( .IN1(\mem2[168][18] ), .IN2(n1092), .S(n8051), .Q(n11758)
         );
  MUX21X1 U14863 ( .IN1(\mem2[168][17] ), .IN2(n1070), .S(n8051), .Q(n11757)
         );
  MUX21X1 U14864 ( .IN1(\mem2[168][16] ), .IN2(n1048), .S(n8051), .Q(n11756)
         );
  AND2X1 U14865 ( .IN1(n8044), .IN2(n7114), .Q(n8051) );
  MUX21X1 U14866 ( .IN1(\mem2[167][23] ), .IN2(n1202), .S(n8052), .Q(n11755)
         );
  MUX21X1 U14867 ( .IN1(\mem2[167][22] ), .IN2(n1180), .S(n8052), .Q(n11754)
         );
  MUX21X1 U14868 ( .IN1(\mem2[167][21] ), .IN2(n1158), .S(n8052), .Q(n11753)
         );
  MUX21X1 U14869 ( .IN1(\mem2[167][20] ), .IN2(n1136), .S(n8052), .Q(n11752)
         );
  MUX21X1 U14870 ( .IN1(\mem2[167][19] ), .IN2(n1114), .S(n8052), .Q(n11751)
         );
  MUX21X1 U14871 ( .IN1(\mem2[167][18] ), .IN2(n1092), .S(n8052), .Q(n11750)
         );
  MUX21X1 U14872 ( .IN1(\mem2[167][17] ), .IN2(n1070), .S(n8052), .Q(n11749)
         );
  MUX21X1 U14873 ( .IN1(\mem2[167][16] ), .IN2(n1048), .S(n8052), .Q(n11748)
         );
  AND2X1 U14874 ( .IN1(n8044), .IN2(n7116), .Q(n8052) );
  MUX21X1 U14875 ( .IN1(\mem2[166][23] ), .IN2(n1202), .S(n8053), .Q(n11747)
         );
  MUX21X1 U14876 ( .IN1(\mem2[166][22] ), .IN2(n1180), .S(n8053), .Q(n11746)
         );
  MUX21X1 U14877 ( .IN1(\mem2[166][21] ), .IN2(n1158), .S(n8053), .Q(n11745)
         );
  MUX21X1 U14878 ( .IN1(\mem2[166][20] ), .IN2(n1136), .S(n8053), .Q(n11744)
         );
  MUX21X1 U14879 ( .IN1(\mem2[166][19] ), .IN2(n1114), .S(n8053), .Q(n11743)
         );
  MUX21X1 U14880 ( .IN1(\mem2[166][18] ), .IN2(n1092), .S(n8053), .Q(n11742)
         );
  MUX21X1 U14881 ( .IN1(\mem2[166][17] ), .IN2(n1070), .S(n8053), .Q(n11741)
         );
  MUX21X1 U14882 ( .IN1(\mem2[166][16] ), .IN2(n1048), .S(n8053), .Q(n11740)
         );
  AND2X1 U14883 ( .IN1(n8044), .IN2(n7118), .Q(n8053) );
  MUX21X1 U14884 ( .IN1(\mem2[165][23] ), .IN2(n1202), .S(n8054), .Q(n11739)
         );
  MUX21X1 U14885 ( .IN1(\mem2[165][22] ), .IN2(n1180), .S(n8054), .Q(n11738)
         );
  MUX21X1 U14886 ( .IN1(\mem2[165][21] ), .IN2(n1158), .S(n8054), .Q(n11737)
         );
  MUX21X1 U14887 ( .IN1(\mem2[165][20] ), .IN2(n1136), .S(n8054), .Q(n11736)
         );
  MUX21X1 U14888 ( .IN1(\mem2[165][19] ), .IN2(n1114), .S(n8054), .Q(n11735)
         );
  MUX21X1 U14889 ( .IN1(\mem2[165][18] ), .IN2(n1092), .S(n8054), .Q(n11734)
         );
  MUX21X1 U14890 ( .IN1(\mem2[165][17] ), .IN2(n1070), .S(n8054), .Q(n11733)
         );
  MUX21X1 U14891 ( .IN1(\mem2[165][16] ), .IN2(n1048), .S(n8054), .Q(n11732)
         );
  AND2X1 U14892 ( .IN1(n8044), .IN2(n7120), .Q(n8054) );
  MUX21X1 U14893 ( .IN1(\mem2[164][23] ), .IN2(n1202), .S(n8055), .Q(n11731)
         );
  MUX21X1 U14894 ( .IN1(\mem2[164][22] ), .IN2(n1180), .S(n8055), .Q(n11730)
         );
  MUX21X1 U14895 ( .IN1(\mem2[164][21] ), .IN2(n1158), .S(n8055), .Q(n11729)
         );
  MUX21X1 U14896 ( .IN1(\mem2[164][20] ), .IN2(n1136), .S(n8055), .Q(n11728)
         );
  MUX21X1 U14897 ( .IN1(\mem2[164][19] ), .IN2(n1114), .S(n8055), .Q(n11727)
         );
  MUX21X1 U14898 ( .IN1(\mem2[164][18] ), .IN2(n1092), .S(n8055), .Q(n11726)
         );
  MUX21X1 U14899 ( .IN1(\mem2[164][17] ), .IN2(n1070), .S(n8055), .Q(n11725)
         );
  MUX21X1 U14900 ( .IN1(\mem2[164][16] ), .IN2(n1048), .S(n8055), .Q(n11724)
         );
  AND2X1 U14901 ( .IN1(n8044), .IN2(n7122), .Q(n8055) );
  MUX21X1 U14902 ( .IN1(\mem2[163][23] ), .IN2(n1202), .S(n8056), .Q(n11723)
         );
  MUX21X1 U14903 ( .IN1(\mem2[163][22] ), .IN2(n1180), .S(n8056), .Q(n11722)
         );
  MUX21X1 U14904 ( .IN1(\mem2[163][21] ), .IN2(n1158), .S(n8056), .Q(n11721)
         );
  MUX21X1 U14905 ( .IN1(\mem2[163][20] ), .IN2(n1136), .S(n8056), .Q(n11720)
         );
  MUX21X1 U14906 ( .IN1(\mem2[163][19] ), .IN2(n1114), .S(n8056), .Q(n11719)
         );
  MUX21X1 U14907 ( .IN1(\mem2[163][18] ), .IN2(n1092), .S(n8056), .Q(n11718)
         );
  MUX21X1 U14908 ( .IN1(\mem2[163][17] ), .IN2(n1070), .S(n8056), .Q(n11717)
         );
  MUX21X1 U14909 ( .IN1(\mem2[163][16] ), .IN2(n1048), .S(n8056), .Q(n11716)
         );
  AND2X1 U14910 ( .IN1(n8044), .IN2(n7124), .Q(n8056) );
  MUX21X1 U14911 ( .IN1(\mem2[162][23] ), .IN2(n1202), .S(n8057), .Q(n11715)
         );
  MUX21X1 U14912 ( .IN1(\mem2[162][22] ), .IN2(n1180), .S(n8057), .Q(n11714)
         );
  MUX21X1 U14913 ( .IN1(\mem2[162][21] ), .IN2(n1158), .S(n8057), .Q(n11713)
         );
  MUX21X1 U14914 ( .IN1(\mem2[162][20] ), .IN2(n1136), .S(n8057), .Q(n11712)
         );
  MUX21X1 U14915 ( .IN1(\mem2[162][19] ), .IN2(n1114), .S(n8057), .Q(n11711)
         );
  MUX21X1 U14916 ( .IN1(\mem2[162][18] ), .IN2(n1092), .S(n8057), .Q(n11710)
         );
  MUX21X1 U14917 ( .IN1(\mem2[162][17] ), .IN2(n1070), .S(n8057), .Q(n11709)
         );
  MUX21X1 U14918 ( .IN1(\mem2[162][16] ), .IN2(n1048), .S(n8057), .Q(n11708)
         );
  AND2X1 U14919 ( .IN1(n8044), .IN2(n7126), .Q(n8057) );
  MUX21X1 U14920 ( .IN1(\mem2[161][23] ), .IN2(n1202), .S(n8058), .Q(n11707)
         );
  MUX21X1 U14921 ( .IN1(\mem2[161][22] ), .IN2(n1180), .S(n8058), .Q(n11706)
         );
  MUX21X1 U14922 ( .IN1(\mem2[161][21] ), .IN2(n1158), .S(n8058), .Q(n11705)
         );
  MUX21X1 U14923 ( .IN1(\mem2[161][20] ), .IN2(n1136), .S(n8058), .Q(n11704)
         );
  MUX21X1 U14924 ( .IN1(\mem2[161][19] ), .IN2(n1114), .S(n8058), .Q(n11703)
         );
  MUX21X1 U14925 ( .IN1(\mem2[161][18] ), .IN2(n1092), .S(n8058), .Q(n11702)
         );
  MUX21X1 U14926 ( .IN1(\mem2[161][17] ), .IN2(n1070), .S(n8058), .Q(n11701)
         );
  MUX21X1 U14927 ( .IN1(\mem2[161][16] ), .IN2(n1048), .S(n8058), .Q(n11700)
         );
  AND2X1 U14928 ( .IN1(n8044), .IN2(n7128), .Q(n8058) );
  MUX21X1 U14929 ( .IN1(\mem2[160][23] ), .IN2(n1202), .S(n8059), .Q(n11699)
         );
  MUX21X1 U14930 ( .IN1(\mem2[160][22] ), .IN2(n1180), .S(n8059), .Q(n11698)
         );
  MUX21X1 U14931 ( .IN1(\mem2[160][21] ), .IN2(n1158), .S(n8059), .Q(n11697)
         );
  MUX21X1 U14932 ( .IN1(\mem2[160][20] ), .IN2(n1136), .S(n8059), .Q(n11696)
         );
  MUX21X1 U14933 ( .IN1(\mem2[160][19] ), .IN2(n1114), .S(n8059), .Q(n11695)
         );
  MUX21X1 U14934 ( .IN1(\mem2[160][18] ), .IN2(n1092), .S(n8059), .Q(n11694)
         );
  MUX21X1 U14935 ( .IN1(\mem2[160][17] ), .IN2(n1070), .S(n8059), .Q(n11693)
         );
  MUX21X1 U14936 ( .IN1(\mem2[160][16] ), .IN2(n1048), .S(n8059), .Q(n11692)
         );
  AND2X1 U14937 ( .IN1(n8044), .IN2(n7130), .Q(n8059) );
  AND2X1 U14938 ( .IN1(n7966), .IN2(n7222), .Q(n8044) );
  AND2X1 U14939 ( .IN1(n8042), .IN2(n7986), .Q(n7222) );
  MUX21X1 U14940 ( .IN1(\mem2[159][23] ), .IN2(n1203), .S(n8060), .Q(n11691)
         );
  MUX21X1 U14941 ( .IN1(\mem2[159][22] ), .IN2(n1181), .S(n8060), .Q(n11690)
         );
  MUX21X1 U14942 ( .IN1(\mem2[159][21] ), .IN2(n1159), .S(n8060), .Q(n11689)
         );
  MUX21X1 U14943 ( .IN1(\mem2[159][20] ), .IN2(n1137), .S(n8060), .Q(n11688)
         );
  MUX21X1 U14944 ( .IN1(\mem2[159][19] ), .IN2(n1115), .S(n8060), .Q(n11687)
         );
  MUX21X1 U14945 ( .IN1(\mem2[159][18] ), .IN2(n1093), .S(n8060), .Q(n11686)
         );
  MUX21X1 U14946 ( .IN1(\mem2[159][17] ), .IN2(n1071), .S(n8060), .Q(n11685)
         );
  MUX21X1 U14947 ( .IN1(\mem2[159][16] ), .IN2(n1049), .S(n8060), .Q(n11684)
         );
  AND2X1 U14948 ( .IN1(n8061), .IN2(n7099), .Q(n8060) );
  MUX21X1 U14949 ( .IN1(\mem2[158][23] ), .IN2(n1203), .S(n8062), .Q(n11683)
         );
  MUX21X1 U14950 ( .IN1(\mem2[158][22] ), .IN2(n1181), .S(n8062), .Q(n11682)
         );
  MUX21X1 U14951 ( .IN1(\mem2[158][21] ), .IN2(n1159), .S(n8062), .Q(n11681)
         );
  MUX21X1 U14952 ( .IN1(\mem2[158][20] ), .IN2(n1137), .S(n8062), .Q(n11680)
         );
  MUX21X1 U14953 ( .IN1(\mem2[158][19] ), .IN2(n1115), .S(n8062), .Q(n11679)
         );
  MUX21X1 U14954 ( .IN1(\mem2[158][18] ), .IN2(n1093), .S(n8062), .Q(n11678)
         );
  MUX21X1 U14955 ( .IN1(\mem2[158][17] ), .IN2(n1071), .S(n8062), .Q(n11677)
         );
  MUX21X1 U14956 ( .IN1(\mem2[158][16] ), .IN2(n1049), .S(n8062), .Q(n11676)
         );
  AND2X1 U14957 ( .IN1(n8061), .IN2(n7102), .Q(n8062) );
  MUX21X1 U14958 ( .IN1(\mem2[157][23] ), .IN2(n1203), .S(n8063), .Q(n11675)
         );
  MUX21X1 U14959 ( .IN1(\mem2[157][22] ), .IN2(n1181), .S(n8063), .Q(n11674)
         );
  MUX21X1 U14960 ( .IN1(\mem2[157][21] ), .IN2(n1159), .S(n8063), .Q(n11673)
         );
  MUX21X1 U14961 ( .IN1(\mem2[157][20] ), .IN2(n1137), .S(n8063), .Q(n11672)
         );
  MUX21X1 U14962 ( .IN1(\mem2[157][19] ), .IN2(n1115), .S(n8063), .Q(n11671)
         );
  MUX21X1 U14963 ( .IN1(\mem2[157][18] ), .IN2(n1093), .S(n8063), .Q(n11670)
         );
  MUX21X1 U14964 ( .IN1(\mem2[157][17] ), .IN2(n1071), .S(n8063), .Q(n11669)
         );
  MUX21X1 U14965 ( .IN1(\mem2[157][16] ), .IN2(n1049), .S(n8063), .Q(n11668)
         );
  AND2X1 U14966 ( .IN1(n8061), .IN2(n7104), .Q(n8063) );
  MUX21X1 U14967 ( .IN1(\mem2[156][23] ), .IN2(n1203), .S(n8064), .Q(n11667)
         );
  MUX21X1 U14968 ( .IN1(\mem2[156][22] ), .IN2(n1181), .S(n8064), .Q(n11666)
         );
  MUX21X1 U14969 ( .IN1(\mem2[156][21] ), .IN2(n1159), .S(n8064), .Q(n11665)
         );
  MUX21X1 U14970 ( .IN1(\mem2[156][20] ), .IN2(n1137), .S(n8064), .Q(n11664)
         );
  MUX21X1 U14971 ( .IN1(\mem2[156][19] ), .IN2(n1115), .S(n8064), .Q(n11663)
         );
  MUX21X1 U14972 ( .IN1(\mem2[156][18] ), .IN2(n1093), .S(n8064), .Q(n11662)
         );
  MUX21X1 U14973 ( .IN1(\mem2[156][17] ), .IN2(n1071), .S(n8064), .Q(n11661)
         );
  MUX21X1 U14974 ( .IN1(\mem2[156][16] ), .IN2(n1049), .S(n8064), .Q(n11660)
         );
  AND2X1 U14975 ( .IN1(n8061), .IN2(n7106), .Q(n8064) );
  MUX21X1 U14976 ( .IN1(\mem2[155][23] ), .IN2(n1203), .S(n8065), .Q(n11659)
         );
  MUX21X1 U14977 ( .IN1(\mem2[155][22] ), .IN2(n1181), .S(n8065), .Q(n11658)
         );
  MUX21X1 U14978 ( .IN1(\mem2[155][21] ), .IN2(n1159), .S(n8065), .Q(n11657)
         );
  MUX21X1 U14979 ( .IN1(\mem2[155][20] ), .IN2(n1137), .S(n8065), .Q(n11656)
         );
  MUX21X1 U14980 ( .IN1(\mem2[155][19] ), .IN2(n1115), .S(n8065), .Q(n11655)
         );
  MUX21X1 U14981 ( .IN1(\mem2[155][18] ), .IN2(n1093), .S(n8065), .Q(n11654)
         );
  MUX21X1 U14982 ( .IN1(\mem2[155][17] ), .IN2(n1071), .S(n8065), .Q(n11653)
         );
  MUX21X1 U14983 ( .IN1(\mem2[155][16] ), .IN2(n1049), .S(n8065), .Q(n11652)
         );
  AND2X1 U14984 ( .IN1(n8061), .IN2(n7108), .Q(n8065) );
  MUX21X1 U14985 ( .IN1(\mem2[154][23] ), .IN2(n1203), .S(n8066), .Q(n11651)
         );
  MUX21X1 U14986 ( .IN1(\mem2[154][22] ), .IN2(n1181), .S(n8066), .Q(n11650)
         );
  MUX21X1 U14987 ( .IN1(\mem2[154][21] ), .IN2(n1159), .S(n8066), .Q(n11649)
         );
  MUX21X1 U14988 ( .IN1(\mem2[154][20] ), .IN2(n1137), .S(n8066), .Q(n11648)
         );
  MUX21X1 U14989 ( .IN1(\mem2[154][19] ), .IN2(n1115), .S(n8066), .Q(n11647)
         );
  MUX21X1 U14990 ( .IN1(\mem2[154][18] ), .IN2(n1093), .S(n8066), .Q(n11646)
         );
  MUX21X1 U14991 ( .IN1(\mem2[154][17] ), .IN2(n1071), .S(n8066), .Q(n11645)
         );
  MUX21X1 U14992 ( .IN1(\mem2[154][16] ), .IN2(n1049), .S(n8066), .Q(n11644)
         );
  AND2X1 U14993 ( .IN1(n8061), .IN2(n7110), .Q(n8066) );
  MUX21X1 U14994 ( .IN1(\mem2[153][23] ), .IN2(n1203), .S(n8067), .Q(n11643)
         );
  MUX21X1 U14995 ( .IN1(\mem2[153][22] ), .IN2(n1181), .S(n8067), .Q(n11642)
         );
  MUX21X1 U14996 ( .IN1(\mem2[153][21] ), .IN2(n1159), .S(n8067), .Q(n11641)
         );
  MUX21X1 U14997 ( .IN1(\mem2[153][20] ), .IN2(n1137), .S(n8067), .Q(n11640)
         );
  MUX21X1 U14998 ( .IN1(\mem2[153][19] ), .IN2(n1115), .S(n8067), .Q(n11639)
         );
  MUX21X1 U14999 ( .IN1(\mem2[153][18] ), .IN2(n1093), .S(n8067), .Q(n11638)
         );
  MUX21X1 U15000 ( .IN1(\mem2[153][17] ), .IN2(n1071), .S(n8067), .Q(n11637)
         );
  MUX21X1 U15001 ( .IN1(\mem2[153][16] ), .IN2(n1049), .S(n8067), .Q(n11636)
         );
  AND2X1 U15002 ( .IN1(n8061), .IN2(n7112), .Q(n8067) );
  MUX21X1 U15003 ( .IN1(\mem2[152][23] ), .IN2(n1203), .S(n8068), .Q(n11635)
         );
  MUX21X1 U15004 ( .IN1(\mem2[152][22] ), .IN2(n1181), .S(n8068), .Q(n11634)
         );
  MUX21X1 U15005 ( .IN1(\mem2[152][21] ), .IN2(n1159), .S(n8068), .Q(n11633)
         );
  MUX21X1 U15006 ( .IN1(\mem2[152][20] ), .IN2(n1137), .S(n8068), .Q(n11632)
         );
  MUX21X1 U15007 ( .IN1(\mem2[152][19] ), .IN2(n1115), .S(n8068), .Q(n11631)
         );
  MUX21X1 U15008 ( .IN1(\mem2[152][18] ), .IN2(n1093), .S(n8068), .Q(n11630)
         );
  MUX21X1 U15009 ( .IN1(\mem2[152][17] ), .IN2(n1071), .S(n8068), .Q(n11629)
         );
  MUX21X1 U15010 ( .IN1(\mem2[152][16] ), .IN2(n1049), .S(n8068), .Q(n11628)
         );
  AND2X1 U15011 ( .IN1(n8061), .IN2(n7114), .Q(n8068) );
  MUX21X1 U15012 ( .IN1(\mem2[151][23] ), .IN2(n1203), .S(n8069), .Q(n11627)
         );
  MUX21X1 U15013 ( .IN1(\mem2[151][22] ), .IN2(n1181), .S(n8069), .Q(n11626)
         );
  MUX21X1 U15014 ( .IN1(\mem2[151][21] ), .IN2(n1159), .S(n8069), .Q(n11625)
         );
  MUX21X1 U15015 ( .IN1(\mem2[151][20] ), .IN2(n1137), .S(n8069), .Q(n11624)
         );
  MUX21X1 U15016 ( .IN1(\mem2[151][19] ), .IN2(n1115), .S(n8069), .Q(n11623)
         );
  MUX21X1 U15017 ( .IN1(\mem2[151][18] ), .IN2(n1093), .S(n8069), .Q(n11622)
         );
  MUX21X1 U15018 ( .IN1(\mem2[151][17] ), .IN2(n1071), .S(n8069), .Q(n11621)
         );
  MUX21X1 U15019 ( .IN1(\mem2[151][16] ), .IN2(n1049), .S(n8069), .Q(n11620)
         );
  AND2X1 U15020 ( .IN1(n8061), .IN2(n7116), .Q(n8069) );
  MUX21X1 U15021 ( .IN1(\mem2[150][23] ), .IN2(n1203), .S(n8070), .Q(n11619)
         );
  MUX21X1 U15022 ( .IN1(\mem2[150][22] ), .IN2(n1181), .S(n8070), .Q(n11618)
         );
  MUX21X1 U15023 ( .IN1(\mem2[150][21] ), .IN2(n1159), .S(n8070), .Q(n11617)
         );
  MUX21X1 U15024 ( .IN1(\mem2[150][20] ), .IN2(n1137), .S(n8070), .Q(n11616)
         );
  MUX21X1 U15025 ( .IN1(\mem2[150][19] ), .IN2(n1115), .S(n8070), .Q(n11615)
         );
  MUX21X1 U15026 ( .IN1(\mem2[150][18] ), .IN2(n1093), .S(n8070), .Q(n11614)
         );
  MUX21X1 U15027 ( .IN1(\mem2[150][17] ), .IN2(n1071), .S(n8070), .Q(n11613)
         );
  MUX21X1 U15028 ( .IN1(\mem2[150][16] ), .IN2(n1049), .S(n8070), .Q(n11612)
         );
  AND2X1 U15029 ( .IN1(n8061), .IN2(n7118), .Q(n8070) );
  MUX21X1 U15030 ( .IN1(\mem2[149][23] ), .IN2(n1203), .S(n8071), .Q(n11611)
         );
  MUX21X1 U15031 ( .IN1(\mem2[149][22] ), .IN2(n1181), .S(n8071), .Q(n11610)
         );
  MUX21X1 U15032 ( .IN1(\mem2[149][21] ), .IN2(n1159), .S(n8071), .Q(n11609)
         );
  MUX21X1 U15033 ( .IN1(\mem2[149][20] ), .IN2(n1137), .S(n8071), .Q(n11608)
         );
  MUX21X1 U15034 ( .IN1(\mem2[149][19] ), .IN2(n1115), .S(n8071), .Q(n11607)
         );
  MUX21X1 U15035 ( .IN1(\mem2[149][18] ), .IN2(n1093), .S(n8071), .Q(n11606)
         );
  MUX21X1 U15036 ( .IN1(\mem2[149][17] ), .IN2(n1071), .S(n8071), .Q(n11605)
         );
  MUX21X1 U15037 ( .IN1(\mem2[149][16] ), .IN2(n1049), .S(n8071), .Q(n11604)
         );
  AND2X1 U15038 ( .IN1(n8061), .IN2(n7120), .Q(n8071) );
  MUX21X1 U15039 ( .IN1(\mem2[148][23] ), .IN2(n1203), .S(n8072), .Q(n11603)
         );
  MUX21X1 U15040 ( .IN1(\mem2[148][22] ), .IN2(n1181), .S(n8072), .Q(n11602)
         );
  MUX21X1 U15041 ( .IN1(\mem2[148][21] ), .IN2(n1159), .S(n8072), .Q(n11601)
         );
  MUX21X1 U15042 ( .IN1(\mem2[148][20] ), .IN2(n1137), .S(n8072), .Q(n11600)
         );
  MUX21X1 U15043 ( .IN1(\mem2[148][19] ), .IN2(n1115), .S(n8072), .Q(n11599)
         );
  MUX21X1 U15044 ( .IN1(\mem2[148][18] ), .IN2(n1093), .S(n8072), .Q(n11598)
         );
  MUX21X1 U15045 ( .IN1(\mem2[148][17] ), .IN2(n1071), .S(n8072), .Q(n11597)
         );
  MUX21X1 U15046 ( .IN1(\mem2[148][16] ), .IN2(n1049), .S(n8072), .Q(n11596)
         );
  AND2X1 U15047 ( .IN1(n8061), .IN2(n7122), .Q(n8072) );
  MUX21X1 U15048 ( .IN1(\mem2[147][23] ), .IN2(n1204), .S(n8073), .Q(n11595)
         );
  MUX21X1 U15049 ( .IN1(\mem2[147][22] ), .IN2(n1182), .S(n8073), .Q(n11594)
         );
  MUX21X1 U15050 ( .IN1(\mem2[147][21] ), .IN2(n1160), .S(n8073), .Q(n11593)
         );
  MUX21X1 U15051 ( .IN1(\mem2[147][20] ), .IN2(n1138), .S(n8073), .Q(n11592)
         );
  MUX21X1 U15052 ( .IN1(\mem2[147][19] ), .IN2(n1116), .S(n8073), .Q(n11591)
         );
  MUX21X1 U15053 ( .IN1(\mem2[147][18] ), .IN2(n1094), .S(n8073), .Q(n11590)
         );
  MUX21X1 U15054 ( .IN1(\mem2[147][17] ), .IN2(n1072), .S(n8073), .Q(n11589)
         );
  MUX21X1 U15055 ( .IN1(\mem2[147][16] ), .IN2(n1050), .S(n8073), .Q(n11588)
         );
  AND2X1 U15056 ( .IN1(n8061), .IN2(n7124), .Q(n8073) );
  MUX21X1 U15057 ( .IN1(\mem2[146][23] ), .IN2(n1204), .S(n8074), .Q(n11587)
         );
  MUX21X1 U15058 ( .IN1(\mem2[146][22] ), .IN2(n1182), .S(n8074), .Q(n11586)
         );
  MUX21X1 U15059 ( .IN1(\mem2[146][21] ), .IN2(n1160), .S(n8074), .Q(n11585)
         );
  MUX21X1 U15060 ( .IN1(\mem2[146][20] ), .IN2(n1138), .S(n8074), .Q(n11584)
         );
  MUX21X1 U15061 ( .IN1(\mem2[146][19] ), .IN2(n1116), .S(n8074), .Q(n11583)
         );
  MUX21X1 U15062 ( .IN1(\mem2[146][18] ), .IN2(n1094), .S(n8074), .Q(n11582)
         );
  MUX21X1 U15063 ( .IN1(\mem2[146][17] ), .IN2(n1072), .S(n8074), .Q(n11581)
         );
  MUX21X1 U15064 ( .IN1(\mem2[146][16] ), .IN2(n1050), .S(n8074), .Q(n11580)
         );
  AND2X1 U15065 ( .IN1(n8061), .IN2(n7126), .Q(n8074) );
  MUX21X1 U15066 ( .IN1(\mem2[145][23] ), .IN2(n1204), .S(n8075), .Q(n11579)
         );
  MUX21X1 U15067 ( .IN1(\mem2[145][22] ), .IN2(n1182), .S(n8075), .Q(n11578)
         );
  MUX21X1 U15068 ( .IN1(\mem2[145][21] ), .IN2(n1160), .S(n8075), .Q(n11577)
         );
  MUX21X1 U15069 ( .IN1(\mem2[145][20] ), .IN2(n1138), .S(n8075), .Q(n11576)
         );
  MUX21X1 U15070 ( .IN1(\mem2[145][19] ), .IN2(n1116), .S(n8075), .Q(n11575)
         );
  MUX21X1 U15071 ( .IN1(\mem2[145][18] ), .IN2(n1094), .S(n8075), .Q(n11574)
         );
  MUX21X1 U15072 ( .IN1(\mem2[145][17] ), .IN2(n1072), .S(n8075), .Q(n11573)
         );
  MUX21X1 U15073 ( .IN1(\mem2[145][16] ), .IN2(n1050), .S(n8075), .Q(n11572)
         );
  AND2X1 U15074 ( .IN1(n8061), .IN2(n7128), .Q(n8075) );
  MUX21X1 U15075 ( .IN1(\mem2[144][23] ), .IN2(n1204), .S(n8076), .Q(n11571)
         );
  MUX21X1 U15076 ( .IN1(\mem2[144][22] ), .IN2(n1182), .S(n8076), .Q(n11570)
         );
  MUX21X1 U15077 ( .IN1(\mem2[144][21] ), .IN2(n1160), .S(n8076), .Q(n11569)
         );
  MUX21X1 U15078 ( .IN1(\mem2[144][20] ), .IN2(n1138), .S(n8076), .Q(n11568)
         );
  MUX21X1 U15079 ( .IN1(\mem2[144][19] ), .IN2(n1116), .S(n8076), .Q(n11567)
         );
  MUX21X1 U15080 ( .IN1(\mem2[144][18] ), .IN2(n1094), .S(n8076), .Q(n11566)
         );
  MUX21X1 U15081 ( .IN1(\mem2[144][17] ), .IN2(n1072), .S(n8076), .Q(n11565)
         );
  MUX21X1 U15082 ( .IN1(\mem2[144][16] ), .IN2(n1050), .S(n8076), .Q(n11564)
         );
  AND2X1 U15083 ( .IN1(n8061), .IN2(n7130), .Q(n8076) );
  AND2X1 U15084 ( .IN1(n7966), .IN2(n7240), .Q(n8061) );
  AND2X1 U15085 ( .IN1(n8042), .IN2(n8004), .Q(n7240) );
  MUX21X1 U15086 ( .IN1(\mem2[143][23] ), .IN2(n1204), .S(n8077), .Q(n11563)
         );
  MUX21X1 U15087 ( .IN1(\mem2[143][22] ), .IN2(n1182), .S(n8077), .Q(n11562)
         );
  MUX21X1 U15088 ( .IN1(\mem2[143][21] ), .IN2(n1160), .S(n8077), .Q(n11561)
         );
  MUX21X1 U15089 ( .IN1(\mem2[143][20] ), .IN2(n1138), .S(n8077), .Q(n11560)
         );
  MUX21X1 U15090 ( .IN1(\mem2[143][19] ), .IN2(n1116), .S(n8077), .Q(n11559)
         );
  MUX21X1 U15091 ( .IN1(\mem2[143][18] ), .IN2(n1094), .S(n8077), .Q(n11558)
         );
  MUX21X1 U15092 ( .IN1(\mem2[143][17] ), .IN2(n1072), .S(n8077), .Q(n11557)
         );
  MUX21X1 U15093 ( .IN1(\mem2[143][16] ), .IN2(n1050), .S(n8077), .Q(n11556)
         );
  AND2X1 U15094 ( .IN1(n8078), .IN2(n7099), .Q(n8077) );
  MUX21X1 U15095 ( .IN1(\mem2[142][23] ), .IN2(n1204), .S(n8079), .Q(n11555)
         );
  MUX21X1 U15096 ( .IN1(\mem2[142][22] ), .IN2(n1182), .S(n8079), .Q(n11554)
         );
  MUX21X1 U15097 ( .IN1(\mem2[142][21] ), .IN2(n1160), .S(n8079), .Q(n11553)
         );
  MUX21X1 U15098 ( .IN1(\mem2[142][20] ), .IN2(n1138), .S(n8079), .Q(n11552)
         );
  MUX21X1 U15099 ( .IN1(\mem2[142][19] ), .IN2(n1116), .S(n8079), .Q(n11551)
         );
  MUX21X1 U15100 ( .IN1(\mem2[142][18] ), .IN2(n1094), .S(n8079), .Q(n11550)
         );
  MUX21X1 U15101 ( .IN1(\mem2[142][17] ), .IN2(n1072), .S(n8079), .Q(n11549)
         );
  MUX21X1 U15102 ( .IN1(\mem2[142][16] ), .IN2(n1050), .S(n8079), .Q(n11548)
         );
  AND2X1 U15103 ( .IN1(n8078), .IN2(n7102), .Q(n8079) );
  MUX21X1 U15104 ( .IN1(\mem2[141][23] ), .IN2(n1204), .S(n8080), .Q(n11547)
         );
  MUX21X1 U15105 ( .IN1(\mem2[141][22] ), .IN2(n1182), .S(n8080), .Q(n11546)
         );
  MUX21X1 U15106 ( .IN1(\mem2[141][21] ), .IN2(n1160), .S(n8080), .Q(n11545)
         );
  MUX21X1 U15107 ( .IN1(\mem2[141][20] ), .IN2(n1138), .S(n8080), .Q(n11544)
         );
  MUX21X1 U15108 ( .IN1(\mem2[141][19] ), .IN2(n1116), .S(n8080), .Q(n11543)
         );
  MUX21X1 U15109 ( .IN1(\mem2[141][18] ), .IN2(n1094), .S(n8080), .Q(n11542)
         );
  MUX21X1 U15110 ( .IN1(\mem2[141][17] ), .IN2(n1072), .S(n8080), .Q(n11541)
         );
  MUX21X1 U15111 ( .IN1(\mem2[141][16] ), .IN2(n1050), .S(n8080), .Q(n11540)
         );
  AND2X1 U15112 ( .IN1(n8078), .IN2(n7104), .Q(n8080) );
  MUX21X1 U15113 ( .IN1(\mem2[140][23] ), .IN2(n1204), .S(n8081), .Q(n11539)
         );
  MUX21X1 U15114 ( .IN1(\mem2[140][22] ), .IN2(n1182), .S(n8081), .Q(n11538)
         );
  MUX21X1 U15115 ( .IN1(\mem2[140][21] ), .IN2(n1160), .S(n8081), .Q(n11537)
         );
  MUX21X1 U15116 ( .IN1(\mem2[140][20] ), .IN2(n1138), .S(n8081), .Q(n11536)
         );
  MUX21X1 U15117 ( .IN1(\mem2[140][19] ), .IN2(n1116), .S(n8081), .Q(n11535)
         );
  MUX21X1 U15118 ( .IN1(\mem2[140][18] ), .IN2(n1094), .S(n8081), .Q(n11534)
         );
  MUX21X1 U15119 ( .IN1(\mem2[140][17] ), .IN2(n1072), .S(n8081), .Q(n11533)
         );
  MUX21X1 U15120 ( .IN1(\mem2[140][16] ), .IN2(n1050), .S(n8081), .Q(n11532)
         );
  AND2X1 U15121 ( .IN1(n8078), .IN2(n7106), .Q(n8081) );
  MUX21X1 U15122 ( .IN1(\mem2[139][23] ), .IN2(n1204), .S(n8082), .Q(n11531)
         );
  MUX21X1 U15123 ( .IN1(\mem2[139][22] ), .IN2(n1182), .S(n8082), .Q(n11530)
         );
  MUX21X1 U15124 ( .IN1(\mem2[139][21] ), .IN2(n1160), .S(n8082), .Q(n11529)
         );
  MUX21X1 U15125 ( .IN1(\mem2[139][20] ), .IN2(n1138), .S(n8082), .Q(n11528)
         );
  MUX21X1 U15126 ( .IN1(\mem2[139][19] ), .IN2(n1116), .S(n8082), .Q(n11527)
         );
  MUX21X1 U15127 ( .IN1(\mem2[139][18] ), .IN2(n1094), .S(n8082), .Q(n11526)
         );
  MUX21X1 U15128 ( .IN1(\mem2[139][17] ), .IN2(n1072), .S(n8082), .Q(n11525)
         );
  MUX21X1 U15129 ( .IN1(\mem2[139][16] ), .IN2(n1050), .S(n8082), .Q(n11524)
         );
  AND2X1 U15130 ( .IN1(n8078), .IN2(n7108), .Q(n8082) );
  MUX21X1 U15131 ( .IN1(\mem2[138][23] ), .IN2(n1204), .S(n8083), .Q(n11523)
         );
  MUX21X1 U15132 ( .IN1(\mem2[138][22] ), .IN2(n1182), .S(n8083), .Q(n11522)
         );
  MUX21X1 U15133 ( .IN1(\mem2[138][21] ), .IN2(n1160), .S(n8083), .Q(n11521)
         );
  MUX21X1 U15134 ( .IN1(\mem2[138][20] ), .IN2(n1138), .S(n8083), .Q(n11520)
         );
  MUX21X1 U15135 ( .IN1(\mem2[138][19] ), .IN2(n1116), .S(n8083), .Q(n11519)
         );
  MUX21X1 U15136 ( .IN1(\mem2[138][18] ), .IN2(n1094), .S(n8083), .Q(n11518)
         );
  MUX21X1 U15137 ( .IN1(\mem2[138][17] ), .IN2(n1072), .S(n8083), .Q(n11517)
         );
  MUX21X1 U15138 ( .IN1(\mem2[138][16] ), .IN2(n1050), .S(n8083), .Q(n11516)
         );
  AND2X1 U15139 ( .IN1(n8078), .IN2(n7110), .Q(n8083) );
  MUX21X1 U15140 ( .IN1(\mem2[137][23] ), .IN2(n1204), .S(n8084), .Q(n11515)
         );
  MUX21X1 U15141 ( .IN1(\mem2[137][22] ), .IN2(n1182), .S(n8084), .Q(n11514)
         );
  MUX21X1 U15142 ( .IN1(\mem2[137][21] ), .IN2(n1160), .S(n8084), .Q(n11513)
         );
  MUX21X1 U15143 ( .IN1(\mem2[137][20] ), .IN2(n1138), .S(n8084), .Q(n11512)
         );
  MUX21X1 U15144 ( .IN1(\mem2[137][19] ), .IN2(n1116), .S(n8084), .Q(n11511)
         );
  MUX21X1 U15145 ( .IN1(\mem2[137][18] ), .IN2(n1094), .S(n8084), .Q(n11510)
         );
  MUX21X1 U15146 ( .IN1(\mem2[137][17] ), .IN2(n1072), .S(n8084), .Q(n11509)
         );
  MUX21X1 U15147 ( .IN1(\mem2[137][16] ), .IN2(n1050), .S(n8084), .Q(n11508)
         );
  AND2X1 U15148 ( .IN1(n8078), .IN2(n7112), .Q(n8084) );
  MUX21X1 U15149 ( .IN1(\mem2[136][23] ), .IN2(n1204), .S(n8085), .Q(n11507)
         );
  MUX21X1 U15150 ( .IN1(\mem2[136][22] ), .IN2(n1182), .S(n8085), .Q(n11506)
         );
  MUX21X1 U15151 ( .IN1(\mem2[136][21] ), .IN2(n1160), .S(n8085), .Q(n11505)
         );
  MUX21X1 U15152 ( .IN1(\mem2[136][20] ), .IN2(n1138), .S(n8085), .Q(n11504)
         );
  MUX21X1 U15153 ( .IN1(\mem2[136][19] ), .IN2(n1116), .S(n8085), .Q(n11503)
         );
  MUX21X1 U15154 ( .IN1(\mem2[136][18] ), .IN2(n1094), .S(n8085), .Q(n11502)
         );
  MUX21X1 U15155 ( .IN1(\mem2[136][17] ), .IN2(n1072), .S(n8085), .Q(n11501)
         );
  MUX21X1 U15156 ( .IN1(\mem2[136][16] ), .IN2(n1050), .S(n8085), .Q(n11500)
         );
  AND2X1 U15157 ( .IN1(n8078), .IN2(n7114), .Q(n8085) );
  MUX21X1 U15158 ( .IN1(\mem2[135][23] ), .IN2(n1205), .S(n8086), .Q(n11499)
         );
  MUX21X1 U15159 ( .IN1(\mem2[135][22] ), .IN2(n1183), .S(n8086), .Q(n11498)
         );
  MUX21X1 U15160 ( .IN1(\mem2[135][21] ), .IN2(n1161), .S(n8086), .Q(n11497)
         );
  MUX21X1 U15161 ( .IN1(\mem2[135][20] ), .IN2(n1139), .S(n8086), .Q(n11496)
         );
  MUX21X1 U15162 ( .IN1(\mem2[135][19] ), .IN2(n1117), .S(n8086), .Q(n11495)
         );
  MUX21X1 U15163 ( .IN1(\mem2[135][18] ), .IN2(n1095), .S(n8086), .Q(n11494)
         );
  MUX21X1 U15164 ( .IN1(\mem2[135][17] ), .IN2(n1073), .S(n8086), .Q(n11493)
         );
  MUX21X1 U15165 ( .IN1(\mem2[135][16] ), .IN2(n1051), .S(n8086), .Q(n11492)
         );
  AND2X1 U15166 ( .IN1(n8078), .IN2(n7116), .Q(n8086) );
  MUX21X1 U15167 ( .IN1(\mem2[134][23] ), .IN2(n1205), .S(n8087), .Q(n11491)
         );
  MUX21X1 U15168 ( .IN1(\mem2[134][22] ), .IN2(n1183), .S(n8087), .Q(n11490)
         );
  MUX21X1 U15169 ( .IN1(\mem2[134][21] ), .IN2(n1161), .S(n8087), .Q(n11489)
         );
  MUX21X1 U15170 ( .IN1(\mem2[134][20] ), .IN2(n1139), .S(n8087), .Q(n11488)
         );
  MUX21X1 U15171 ( .IN1(\mem2[134][19] ), .IN2(n1117), .S(n8087), .Q(n11487)
         );
  MUX21X1 U15172 ( .IN1(\mem2[134][18] ), .IN2(n1095), .S(n8087), .Q(n11486)
         );
  MUX21X1 U15173 ( .IN1(\mem2[134][17] ), .IN2(n1073), .S(n8087), .Q(n11485)
         );
  MUX21X1 U15174 ( .IN1(\mem2[134][16] ), .IN2(n1051), .S(n8087), .Q(n11484)
         );
  AND2X1 U15175 ( .IN1(n8078), .IN2(n7118), .Q(n8087) );
  MUX21X1 U15176 ( .IN1(\mem2[133][23] ), .IN2(n1205), .S(n8088), .Q(n11483)
         );
  MUX21X1 U15177 ( .IN1(\mem2[133][22] ), .IN2(n1183), .S(n8088), .Q(n11482)
         );
  MUX21X1 U15178 ( .IN1(\mem2[133][21] ), .IN2(n1161), .S(n8088), .Q(n11481)
         );
  MUX21X1 U15179 ( .IN1(\mem2[133][20] ), .IN2(n1139), .S(n8088), .Q(n11480)
         );
  MUX21X1 U15180 ( .IN1(\mem2[133][19] ), .IN2(n1117), .S(n8088), .Q(n11479)
         );
  MUX21X1 U15181 ( .IN1(\mem2[133][18] ), .IN2(n1095), .S(n8088), .Q(n11478)
         );
  MUX21X1 U15182 ( .IN1(\mem2[133][17] ), .IN2(n1073), .S(n8088), .Q(n11477)
         );
  MUX21X1 U15183 ( .IN1(\mem2[133][16] ), .IN2(n1051), .S(n8088), .Q(n11476)
         );
  AND2X1 U15184 ( .IN1(n8078), .IN2(n7120), .Q(n8088) );
  MUX21X1 U15185 ( .IN1(\mem2[132][23] ), .IN2(n1205), .S(n8089), .Q(n11475)
         );
  MUX21X1 U15186 ( .IN1(\mem2[132][22] ), .IN2(n1183), .S(n8089), .Q(n11474)
         );
  MUX21X1 U15187 ( .IN1(\mem2[132][21] ), .IN2(n1161), .S(n8089), .Q(n11473)
         );
  MUX21X1 U15188 ( .IN1(\mem2[132][20] ), .IN2(n1139), .S(n8089), .Q(n11472)
         );
  MUX21X1 U15189 ( .IN1(\mem2[132][19] ), .IN2(n1117), .S(n8089), .Q(n11471)
         );
  MUX21X1 U15190 ( .IN1(\mem2[132][18] ), .IN2(n1095), .S(n8089), .Q(n11470)
         );
  MUX21X1 U15191 ( .IN1(\mem2[132][17] ), .IN2(n1073), .S(n8089), .Q(n11469)
         );
  MUX21X1 U15192 ( .IN1(\mem2[132][16] ), .IN2(n1051), .S(n8089), .Q(n11468)
         );
  AND2X1 U15193 ( .IN1(n8078), .IN2(n7122), .Q(n8089) );
  MUX21X1 U15194 ( .IN1(\mem2[131][23] ), .IN2(n1205), .S(n8090), .Q(n11467)
         );
  MUX21X1 U15195 ( .IN1(\mem2[131][22] ), .IN2(n1183), .S(n8090), .Q(n11466)
         );
  MUX21X1 U15196 ( .IN1(\mem2[131][21] ), .IN2(n1161), .S(n8090), .Q(n11465)
         );
  MUX21X1 U15197 ( .IN1(\mem2[131][20] ), .IN2(n1139), .S(n8090), .Q(n11464)
         );
  MUX21X1 U15198 ( .IN1(\mem2[131][19] ), .IN2(n1117), .S(n8090), .Q(n11463)
         );
  MUX21X1 U15199 ( .IN1(\mem2[131][18] ), .IN2(n1095), .S(n8090), .Q(n11462)
         );
  MUX21X1 U15200 ( .IN1(\mem2[131][17] ), .IN2(n1073), .S(n8090), .Q(n11461)
         );
  MUX21X1 U15201 ( .IN1(\mem2[131][16] ), .IN2(n1051), .S(n8090), .Q(n11460)
         );
  AND2X1 U15202 ( .IN1(n8078), .IN2(n7124), .Q(n8090) );
  MUX21X1 U15203 ( .IN1(\mem2[130][23] ), .IN2(n1205), .S(n8091), .Q(n11459)
         );
  MUX21X1 U15204 ( .IN1(\mem2[130][22] ), .IN2(n1183), .S(n8091), .Q(n11458)
         );
  MUX21X1 U15205 ( .IN1(\mem2[130][21] ), .IN2(n1161), .S(n8091), .Q(n11457)
         );
  MUX21X1 U15206 ( .IN1(\mem2[130][20] ), .IN2(n1139), .S(n8091), .Q(n11456)
         );
  MUX21X1 U15207 ( .IN1(\mem2[130][19] ), .IN2(n1117), .S(n8091), .Q(n11455)
         );
  MUX21X1 U15208 ( .IN1(\mem2[130][18] ), .IN2(n1095), .S(n8091), .Q(n11454)
         );
  MUX21X1 U15209 ( .IN1(\mem2[130][17] ), .IN2(n1073), .S(n8091), .Q(n11453)
         );
  MUX21X1 U15210 ( .IN1(\mem2[130][16] ), .IN2(n1051), .S(n8091), .Q(n11452)
         );
  AND2X1 U15211 ( .IN1(n8078), .IN2(n7126), .Q(n8091) );
  MUX21X1 U15212 ( .IN1(\mem2[129][23] ), .IN2(n1205), .S(n8092), .Q(n11451)
         );
  MUX21X1 U15213 ( .IN1(\mem2[129][22] ), .IN2(n1183), .S(n8092), .Q(n11450)
         );
  MUX21X1 U15214 ( .IN1(\mem2[129][21] ), .IN2(n1161), .S(n8092), .Q(n11449)
         );
  MUX21X1 U15215 ( .IN1(\mem2[129][20] ), .IN2(n1139), .S(n8092), .Q(n11448)
         );
  MUX21X1 U15216 ( .IN1(\mem2[129][19] ), .IN2(n1117), .S(n8092), .Q(n11447)
         );
  MUX21X1 U15217 ( .IN1(\mem2[129][18] ), .IN2(n1095), .S(n8092), .Q(n11446)
         );
  MUX21X1 U15218 ( .IN1(\mem2[129][17] ), .IN2(n1073), .S(n8092), .Q(n11445)
         );
  MUX21X1 U15219 ( .IN1(\mem2[129][16] ), .IN2(n1051), .S(n8092), .Q(n11444)
         );
  AND2X1 U15220 ( .IN1(n8078), .IN2(n7128), .Q(n8092) );
  MUX21X1 U15221 ( .IN1(\mem2[128][23] ), .IN2(n1205), .S(n8093), .Q(n11443)
         );
  MUX21X1 U15222 ( .IN1(\mem2[128][22] ), .IN2(n1183), .S(n8093), .Q(n11442)
         );
  MUX21X1 U15223 ( .IN1(\mem2[128][21] ), .IN2(n1161), .S(n8093), .Q(n11441)
         );
  MUX21X1 U15224 ( .IN1(\mem2[128][20] ), .IN2(n1139), .S(n8093), .Q(n11440)
         );
  MUX21X1 U15225 ( .IN1(\mem2[128][19] ), .IN2(n1117), .S(n8093), .Q(n11439)
         );
  MUX21X1 U15226 ( .IN1(\mem2[128][18] ), .IN2(n1095), .S(n8093), .Q(n11438)
         );
  MUX21X1 U15227 ( .IN1(\mem2[128][17] ), .IN2(n1073), .S(n8093), .Q(n11437)
         );
  MUX21X1 U15228 ( .IN1(\mem2[128][16] ), .IN2(n1051), .S(n8093), .Q(n11436)
         );
  AND2X1 U15229 ( .IN1(n8078), .IN2(n7130), .Q(n8093) );
  AND2X1 U15230 ( .IN1(n7966), .IN2(n7258), .Q(n8078) );
  AND2X1 U15231 ( .IN1(n8042), .IN2(n8022), .Q(n7258) );
  NOR2X0 U15232 ( .IN1(n8023), .IN2(addr[6]), .QN(n8042) );
  INVX0 U15233 ( .INP(addr[7]), .ZN(n8023) );
  MUX21X1 U15234 ( .IN1(\mem2[127][23] ), .IN2(n1205), .S(n8094), .Q(n11435)
         );
  MUX21X1 U15235 ( .IN1(\mem2[127][22] ), .IN2(n1183), .S(n8094), .Q(n11434)
         );
  MUX21X1 U15236 ( .IN1(\mem2[127][21] ), .IN2(n1161), .S(n8094), .Q(n11433)
         );
  MUX21X1 U15237 ( .IN1(\mem2[127][20] ), .IN2(n1139), .S(n8094), .Q(n11432)
         );
  MUX21X1 U15238 ( .IN1(\mem2[127][19] ), .IN2(n1117), .S(n8094), .Q(n11431)
         );
  MUX21X1 U15239 ( .IN1(\mem2[127][18] ), .IN2(n1095), .S(n8094), .Q(n11430)
         );
  MUX21X1 U15240 ( .IN1(\mem2[127][17] ), .IN2(n1073), .S(n8094), .Q(n11429)
         );
  MUX21X1 U15241 ( .IN1(\mem2[127][16] ), .IN2(n1051), .S(n8094), .Q(n11428)
         );
  AND2X1 U15242 ( .IN1(n8095), .IN2(n7099), .Q(n8094) );
  MUX21X1 U15243 ( .IN1(\mem2[126][23] ), .IN2(n1205), .S(n8096), .Q(n11427)
         );
  MUX21X1 U15244 ( .IN1(\mem2[126][22] ), .IN2(n1183), .S(n8096), .Q(n11426)
         );
  MUX21X1 U15245 ( .IN1(\mem2[126][21] ), .IN2(n1161), .S(n8096), .Q(n11425)
         );
  MUX21X1 U15246 ( .IN1(\mem2[126][20] ), .IN2(n1139), .S(n8096), .Q(n11424)
         );
  MUX21X1 U15247 ( .IN1(\mem2[126][19] ), .IN2(n1117), .S(n8096), .Q(n11423)
         );
  MUX21X1 U15248 ( .IN1(\mem2[126][18] ), .IN2(n1095), .S(n8096), .Q(n11422)
         );
  MUX21X1 U15249 ( .IN1(\mem2[126][17] ), .IN2(n1073), .S(n8096), .Q(n11421)
         );
  MUX21X1 U15250 ( .IN1(\mem2[126][16] ), .IN2(n1051), .S(n8096), .Q(n11420)
         );
  AND2X1 U15251 ( .IN1(n8095), .IN2(n7102), .Q(n8096) );
  MUX21X1 U15252 ( .IN1(\mem2[125][23] ), .IN2(n1205), .S(n8097), .Q(n11419)
         );
  MUX21X1 U15253 ( .IN1(\mem2[125][22] ), .IN2(n1183), .S(n8097), .Q(n11418)
         );
  MUX21X1 U15254 ( .IN1(\mem2[125][21] ), .IN2(n1161), .S(n8097), .Q(n11417)
         );
  MUX21X1 U15255 ( .IN1(\mem2[125][20] ), .IN2(n1139), .S(n8097), .Q(n11416)
         );
  MUX21X1 U15256 ( .IN1(\mem2[125][19] ), .IN2(n1117), .S(n8097), .Q(n11415)
         );
  MUX21X1 U15257 ( .IN1(\mem2[125][18] ), .IN2(n1095), .S(n8097), .Q(n11414)
         );
  MUX21X1 U15258 ( .IN1(\mem2[125][17] ), .IN2(n1073), .S(n8097), .Q(n11413)
         );
  MUX21X1 U15259 ( .IN1(\mem2[125][16] ), .IN2(n1051), .S(n8097), .Q(n11412)
         );
  AND2X1 U15260 ( .IN1(n8095), .IN2(n7104), .Q(n8097) );
  MUX21X1 U15261 ( .IN1(\mem2[124][23] ), .IN2(n1205), .S(n8098), .Q(n11411)
         );
  MUX21X1 U15262 ( .IN1(\mem2[124][22] ), .IN2(n1183), .S(n8098), .Q(n11410)
         );
  MUX21X1 U15263 ( .IN1(\mem2[124][21] ), .IN2(n1161), .S(n8098), .Q(n11409)
         );
  MUX21X1 U15264 ( .IN1(\mem2[124][20] ), .IN2(n1139), .S(n8098), .Q(n11408)
         );
  MUX21X1 U15265 ( .IN1(\mem2[124][19] ), .IN2(n1117), .S(n8098), .Q(n11407)
         );
  MUX21X1 U15266 ( .IN1(\mem2[124][18] ), .IN2(n1095), .S(n8098), .Q(n11406)
         );
  MUX21X1 U15267 ( .IN1(\mem2[124][17] ), .IN2(n1073), .S(n8098), .Q(n11405)
         );
  MUX21X1 U15268 ( .IN1(\mem2[124][16] ), .IN2(n1051), .S(n8098), .Q(n11404)
         );
  AND2X1 U15269 ( .IN1(n8095), .IN2(n7106), .Q(n8098) );
  MUX21X1 U15270 ( .IN1(\mem2[123][23] ), .IN2(n1206), .S(n8099), .Q(n11403)
         );
  MUX21X1 U15271 ( .IN1(\mem2[123][22] ), .IN2(n1184), .S(n8099), .Q(n11402)
         );
  MUX21X1 U15272 ( .IN1(\mem2[123][21] ), .IN2(n1162), .S(n8099), .Q(n11401)
         );
  MUX21X1 U15273 ( .IN1(\mem2[123][20] ), .IN2(n1140), .S(n8099), .Q(n11400)
         );
  MUX21X1 U15274 ( .IN1(\mem2[123][19] ), .IN2(n1118), .S(n8099), .Q(n11399)
         );
  MUX21X1 U15275 ( .IN1(\mem2[123][18] ), .IN2(n1096), .S(n8099), .Q(n11398)
         );
  MUX21X1 U15276 ( .IN1(\mem2[123][17] ), .IN2(n1074), .S(n8099), .Q(n11397)
         );
  MUX21X1 U15277 ( .IN1(\mem2[123][16] ), .IN2(n1052), .S(n8099), .Q(n11396)
         );
  AND2X1 U15278 ( .IN1(n8095), .IN2(n7108), .Q(n8099) );
  MUX21X1 U15279 ( .IN1(\mem2[122][23] ), .IN2(n1206), .S(n8100), .Q(n11395)
         );
  MUX21X1 U15280 ( .IN1(\mem2[122][22] ), .IN2(n1184), .S(n8100), .Q(n11394)
         );
  MUX21X1 U15281 ( .IN1(\mem2[122][21] ), .IN2(n1162), .S(n8100), .Q(n11393)
         );
  MUX21X1 U15282 ( .IN1(\mem2[122][20] ), .IN2(n1140), .S(n8100), .Q(n11392)
         );
  MUX21X1 U15283 ( .IN1(\mem2[122][19] ), .IN2(n1118), .S(n8100), .Q(n11391)
         );
  MUX21X1 U15284 ( .IN1(\mem2[122][18] ), .IN2(n1096), .S(n8100), .Q(n11390)
         );
  MUX21X1 U15285 ( .IN1(\mem2[122][17] ), .IN2(n1074), .S(n8100), .Q(n11389)
         );
  MUX21X1 U15286 ( .IN1(\mem2[122][16] ), .IN2(n1052), .S(n8100), .Q(n11388)
         );
  AND2X1 U15287 ( .IN1(n8095), .IN2(n7110), .Q(n8100) );
  MUX21X1 U15288 ( .IN1(\mem2[121][23] ), .IN2(n1206), .S(n8101), .Q(n11387)
         );
  MUX21X1 U15289 ( .IN1(\mem2[121][22] ), .IN2(n1184), .S(n8101), .Q(n11386)
         );
  MUX21X1 U15290 ( .IN1(\mem2[121][21] ), .IN2(n1162), .S(n8101), .Q(n11385)
         );
  MUX21X1 U15291 ( .IN1(\mem2[121][20] ), .IN2(n1140), .S(n8101), .Q(n11384)
         );
  MUX21X1 U15292 ( .IN1(\mem2[121][19] ), .IN2(n1118), .S(n8101), .Q(n11383)
         );
  MUX21X1 U15293 ( .IN1(\mem2[121][18] ), .IN2(n1096), .S(n8101), .Q(n11382)
         );
  MUX21X1 U15294 ( .IN1(\mem2[121][17] ), .IN2(n1074), .S(n8101), .Q(n11381)
         );
  MUX21X1 U15295 ( .IN1(\mem2[121][16] ), .IN2(n1052), .S(n8101), .Q(n11380)
         );
  AND2X1 U15296 ( .IN1(n8095), .IN2(n7112), .Q(n8101) );
  MUX21X1 U15297 ( .IN1(\mem2[120][23] ), .IN2(n1206), .S(n8102), .Q(n11379)
         );
  MUX21X1 U15298 ( .IN1(\mem2[120][22] ), .IN2(n1184), .S(n8102), .Q(n11378)
         );
  MUX21X1 U15299 ( .IN1(\mem2[120][21] ), .IN2(n1162), .S(n8102), .Q(n11377)
         );
  MUX21X1 U15300 ( .IN1(\mem2[120][20] ), .IN2(n1140), .S(n8102), .Q(n11376)
         );
  MUX21X1 U15301 ( .IN1(\mem2[120][19] ), .IN2(n1118), .S(n8102), .Q(n11375)
         );
  MUX21X1 U15302 ( .IN1(\mem2[120][18] ), .IN2(n1096), .S(n8102), .Q(n11374)
         );
  MUX21X1 U15303 ( .IN1(\mem2[120][17] ), .IN2(n1074), .S(n8102), .Q(n11373)
         );
  MUX21X1 U15304 ( .IN1(\mem2[120][16] ), .IN2(n1052), .S(n8102), .Q(n11372)
         );
  AND2X1 U15305 ( .IN1(n8095), .IN2(n7114), .Q(n8102) );
  MUX21X1 U15306 ( .IN1(\mem2[119][23] ), .IN2(n1206), .S(n8103), .Q(n11371)
         );
  MUX21X1 U15307 ( .IN1(\mem2[119][22] ), .IN2(n1184), .S(n8103), .Q(n11370)
         );
  MUX21X1 U15308 ( .IN1(\mem2[119][21] ), .IN2(n1162), .S(n8103), .Q(n11369)
         );
  MUX21X1 U15309 ( .IN1(\mem2[119][20] ), .IN2(n1140), .S(n8103), .Q(n11368)
         );
  MUX21X1 U15310 ( .IN1(\mem2[119][19] ), .IN2(n1118), .S(n8103), .Q(n11367)
         );
  MUX21X1 U15311 ( .IN1(\mem2[119][18] ), .IN2(n1096), .S(n8103), .Q(n11366)
         );
  MUX21X1 U15312 ( .IN1(\mem2[119][17] ), .IN2(n1074), .S(n8103), .Q(n11365)
         );
  MUX21X1 U15313 ( .IN1(\mem2[119][16] ), .IN2(n1052), .S(n8103), .Q(n11364)
         );
  AND2X1 U15314 ( .IN1(n8095), .IN2(n7116), .Q(n8103) );
  MUX21X1 U15315 ( .IN1(\mem2[118][23] ), .IN2(n1206), .S(n8104), .Q(n11363)
         );
  MUX21X1 U15316 ( .IN1(\mem2[118][22] ), .IN2(n1184), .S(n8104), .Q(n11362)
         );
  MUX21X1 U15317 ( .IN1(\mem2[118][21] ), .IN2(n1162), .S(n8104), .Q(n11361)
         );
  MUX21X1 U15318 ( .IN1(\mem2[118][20] ), .IN2(n1140), .S(n8104), .Q(n11360)
         );
  MUX21X1 U15319 ( .IN1(\mem2[118][19] ), .IN2(n1118), .S(n8104), .Q(n11359)
         );
  MUX21X1 U15320 ( .IN1(\mem2[118][18] ), .IN2(n1096), .S(n8104), .Q(n11358)
         );
  MUX21X1 U15321 ( .IN1(\mem2[118][17] ), .IN2(n1074), .S(n8104), .Q(n11357)
         );
  MUX21X1 U15322 ( .IN1(\mem2[118][16] ), .IN2(n1052), .S(n8104), .Q(n11356)
         );
  AND2X1 U15323 ( .IN1(n8095), .IN2(n7118), .Q(n8104) );
  MUX21X1 U15324 ( .IN1(\mem2[117][23] ), .IN2(n1206), .S(n8105), .Q(n11355)
         );
  MUX21X1 U15325 ( .IN1(\mem2[117][22] ), .IN2(n1184), .S(n8105), .Q(n11354)
         );
  MUX21X1 U15326 ( .IN1(\mem2[117][21] ), .IN2(n1162), .S(n8105), .Q(n11353)
         );
  MUX21X1 U15327 ( .IN1(\mem2[117][20] ), .IN2(n1140), .S(n8105), .Q(n11352)
         );
  MUX21X1 U15328 ( .IN1(\mem2[117][19] ), .IN2(n1118), .S(n8105), .Q(n11351)
         );
  MUX21X1 U15329 ( .IN1(\mem2[117][18] ), .IN2(n1096), .S(n8105), .Q(n11350)
         );
  MUX21X1 U15330 ( .IN1(\mem2[117][17] ), .IN2(n1074), .S(n8105), .Q(n11349)
         );
  MUX21X1 U15331 ( .IN1(\mem2[117][16] ), .IN2(n1052), .S(n8105), .Q(n11348)
         );
  AND2X1 U15332 ( .IN1(n8095), .IN2(n7120), .Q(n8105) );
  MUX21X1 U15333 ( .IN1(\mem2[116][23] ), .IN2(n1206), .S(n8106), .Q(n11347)
         );
  MUX21X1 U15334 ( .IN1(\mem2[116][22] ), .IN2(n1184), .S(n8106), .Q(n11346)
         );
  MUX21X1 U15335 ( .IN1(\mem2[116][21] ), .IN2(n1162), .S(n8106), .Q(n11345)
         );
  MUX21X1 U15336 ( .IN1(\mem2[116][20] ), .IN2(n1140), .S(n8106), .Q(n11344)
         );
  MUX21X1 U15337 ( .IN1(\mem2[116][19] ), .IN2(n1118), .S(n8106), .Q(n11343)
         );
  MUX21X1 U15338 ( .IN1(\mem2[116][18] ), .IN2(n1096), .S(n8106), .Q(n11342)
         );
  MUX21X1 U15339 ( .IN1(\mem2[116][17] ), .IN2(n1074), .S(n8106), .Q(n11341)
         );
  MUX21X1 U15340 ( .IN1(\mem2[116][16] ), .IN2(n1052), .S(n8106), .Q(n11340)
         );
  AND2X1 U15341 ( .IN1(n8095), .IN2(n7122), .Q(n8106) );
  MUX21X1 U15342 ( .IN1(\mem2[115][23] ), .IN2(n1206), .S(n8107), .Q(n11339)
         );
  MUX21X1 U15343 ( .IN1(\mem2[115][22] ), .IN2(n1184), .S(n8107), .Q(n11338)
         );
  MUX21X1 U15344 ( .IN1(\mem2[115][21] ), .IN2(n1162), .S(n8107), .Q(n11337)
         );
  MUX21X1 U15345 ( .IN1(\mem2[115][20] ), .IN2(n1140), .S(n8107), .Q(n11336)
         );
  MUX21X1 U15346 ( .IN1(\mem2[115][19] ), .IN2(n1118), .S(n8107), .Q(n11335)
         );
  MUX21X1 U15347 ( .IN1(\mem2[115][18] ), .IN2(n1096), .S(n8107), .Q(n11334)
         );
  MUX21X1 U15348 ( .IN1(\mem2[115][17] ), .IN2(n1074), .S(n8107), .Q(n11333)
         );
  MUX21X1 U15349 ( .IN1(\mem2[115][16] ), .IN2(n1052), .S(n8107), .Q(n11332)
         );
  AND2X1 U15350 ( .IN1(n8095), .IN2(n7124), .Q(n8107) );
  MUX21X1 U15351 ( .IN1(\mem2[114][23] ), .IN2(n1206), .S(n8108), .Q(n11331)
         );
  MUX21X1 U15352 ( .IN1(\mem2[114][22] ), .IN2(n1184), .S(n8108), .Q(n11330)
         );
  MUX21X1 U15353 ( .IN1(\mem2[114][21] ), .IN2(n1162), .S(n8108), .Q(n11329)
         );
  MUX21X1 U15354 ( .IN1(\mem2[114][20] ), .IN2(n1140), .S(n8108), .Q(n11328)
         );
  MUX21X1 U15355 ( .IN1(\mem2[114][19] ), .IN2(n1118), .S(n8108), .Q(n11327)
         );
  MUX21X1 U15356 ( .IN1(\mem2[114][18] ), .IN2(n1096), .S(n8108), .Q(n11326)
         );
  MUX21X1 U15357 ( .IN1(\mem2[114][17] ), .IN2(n1074), .S(n8108), .Q(n11325)
         );
  MUX21X1 U15358 ( .IN1(\mem2[114][16] ), .IN2(n1052), .S(n8108), .Q(n11324)
         );
  AND2X1 U15359 ( .IN1(n8095), .IN2(n7126), .Q(n8108) );
  MUX21X1 U15360 ( .IN1(\mem2[113][23] ), .IN2(n1206), .S(n8109), .Q(n11323)
         );
  MUX21X1 U15361 ( .IN1(\mem2[113][22] ), .IN2(n1184), .S(n8109), .Q(n11322)
         );
  MUX21X1 U15362 ( .IN1(\mem2[113][21] ), .IN2(n1162), .S(n8109), .Q(n11321)
         );
  MUX21X1 U15363 ( .IN1(\mem2[113][20] ), .IN2(n1140), .S(n8109), .Q(n11320)
         );
  MUX21X1 U15364 ( .IN1(\mem2[113][19] ), .IN2(n1118), .S(n8109), .Q(n11319)
         );
  MUX21X1 U15365 ( .IN1(\mem2[113][18] ), .IN2(n1096), .S(n8109), .Q(n11318)
         );
  MUX21X1 U15366 ( .IN1(\mem2[113][17] ), .IN2(n1074), .S(n8109), .Q(n11317)
         );
  MUX21X1 U15367 ( .IN1(\mem2[113][16] ), .IN2(n1052), .S(n8109), .Q(n11316)
         );
  AND2X1 U15368 ( .IN1(n8095), .IN2(n7128), .Q(n8109) );
  MUX21X1 U15369 ( .IN1(\mem2[112][23] ), .IN2(n1206), .S(n8110), .Q(n11315)
         );
  MUX21X1 U15370 ( .IN1(\mem2[112][22] ), .IN2(n1184), .S(n8110), .Q(n11314)
         );
  MUX21X1 U15371 ( .IN1(\mem2[112][21] ), .IN2(n1162), .S(n8110), .Q(n11313)
         );
  MUX21X1 U15372 ( .IN1(\mem2[112][20] ), .IN2(n1140), .S(n8110), .Q(n11312)
         );
  MUX21X1 U15373 ( .IN1(\mem2[112][19] ), .IN2(n1118), .S(n8110), .Q(n11311)
         );
  MUX21X1 U15374 ( .IN1(\mem2[112][18] ), .IN2(n1096), .S(n8110), .Q(n11310)
         );
  MUX21X1 U15375 ( .IN1(\mem2[112][17] ), .IN2(n1074), .S(n8110), .Q(n11309)
         );
  MUX21X1 U15376 ( .IN1(\mem2[112][16] ), .IN2(n1052), .S(n8110), .Q(n11308)
         );
  AND2X1 U15377 ( .IN1(n8095), .IN2(n7130), .Q(n8110) );
  AND2X1 U15378 ( .IN1(n7966), .IN2(n7276), .Q(n8095) );
  AND2X1 U15379 ( .IN1(n8111), .IN2(n7968), .Q(n7276) );
  MUX21X1 U15380 ( .IN1(\mem2[111][23] ), .IN2(n1207), .S(n8112), .Q(n11307)
         );
  MUX21X1 U15381 ( .IN1(\mem2[111][22] ), .IN2(n1185), .S(n8112), .Q(n11306)
         );
  MUX21X1 U15382 ( .IN1(\mem2[111][21] ), .IN2(n1163), .S(n8112), .Q(n11305)
         );
  MUX21X1 U15383 ( .IN1(\mem2[111][20] ), .IN2(n1141), .S(n8112), .Q(n11304)
         );
  MUX21X1 U15384 ( .IN1(\mem2[111][19] ), .IN2(n1119), .S(n8112), .Q(n11303)
         );
  MUX21X1 U15385 ( .IN1(\mem2[111][18] ), .IN2(n1097), .S(n8112), .Q(n11302)
         );
  MUX21X1 U15386 ( .IN1(\mem2[111][17] ), .IN2(n1075), .S(n8112), .Q(n11301)
         );
  MUX21X1 U15387 ( .IN1(\mem2[111][16] ), .IN2(n1053), .S(n8112), .Q(n11300)
         );
  AND2X1 U15388 ( .IN1(n8113), .IN2(n7099), .Q(n8112) );
  MUX21X1 U15389 ( .IN1(\mem2[110][23] ), .IN2(n1207), .S(n8114), .Q(n11299)
         );
  MUX21X1 U15390 ( .IN1(\mem2[110][22] ), .IN2(n1185), .S(n8114), .Q(n11298)
         );
  MUX21X1 U15391 ( .IN1(\mem2[110][21] ), .IN2(n1163), .S(n8114), .Q(n11297)
         );
  MUX21X1 U15392 ( .IN1(\mem2[110][20] ), .IN2(n1141), .S(n8114), .Q(n11296)
         );
  MUX21X1 U15393 ( .IN1(\mem2[110][19] ), .IN2(n1119), .S(n8114), .Q(n11295)
         );
  MUX21X1 U15394 ( .IN1(\mem2[110][18] ), .IN2(n1097), .S(n8114), .Q(n11294)
         );
  MUX21X1 U15395 ( .IN1(\mem2[110][17] ), .IN2(n1075), .S(n8114), .Q(n11293)
         );
  MUX21X1 U15396 ( .IN1(\mem2[110][16] ), .IN2(n1053), .S(n8114), .Q(n11292)
         );
  AND2X1 U15397 ( .IN1(n8113), .IN2(n7102), .Q(n8114) );
  MUX21X1 U15398 ( .IN1(\mem2[109][23] ), .IN2(n1207), .S(n8115), .Q(n11291)
         );
  MUX21X1 U15399 ( .IN1(\mem2[109][22] ), .IN2(n1185), .S(n8115), .Q(n11290)
         );
  MUX21X1 U15400 ( .IN1(\mem2[109][21] ), .IN2(n1163), .S(n8115), .Q(n11289)
         );
  MUX21X1 U15401 ( .IN1(\mem2[109][20] ), .IN2(n1141), .S(n8115), .Q(n11288)
         );
  MUX21X1 U15402 ( .IN1(\mem2[109][19] ), .IN2(n1119), .S(n8115), .Q(n11287)
         );
  MUX21X1 U15403 ( .IN1(\mem2[109][18] ), .IN2(n1097), .S(n8115), .Q(n11286)
         );
  MUX21X1 U15404 ( .IN1(\mem2[109][17] ), .IN2(n1075), .S(n8115), .Q(n11285)
         );
  MUX21X1 U15405 ( .IN1(\mem2[109][16] ), .IN2(n1053), .S(n8115), .Q(n11284)
         );
  AND2X1 U15406 ( .IN1(n8113), .IN2(n7104), .Q(n8115) );
  MUX21X1 U15407 ( .IN1(\mem2[108][23] ), .IN2(n1207), .S(n8116), .Q(n11283)
         );
  MUX21X1 U15408 ( .IN1(\mem2[108][22] ), .IN2(n1185), .S(n8116), .Q(n11282)
         );
  MUX21X1 U15409 ( .IN1(\mem2[108][21] ), .IN2(n1163), .S(n8116), .Q(n11281)
         );
  MUX21X1 U15410 ( .IN1(\mem2[108][20] ), .IN2(n1141), .S(n8116), .Q(n11280)
         );
  MUX21X1 U15411 ( .IN1(\mem2[108][19] ), .IN2(n1119), .S(n8116), .Q(n11279)
         );
  MUX21X1 U15412 ( .IN1(\mem2[108][18] ), .IN2(n1097), .S(n8116), .Q(n11278)
         );
  MUX21X1 U15413 ( .IN1(\mem2[108][17] ), .IN2(n1075), .S(n8116), .Q(n11277)
         );
  MUX21X1 U15414 ( .IN1(\mem2[108][16] ), .IN2(n1053), .S(n8116), .Q(n11276)
         );
  AND2X1 U15415 ( .IN1(n8113), .IN2(n7106), .Q(n8116) );
  MUX21X1 U15416 ( .IN1(\mem2[107][23] ), .IN2(n1207), .S(n8117), .Q(n11275)
         );
  MUX21X1 U15417 ( .IN1(\mem2[107][22] ), .IN2(n1185), .S(n8117), .Q(n11274)
         );
  MUX21X1 U15418 ( .IN1(\mem2[107][21] ), .IN2(n1163), .S(n8117), .Q(n11273)
         );
  MUX21X1 U15419 ( .IN1(\mem2[107][20] ), .IN2(n1141), .S(n8117), .Q(n11272)
         );
  MUX21X1 U15420 ( .IN1(\mem2[107][19] ), .IN2(n1119), .S(n8117), .Q(n11271)
         );
  MUX21X1 U15421 ( .IN1(\mem2[107][18] ), .IN2(n1097), .S(n8117), .Q(n11270)
         );
  MUX21X1 U15422 ( .IN1(\mem2[107][17] ), .IN2(n1075), .S(n8117), .Q(n11269)
         );
  MUX21X1 U15423 ( .IN1(\mem2[107][16] ), .IN2(n1053), .S(n8117), .Q(n11268)
         );
  AND2X1 U15424 ( .IN1(n8113), .IN2(n7108), .Q(n8117) );
  MUX21X1 U15425 ( .IN1(\mem2[106][23] ), .IN2(n1207), .S(n8118), .Q(n11267)
         );
  MUX21X1 U15426 ( .IN1(\mem2[106][22] ), .IN2(n1185), .S(n8118), .Q(n11266)
         );
  MUX21X1 U15427 ( .IN1(\mem2[106][21] ), .IN2(n1163), .S(n8118), .Q(n11265)
         );
  MUX21X1 U15428 ( .IN1(\mem2[106][20] ), .IN2(n1141), .S(n8118), .Q(n11264)
         );
  MUX21X1 U15429 ( .IN1(\mem2[106][19] ), .IN2(n1119), .S(n8118), .Q(n11263)
         );
  MUX21X1 U15430 ( .IN1(\mem2[106][18] ), .IN2(n1097), .S(n8118), .Q(n11262)
         );
  MUX21X1 U15431 ( .IN1(\mem2[106][17] ), .IN2(n1075), .S(n8118), .Q(n11261)
         );
  MUX21X1 U15432 ( .IN1(\mem2[106][16] ), .IN2(n1053), .S(n8118), .Q(n11260)
         );
  AND2X1 U15433 ( .IN1(n8113), .IN2(n7110), .Q(n8118) );
  MUX21X1 U15434 ( .IN1(\mem2[105][23] ), .IN2(n1207), .S(n8119), .Q(n11259)
         );
  MUX21X1 U15435 ( .IN1(\mem2[105][22] ), .IN2(n1185), .S(n8119), .Q(n11258)
         );
  MUX21X1 U15436 ( .IN1(\mem2[105][21] ), .IN2(n1163), .S(n8119), .Q(n11257)
         );
  MUX21X1 U15437 ( .IN1(\mem2[105][20] ), .IN2(n1141), .S(n8119), .Q(n11256)
         );
  MUX21X1 U15438 ( .IN1(\mem2[105][19] ), .IN2(n1119), .S(n8119), .Q(n11255)
         );
  MUX21X1 U15439 ( .IN1(\mem2[105][18] ), .IN2(n1097), .S(n8119), .Q(n11254)
         );
  MUX21X1 U15440 ( .IN1(\mem2[105][17] ), .IN2(n1075), .S(n8119), .Q(n11253)
         );
  MUX21X1 U15441 ( .IN1(\mem2[105][16] ), .IN2(n1053), .S(n8119), .Q(n11252)
         );
  AND2X1 U15442 ( .IN1(n8113), .IN2(n7112), .Q(n8119) );
  MUX21X1 U15443 ( .IN1(\mem2[104][23] ), .IN2(n1207), .S(n8120), .Q(n11251)
         );
  MUX21X1 U15444 ( .IN1(\mem2[104][22] ), .IN2(n1185), .S(n8120), .Q(n11250)
         );
  MUX21X1 U15445 ( .IN1(\mem2[104][21] ), .IN2(n1163), .S(n8120), .Q(n11249)
         );
  MUX21X1 U15446 ( .IN1(\mem2[104][20] ), .IN2(n1141), .S(n8120), .Q(n11248)
         );
  MUX21X1 U15447 ( .IN1(\mem2[104][19] ), .IN2(n1119), .S(n8120), .Q(n11247)
         );
  MUX21X1 U15448 ( .IN1(\mem2[104][18] ), .IN2(n1097), .S(n8120), .Q(n11246)
         );
  MUX21X1 U15449 ( .IN1(\mem2[104][17] ), .IN2(n1075), .S(n8120), .Q(n11245)
         );
  MUX21X1 U15450 ( .IN1(\mem2[104][16] ), .IN2(n1053), .S(n8120), .Q(n11244)
         );
  AND2X1 U15451 ( .IN1(n8113), .IN2(n7114), .Q(n8120) );
  MUX21X1 U15452 ( .IN1(\mem2[103][23] ), .IN2(n1207), .S(n8121), .Q(n11243)
         );
  MUX21X1 U15453 ( .IN1(\mem2[103][22] ), .IN2(n1185), .S(n8121), .Q(n11242)
         );
  MUX21X1 U15454 ( .IN1(\mem2[103][21] ), .IN2(n1163), .S(n8121), .Q(n11241)
         );
  MUX21X1 U15455 ( .IN1(\mem2[103][20] ), .IN2(n1141), .S(n8121), .Q(n11240)
         );
  MUX21X1 U15456 ( .IN1(\mem2[103][19] ), .IN2(n1119), .S(n8121), .Q(n11239)
         );
  MUX21X1 U15457 ( .IN1(\mem2[103][18] ), .IN2(n1097), .S(n8121), .Q(n11238)
         );
  MUX21X1 U15458 ( .IN1(\mem2[103][17] ), .IN2(n1075), .S(n8121), .Q(n11237)
         );
  MUX21X1 U15459 ( .IN1(\mem2[103][16] ), .IN2(n1053), .S(n8121), .Q(n11236)
         );
  AND2X1 U15460 ( .IN1(n8113), .IN2(n7116), .Q(n8121) );
  MUX21X1 U15461 ( .IN1(\mem2[102][23] ), .IN2(n1207), .S(n8122), .Q(n11235)
         );
  MUX21X1 U15462 ( .IN1(\mem2[102][22] ), .IN2(n1185), .S(n8122), .Q(n11234)
         );
  MUX21X1 U15463 ( .IN1(\mem2[102][21] ), .IN2(n1163), .S(n8122), .Q(n11233)
         );
  MUX21X1 U15464 ( .IN1(\mem2[102][20] ), .IN2(n1141), .S(n8122), .Q(n11232)
         );
  MUX21X1 U15465 ( .IN1(\mem2[102][19] ), .IN2(n1119), .S(n8122), .Q(n11231)
         );
  MUX21X1 U15466 ( .IN1(\mem2[102][18] ), .IN2(n1097), .S(n8122), .Q(n11230)
         );
  MUX21X1 U15467 ( .IN1(\mem2[102][17] ), .IN2(n1075), .S(n8122), .Q(n11229)
         );
  MUX21X1 U15468 ( .IN1(\mem2[102][16] ), .IN2(n1053), .S(n8122), .Q(n11228)
         );
  AND2X1 U15469 ( .IN1(n8113), .IN2(n7118), .Q(n8122) );
  MUX21X1 U15470 ( .IN1(\mem2[101][23] ), .IN2(n1207), .S(n8123), .Q(n11227)
         );
  MUX21X1 U15471 ( .IN1(\mem2[101][22] ), .IN2(n1185), .S(n8123), .Q(n11226)
         );
  MUX21X1 U15472 ( .IN1(\mem2[101][21] ), .IN2(n1163), .S(n8123), .Q(n11225)
         );
  MUX21X1 U15473 ( .IN1(\mem2[101][20] ), .IN2(n1141), .S(n8123), .Q(n11224)
         );
  MUX21X1 U15474 ( .IN1(\mem2[101][19] ), .IN2(n1119), .S(n8123), .Q(n11223)
         );
  MUX21X1 U15475 ( .IN1(\mem2[101][18] ), .IN2(n1097), .S(n8123), .Q(n11222)
         );
  MUX21X1 U15476 ( .IN1(\mem2[101][17] ), .IN2(n1075), .S(n8123), .Q(n11221)
         );
  MUX21X1 U15477 ( .IN1(\mem2[101][16] ), .IN2(n1053), .S(n8123), .Q(n11220)
         );
  AND2X1 U15478 ( .IN1(n8113), .IN2(n7120), .Q(n8123) );
  MUX21X1 U15479 ( .IN1(\mem2[100][23] ), .IN2(n1207), .S(n8124), .Q(n11219)
         );
  MUX21X1 U15480 ( .IN1(\mem2[100][22] ), .IN2(n1185), .S(n8124), .Q(n11218)
         );
  MUX21X1 U15481 ( .IN1(\mem2[100][21] ), .IN2(n1163), .S(n8124), .Q(n11217)
         );
  MUX21X1 U15482 ( .IN1(\mem2[100][20] ), .IN2(n1141), .S(n8124), .Q(n11216)
         );
  MUX21X1 U15483 ( .IN1(\mem2[100][19] ), .IN2(n1119), .S(n8124), .Q(n11215)
         );
  MUX21X1 U15484 ( .IN1(\mem2[100][18] ), .IN2(n1097), .S(n8124), .Q(n11214)
         );
  MUX21X1 U15485 ( .IN1(\mem2[100][17] ), .IN2(n1075), .S(n8124), .Q(n11213)
         );
  MUX21X1 U15486 ( .IN1(\mem2[100][16] ), .IN2(n1053), .S(n8124), .Q(n11212)
         );
  AND2X1 U15487 ( .IN1(n8113), .IN2(n7122), .Q(n8124) );
  MUX21X1 U15488 ( .IN1(\mem2[99][23] ), .IN2(n1208), .S(n8125), .Q(n11211) );
  MUX21X1 U15489 ( .IN1(\mem2[99][22] ), .IN2(n1186), .S(n8125), .Q(n11210) );
  MUX21X1 U15490 ( .IN1(\mem2[99][21] ), .IN2(n1164), .S(n8125), .Q(n11209) );
  MUX21X1 U15491 ( .IN1(\mem2[99][20] ), .IN2(n1142), .S(n8125), .Q(n11208) );
  MUX21X1 U15492 ( .IN1(\mem2[99][19] ), .IN2(n1120), .S(n8125), .Q(n11207) );
  MUX21X1 U15493 ( .IN1(\mem2[99][18] ), .IN2(n1098), .S(n8125), .Q(n11206) );
  MUX21X1 U15494 ( .IN1(\mem2[99][17] ), .IN2(n1076), .S(n8125), .Q(n11205) );
  MUX21X1 U15495 ( .IN1(\mem2[99][16] ), .IN2(n1054), .S(n8125), .Q(n11204) );
  AND2X1 U15496 ( .IN1(n8113), .IN2(n7124), .Q(n8125) );
  MUX21X1 U15497 ( .IN1(\mem2[98][23] ), .IN2(n1208), .S(n8126), .Q(n11203) );
  MUX21X1 U15498 ( .IN1(\mem2[98][22] ), .IN2(n1186), .S(n8126), .Q(n11202) );
  MUX21X1 U15499 ( .IN1(\mem2[98][21] ), .IN2(n1164), .S(n8126), .Q(n11201) );
  MUX21X1 U15500 ( .IN1(\mem2[98][20] ), .IN2(n1142), .S(n8126), .Q(n11200) );
  MUX21X1 U15501 ( .IN1(\mem2[98][19] ), .IN2(n1120), .S(n8126), .Q(n11199) );
  MUX21X1 U15502 ( .IN1(\mem2[98][18] ), .IN2(n1098), .S(n8126), .Q(n11198) );
  MUX21X1 U15503 ( .IN1(\mem2[98][17] ), .IN2(n1076), .S(n8126), .Q(n11197) );
  MUX21X1 U15504 ( .IN1(\mem2[98][16] ), .IN2(n1054), .S(n8126), .Q(n11196) );
  AND2X1 U15505 ( .IN1(n8113), .IN2(n7126), .Q(n8126) );
  MUX21X1 U15506 ( .IN1(\mem2[97][23] ), .IN2(n1208), .S(n8127), .Q(n11195) );
  MUX21X1 U15507 ( .IN1(\mem2[97][22] ), .IN2(n1186), .S(n8127), .Q(n11194) );
  MUX21X1 U15508 ( .IN1(\mem2[97][21] ), .IN2(n1164), .S(n8127), .Q(n11193) );
  MUX21X1 U15509 ( .IN1(\mem2[97][20] ), .IN2(n1142), .S(n8127), .Q(n11192) );
  MUX21X1 U15510 ( .IN1(\mem2[97][19] ), .IN2(n1120), .S(n8127), .Q(n11191) );
  MUX21X1 U15511 ( .IN1(\mem2[97][18] ), .IN2(n1098), .S(n8127), .Q(n11190) );
  MUX21X1 U15512 ( .IN1(\mem2[97][17] ), .IN2(n1076), .S(n8127), .Q(n11189) );
  MUX21X1 U15513 ( .IN1(\mem2[97][16] ), .IN2(n1054), .S(n8127), .Q(n11188) );
  AND2X1 U15514 ( .IN1(n8113), .IN2(n7128), .Q(n8127) );
  MUX21X1 U15515 ( .IN1(\mem2[96][23] ), .IN2(n1208), .S(n8128), .Q(n11187) );
  MUX21X1 U15516 ( .IN1(\mem2[96][22] ), .IN2(n1186), .S(n8128), .Q(n11186) );
  MUX21X1 U15517 ( .IN1(\mem2[96][21] ), .IN2(n1164), .S(n8128), .Q(n11185) );
  MUX21X1 U15518 ( .IN1(\mem2[96][20] ), .IN2(n1142), .S(n8128), .Q(n11184) );
  MUX21X1 U15519 ( .IN1(\mem2[96][19] ), .IN2(n1120), .S(n8128), .Q(n11183) );
  MUX21X1 U15520 ( .IN1(\mem2[96][18] ), .IN2(n1098), .S(n8128), .Q(n11182) );
  MUX21X1 U15521 ( .IN1(\mem2[96][17] ), .IN2(n1076), .S(n8128), .Q(n11181) );
  MUX21X1 U15522 ( .IN1(\mem2[96][16] ), .IN2(n1054), .S(n8128), .Q(n11180) );
  AND2X1 U15523 ( .IN1(n8113), .IN2(n7130), .Q(n8128) );
  AND2X1 U15524 ( .IN1(n7966), .IN2(n7294), .Q(n8113) );
  AND2X1 U15525 ( .IN1(n8111), .IN2(n7986), .Q(n7294) );
  MUX21X1 U15526 ( .IN1(\mem2[95][23] ), .IN2(n1208), .S(n8129), .Q(n11179) );
  MUX21X1 U15527 ( .IN1(\mem2[95][22] ), .IN2(n1186), .S(n8129), .Q(n11178) );
  MUX21X1 U15528 ( .IN1(\mem2[95][21] ), .IN2(n1164), .S(n8129), .Q(n11177) );
  MUX21X1 U15529 ( .IN1(\mem2[95][20] ), .IN2(n1142), .S(n8129), .Q(n11176) );
  MUX21X1 U15530 ( .IN1(\mem2[95][19] ), .IN2(n1120), .S(n8129), .Q(n11175) );
  MUX21X1 U15531 ( .IN1(\mem2[95][18] ), .IN2(n1098), .S(n8129), .Q(n11174) );
  MUX21X1 U15532 ( .IN1(\mem2[95][17] ), .IN2(n1076), .S(n8129), .Q(n11173) );
  MUX21X1 U15533 ( .IN1(\mem2[95][16] ), .IN2(n1054), .S(n8129), .Q(n11172) );
  AND2X1 U15534 ( .IN1(n8130), .IN2(n7099), .Q(n8129) );
  MUX21X1 U15535 ( .IN1(\mem2[94][23] ), .IN2(n1208), .S(n8131), .Q(n11171) );
  MUX21X1 U15536 ( .IN1(\mem2[94][22] ), .IN2(n1186), .S(n8131), .Q(n11170) );
  MUX21X1 U15537 ( .IN1(\mem2[94][21] ), .IN2(n1164), .S(n8131), .Q(n11169) );
  MUX21X1 U15538 ( .IN1(\mem2[94][20] ), .IN2(n1142), .S(n8131), .Q(n11168) );
  MUX21X1 U15539 ( .IN1(\mem2[94][19] ), .IN2(n1120), .S(n8131), .Q(n11167) );
  MUX21X1 U15540 ( .IN1(\mem2[94][18] ), .IN2(n1098), .S(n8131), .Q(n11166) );
  MUX21X1 U15541 ( .IN1(\mem2[94][17] ), .IN2(n1076), .S(n8131), .Q(n11165) );
  MUX21X1 U15542 ( .IN1(\mem2[94][16] ), .IN2(n1054), .S(n8131), .Q(n11164) );
  AND2X1 U15543 ( .IN1(n8130), .IN2(n7102), .Q(n8131) );
  MUX21X1 U15544 ( .IN1(\mem2[93][23] ), .IN2(n1208), .S(n8132), .Q(n11163) );
  MUX21X1 U15545 ( .IN1(\mem2[93][22] ), .IN2(n1186), .S(n8132), .Q(n11162) );
  MUX21X1 U15546 ( .IN1(\mem2[93][21] ), .IN2(n1164), .S(n8132), .Q(n11161) );
  MUX21X1 U15547 ( .IN1(\mem2[93][20] ), .IN2(n1142), .S(n8132), .Q(n11160) );
  MUX21X1 U15548 ( .IN1(\mem2[93][19] ), .IN2(n1120), .S(n8132), .Q(n11159) );
  MUX21X1 U15549 ( .IN1(\mem2[93][18] ), .IN2(n1098), .S(n8132), .Q(n11158) );
  MUX21X1 U15550 ( .IN1(\mem2[93][17] ), .IN2(n1076), .S(n8132), .Q(n11157) );
  MUX21X1 U15551 ( .IN1(\mem2[93][16] ), .IN2(n1054), .S(n8132), .Q(n11156) );
  AND2X1 U15552 ( .IN1(n8130), .IN2(n7104), .Q(n8132) );
  MUX21X1 U15553 ( .IN1(\mem2[92][23] ), .IN2(n1208), .S(n8133), .Q(n11155) );
  MUX21X1 U15554 ( .IN1(\mem2[92][22] ), .IN2(n1186), .S(n8133), .Q(n11154) );
  MUX21X1 U15555 ( .IN1(\mem2[92][21] ), .IN2(n1164), .S(n8133), .Q(n11153) );
  MUX21X1 U15556 ( .IN1(\mem2[92][20] ), .IN2(n1142), .S(n8133), .Q(n11152) );
  MUX21X1 U15557 ( .IN1(\mem2[92][19] ), .IN2(n1120), .S(n8133), .Q(n11151) );
  MUX21X1 U15558 ( .IN1(\mem2[92][18] ), .IN2(n1098), .S(n8133), .Q(n11150) );
  MUX21X1 U15559 ( .IN1(\mem2[92][17] ), .IN2(n1076), .S(n8133), .Q(n11149) );
  MUX21X1 U15560 ( .IN1(\mem2[92][16] ), .IN2(n1054), .S(n8133), .Q(n11148) );
  AND2X1 U15561 ( .IN1(n8130), .IN2(n7106), .Q(n8133) );
  MUX21X1 U15562 ( .IN1(\mem2[91][23] ), .IN2(n1208), .S(n8134), .Q(n11147) );
  MUX21X1 U15563 ( .IN1(\mem2[91][22] ), .IN2(n1186), .S(n8134), .Q(n11146) );
  MUX21X1 U15564 ( .IN1(\mem2[91][21] ), .IN2(n1164), .S(n8134), .Q(n11145) );
  MUX21X1 U15565 ( .IN1(\mem2[91][20] ), .IN2(n1142), .S(n8134), .Q(n11144) );
  MUX21X1 U15566 ( .IN1(\mem2[91][19] ), .IN2(n1120), .S(n8134), .Q(n11143) );
  MUX21X1 U15567 ( .IN1(\mem2[91][18] ), .IN2(n1098), .S(n8134), .Q(n11142) );
  MUX21X1 U15568 ( .IN1(\mem2[91][17] ), .IN2(n1076), .S(n8134), .Q(n11141) );
  MUX21X1 U15569 ( .IN1(\mem2[91][16] ), .IN2(n1054), .S(n8134), .Q(n11140) );
  AND2X1 U15570 ( .IN1(n8130), .IN2(n7108), .Q(n8134) );
  MUX21X1 U15571 ( .IN1(\mem2[90][23] ), .IN2(n1208), .S(n8135), .Q(n11139) );
  MUX21X1 U15572 ( .IN1(\mem2[90][22] ), .IN2(n1186), .S(n8135), .Q(n11138) );
  MUX21X1 U15573 ( .IN1(\mem2[90][21] ), .IN2(n1164), .S(n8135), .Q(n11137) );
  MUX21X1 U15574 ( .IN1(\mem2[90][20] ), .IN2(n1142), .S(n8135), .Q(n11136) );
  MUX21X1 U15575 ( .IN1(\mem2[90][19] ), .IN2(n1120), .S(n8135), .Q(n11135) );
  MUX21X1 U15576 ( .IN1(\mem2[90][18] ), .IN2(n1098), .S(n8135), .Q(n11134) );
  MUX21X1 U15577 ( .IN1(\mem2[90][17] ), .IN2(n1076), .S(n8135), .Q(n11133) );
  MUX21X1 U15578 ( .IN1(\mem2[90][16] ), .IN2(n1054), .S(n8135), .Q(n11132) );
  AND2X1 U15579 ( .IN1(n8130), .IN2(n7110), .Q(n8135) );
  MUX21X1 U15580 ( .IN1(\mem2[89][23] ), .IN2(n1208), .S(n8136), .Q(n11131) );
  MUX21X1 U15581 ( .IN1(\mem2[89][22] ), .IN2(n1186), .S(n8136), .Q(n11130) );
  MUX21X1 U15582 ( .IN1(\mem2[89][21] ), .IN2(n1164), .S(n8136), .Q(n11129) );
  MUX21X1 U15583 ( .IN1(\mem2[89][20] ), .IN2(n1142), .S(n8136), .Q(n11128) );
  MUX21X1 U15584 ( .IN1(\mem2[89][19] ), .IN2(n1120), .S(n8136), .Q(n11127) );
  MUX21X1 U15585 ( .IN1(\mem2[89][18] ), .IN2(n1098), .S(n8136), .Q(n11126) );
  MUX21X1 U15586 ( .IN1(\mem2[89][17] ), .IN2(n1076), .S(n8136), .Q(n11125) );
  MUX21X1 U15587 ( .IN1(\mem2[89][16] ), .IN2(n1054), .S(n8136), .Q(n11124) );
  AND2X1 U15588 ( .IN1(n8130), .IN2(n7112), .Q(n8136) );
  MUX21X1 U15589 ( .IN1(\mem2[88][23] ), .IN2(n1208), .S(n8137), .Q(n11123) );
  MUX21X1 U15590 ( .IN1(\mem2[88][22] ), .IN2(n1186), .S(n8137), .Q(n11122) );
  MUX21X1 U15591 ( .IN1(\mem2[88][21] ), .IN2(n1164), .S(n8137), .Q(n11121) );
  MUX21X1 U15592 ( .IN1(\mem2[88][20] ), .IN2(n1142), .S(n8137), .Q(n11120) );
  MUX21X1 U15593 ( .IN1(\mem2[88][19] ), .IN2(n1120), .S(n8137), .Q(n11119) );
  MUX21X1 U15594 ( .IN1(\mem2[88][18] ), .IN2(n1098), .S(n8137), .Q(n11118) );
  MUX21X1 U15595 ( .IN1(\mem2[88][17] ), .IN2(n1076), .S(n8137), .Q(n11117) );
  MUX21X1 U15596 ( .IN1(\mem2[88][16] ), .IN2(n1054), .S(n8137), .Q(n11116) );
  AND2X1 U15597 ( .IN1(n8130), .IN2(n7114), .Q(n8137) );
  MUX21X1 U15598 ( .IN1(\mem2[87][23] ), .IN2(n1209), .S(n8138), .Q(n11115) );
  MUX21X1 U15599 ( .IN1(\mem2[87][22] ), .IN2(n1187), .S(n8138), .Q(n11114) );
  MUX21X1 U15600 ( .IN1(\mem2[87][21] ), .IN2(n1165), .S(n8138), .Q(n11113) );
  MUX21X1 U15601 ( .IN1(\mem2[87][20] ), .IN2(n1143), .S(n8138), .Q(n11112) );
  MUX21X1 U15602 ( .IN1(\mem2[87][19] ), .IN2(n1121), .S(n8138), .Q(n11111) );
  MUX21X1 U15603 ( .IN1(\mem2[87][18] ), .IN2(n1099), .S(n8138), .Q(n11110) );
  MUX21X1 U15604 ( .IN1(\mem2[87][17] ), .IN2(n1077), .S(n8138), .Q(n11109) );
  MUX21X1 U15605 ( .IN1(\mem2[87][16] ), .IN2(n1055), .S(n8138), .Q(n11108) );
  AND2X1 U15606 ( .IN1(n8130), .IN2(n7116), .Q(n8138) );
  MUX21X1 U15607 ( .IN1(\mem2[86][23] ), .IN2(n1209), .S(n8139), .Q(n11107) );
  MUX21X1 U15608 ( .IN1(\mem2[86][22] ), .IN2(n1187), .S(n8139), .Q(n11106) );
  MUX21X1 U15609 ( .IN1(\mem2[86][21] ), .IN2(n1165), .S(n8139), .Q(n11105) );
  MUX21X1 U15610 ( .IN1(\mem2[86][20] ), .IN2(n1143), .S(n8139), .Q(n11104) );
  MUX21X1 U15611 ( .IN1(\mem2[86][19] ), .IN2(n1121), .S(n8139), .Q(n11103) );
  MUX21X1 U15612 ( .IN1(\mem2[86][18] ), .IN2(n1099), .S(n8139), .Q(n11102) );
  MUX21X1 U15613 ( .IN1(\mem2[86][17] ), .IN2(n1077), .S(n8139), .Q(n11101) );
  MUX21X1 U15614 ( .IN1(\mem2[86][16] ), .IN2(n1055), .S(n8139), .Q(n11100) );
  AND2X1 U15615 ( .IN1(n8130), .IN2(n7118), .Q(n8139) );
  MUX21X1 U15616 ( .IN1(\mem2[85][23] ), .IN2(n1209), .S(n8140), .Q(n11099) );
  MUX21X1 U15617 ( .IN1(\mem2[85][22] ), .IN2(n1187), .S(n8140), .Q(n11098) );
  MUX21X1 U15618 ( .IN1(\mem2[85][21] ), .IN2(n1165), .S(n8140), .Q(n11097) );
  MUX21X1 U15619 ( .IN1(\mem2[85][20] ), .IN2(n1143), .S(n8140), .Q(n11096) );
  MUX21X1 U15620 ( .IN1(\mem2[85][19] ), .IN2(n1121), .S(n8140), .Q(n11095) );
  MUX21X1 U15621 ( .IN1(\mem2[85][18] ), .IN2(n1099), .S(n8140), .Q(n11094) );
  MUX21X1 U15622 ( .IN1(\mem2[85][17] ), .IN2(n1077), .S(n8140), .Q(n11093) );
  MUX21X1 U15623 ( .IN1(\mem2[85][16] ), .IN2(n1055), .S(n8140), .Q(n11092) );
  AND2X1 U15624 ( .IN1(n8130), .IN2(n7120), .Q(n8140) );
  MUX21X1 U15625 ( .IN1(\mem2[84][23] ), .IN2(n1209), .S(n8141), .Q(n11091) );
  MUX21X1 U15626 ( .IN1(\mem2[84][22] ), .IN2(n1187), .S(n8141), .Q(n11090) );
  MUX21X1 U15627 ( .IN1(\mem2[84][21] ), .IN2(n1165), .S(n8141), .Q(n11089) );
  MUX21X1 U15628 ( .IN1(\mem2[84][20] ), .IN2(n1143), .S(n8141), .Q(n11088) );
  MUX21X1 U15629 ( .IN1(\mem2[84][19] ), .IN2(n1121), .S(n8141), .Q(n11087) );
  MUX21X1 U15630 ( .IN1(\mem2[84][18] ), .IN2(n1099), .S(n8141), .Q(n11086) );
  MUX21X1 U15631 ( .IN1(\mem2[84][17] ), .IN2(n1077), .S(n8141), .Q(n11085) );
  MUX21X1 U15632 ( .IN1(\mem2[84][16] ), .IN2(n1055), .S(n8141), .Q(n11084) );
  AND2X1 U15633 ( .IN1(n8130), .IN2(n7122), .Q(n8141) );
  MUX21X1 U15634 ( .IN1(\mem2[83][23] ), .IN2(n1209), .S(n8142), .Q(n11083) );
  MUX21X1 U15635 ( .IN1(\mem2[83][22] ), .IN2(n1187), .S(n8142), .Q(n11082) );
  MUX21X1 U15636 ( .IN1(\mem2[83][21] ), .IN2(n1165), .S(n8142), .Q(n11081) );
  MUX21X1 U15637 ( .IN1(\mem2[83][20] ), .IN2(n1143), .S(n8142), .Q(n11080) );
  MUX21X1 U15638 ( .IN1(\mem2[83][19] ), .IN2(n1121), .S(n8142), .Q(n11079) );
  MUX21X1 U15639 ( .IN1(\mem2[83][18] ), .IN2(n1099), .S(n8142), .Q(n11078) );
  MUX21X1 U15640 ( .IN1(\mem2[83][17] ), .IN2(n1077), .S(n8142), .Q(n11077) );
  MUX21X1 U15641 ( .IN1(\mem2[83][16] ), .IN2(n1055), .S(n8142), .Q(n11076) );
  AND2X1 U15642 ( .IN1(n8130), .IN2(n7124), .Q(n8142) );
  MUX21X1 U15643 ( .IN1(\mem2[82][23] ), .IN2(n1209), .S(n8143), .Q(n11075) );
  MUX21X1 U15644 ( .IN1(\mem2[82][22] ), .IN2(n1187), .S(n8143), .Q(n11074) );
  MUX21X1 U15645 ( .IN1(\mem2[82][21] ), .IN2(n1165), .S(n8143), .Q(n11073) );
  MUX21X1 U15646 ( .IN1(\mem2[82][20] ), .IN2(n1143), .S(n8143), .Q(n11072) );
  MUX21X1 U15647 ( .IN1(\mem2[82][19] ), .IN2(n1121), .S(n8143), .Q(n11071) );
  MUX21X1 U15648 ( .IN1(\mem2[82][18] ), .IN2(n1099), .S(n8143), .Q(n11070) );
  MUX21X1 U15649 ( .IN1(\mem2[82][17] ), .IN2(n1077), .S(n8143), .Q(n11069) );
  MUX21X1 U15650 ( .IN1(\mem2[82][16] ), .IN2(n1055), .S(n8143), .Q(n11068) );
  AND2X1 U15651 ( .IN1(n8130), .IN2(n7126), .Q(n8143) );
  MUX21X1 U15652 ( .IN1(\mem2[81][23] ), .IN2(n1209), .S(n8144), .Q(n11067) );
  MUX21X1 U15653 ( .IN1(\mem2[81][22] ), .IN2(n1187), .S(n8144), .Q(n11066) );
  MUX21X1 U15654 ( .IN1(\mem2[81][21] ), .IN2(n1165), .S(n8144), .Q(n11065) );
  MUX21X1 U15655 ( .IN1(\mem2[81][20] ), .IN2(n1143), .S(n8144), .Q(n11064) );
  MUX21X1 U15656 ( .IN1(\mem2[81][19] ), .IN2(n1121), .S(n8144), .Q(n11063) );
  MUX21X1 U15657 ( .IN1(\mem2[81][18] ), .IN2(n1099), .S(n8144), .Q(n11062) );
  MUX21X1 U15658 ( .IN1(\mem2[81][17] ), .IN2(n1077), .S(n8144), .Q(n11061) );
  MUX21X1 U15659 ( .IN1(\mem2[81][16] ), .IN2(n1055), .S(n8144), .Q(n11060) );
  AND2X1 U15660 ( .IN1(n8130), .IN2(n7128), .Q(n8144) );
  MUX21X1 U15661 ( .IN1(\mem2[80][23] ), .IN2(n1209), .S(n8145), .Q(n11059) );
  MUX21X1 U15662 ( .IN1(\mem2[80][22] ), .IN2(n1187), .S(n8145), .Q(n11058) );
  MUX21X1 U15663 ( .IN1(\mem2[80][21] ), .IN2(n1165), .S(n8145), .Q(n11057) );
  MUX21X1 U15664 ( .IN1(\mem2[80][20] ), .IN2(n1143), .S(n8145), .Q(n11056) );
  MUX21X1 U15665 ( .IN1(\mem2[80][19] ), .IN2(n1121), .S(n8145), .Q(n11055) );
  MUX21X1 U15666 ( .IN1(\mem2[80][18] ), .IN2(n1099), .S(n8145), .Q(n11054) );
  MUX21X1 U15667 ( .IN1(\mem2[80][17] ), .IN2(n1077), .S(n8145), .Q(n11053) );
  MUX21X1 U15668 ( .IN1(\mem2[80][16] ), .IN2(n1055), .S(n8145), .Q(n11052) );
  AND2X1 U15669 ( .IN1(n8130), .IN2(n7130), .Q(n8145) );
  AND2X1 U15670 ( .IN1(n7966), .IN2(n7312), .Q(n8130) );
  AND2X1 U15671 ( .IN1(n8111), .IN2(n8004), .Q(n7312) );
  MUX21X1 U15672 ( .IN1(\mem2[79][23] ), .IN2(n1209), .S(n8146), .Q(n11051) );
  MUX21X1 U15673 ( .IN1(\mem2[79][22] ), .IN2(n1187), .S(n8146), .Q(n11050) );
  MUX21X1 U15674 ( .IN1(\mem2[79][21] ), .IN2(n1165), .S(n8146), .Q(n11049) );
  MUX21X1 U15675 ( .IN1(\mem2[79][20] ), .IN2(n1143), .S(n8146), .Q(n11048) );
  MUX21X1 U15676 ( .IN1(\mem2[79][19] ), .IN2(n1121), .S(n8146), .Q(n11047) );
  MUX21X1 U15677 ( .IN1(\mem2[79][18] ), .IN2(n1099), .S(n8146), .Q(n11046) );
  MUX21X1 U15678 ( .IN1(\mem2[79][17] ), .IN2(n1077), .S(n8146), .Q(n11045) );
  MUX21X1 U15679 ( .IN1(\mem2[79][16] ), .IN2(n1055), .S(n8146), .Q(n11044) );
  AND2X1 U15680 ( .IN1(n8147), .IN2(n7099), .Q(n8146) );
  MUX21X1 U15681 ( .IN1(\mem2[78][23] ), .IN2(n1209), .S(n8148), .Q(n11043) );
  MUX21X1 U15682 ( .IN1(\mem2[78][22] ), .IN2(n1187), .S(n8148), .Q(n11042) );
  MUX21X1 U15683 ( .IN1(\mem2[78][21] ), .IN2(n1165), .S(n8148), .Q(n11041) );
  MUX21X1 U15684 ( .IN1(\mem2[78][20] ), .IN2(n1143), .S(n8148), .Q(n11040) );
  MUX21X1 U15685 ( .IN1(\mem2[78][19] ), .IN2(n1121), .S(n8148), .Q(n11039) );
  MUX21X1 U15686 ( .IN1(\mem2[78][18] ), .IN2(n1099), .S(n8148), .Q(n11038) );
  MUX21X1 U15687 ( .IN1(\mem2[78][17] ), .IN2(n1077), .S(n8148), .Q(n11037) );
  MUX21X1 U15688 ( .IN1(\mem2[78][16] ), .IN2(n1055), .S(n8148), .Q(n11036) );
  AND2X1 U15689 ( .IN1(n8147), .IN2(n7102), .Q(n8148) );
  MUX21X1 U15690 ( .IN1(\mem2[77][23] ), .IN2(n1209), .S(n8149), .Q(n11035) );
  MUX21X1 U15691 ( .IN1(\mem2[77][22] ), .IN2(n1187), .S(n8149), .Q(n11034) );
  MUX21X1 U15692 ( .IN1(\mem2[77][21] ), .IN2(n1165), .S(n8149), .Q(n11033) );
  MUX21X1 U15693 ( .IN1(\mem2[77][20] ), .IN2(n1143), .S(n8149), .Q(n11032) );
  MUX21X1 U15694 ( .IN1(\mem2[77][19] ), .IN2(n1121), .S(n8149), .Q(n11031) );
  MUX21X1 U15695 ( .IN1(\mem2[77][18] ), .IN2(n1099), .S(n8149), .Q(n11030) );
  MUX21X1 U15696 ( .IN1(\mem2[77][17] ), .IN2(n1077), .S(n8149), .Q(n11029) );
  MUX21X1 U15697 ( .IN1(\mem2[77][16] ), .IN2(n1055), .S(n8149), .Q(n11028) );
  AND2X1 U15698 ( .IN1(n8147), .IN2(n7104), .Q(n8149) );
  MUX21X1 U15699 ( .IN1(\mem2[76][23] ), .IN2(n1209), .S(n8150), .Q(n11027) );
  MUX21X1 U15700 ( .IN1(\mem2[76][22] ), .IN2(n1187), .S(n8150), .Q(n11026) );
  MUX21X1 U15701 ( .IN1(\mem2[76][21] ), .IN2(n1165), .S(n8150), .Q(n11025) );
  MUX21X1 U15702 ( .IN1(\mem2[76][20] ), .IN2(n1143), .S(n8150), .Q(n11024) );
  MUX21X1 U15703 ( .IN1(\mem2[76][19] ), .IN2(n1121), .S(n8150), .Q(n11023) );
  MUX21X1 U15704 ( .IN1(\mem2[76][18] ), .IN2(n1099), .S(n8150), .Q(n11022) );
  MUX21X1 U15705 ( .IN1(\mem2[76][17] ), .IN2(n1077), .S(n8150), .Q(n11021) );
  MUX21X1 U15706 ( .IN1(\mem2[76][16] ), .IN2(n1055), .S(n8150), .Q(n11020) );
  AND2X1 U15707 ( .IN1(n8147), .IN2(n7106), .Q(n8150) );
  MUX21X1 U15708 ( .IN1(\mem2[75][23] ), .IN2(n1210), .S(n8151), .Q(n11019) );
  MUX21X1 U15709 ( .IN1(\mem2[75][22] ), .IN2(n1188), .S(n8151), .Q(n11018) );
  MUX21X1 U15710 ( .IN1(\mem2[75][21] ), .IN2(n1166), .S(n8151), .Q(n11017) );
  MUX21X1 U15711 ( .IN1(\mem2[75][20] ), .IN2(n1144), .S(n8151), .Q(n11016) );
  MUX21X1 U15712 ( .IN1(\mem2[75][19] ), .IN2(n1122), .S(n8151), .Q(n11015) );
  MUX21X1 U15713 ( .IN1(\mem2[75][18] ), .IN2(n1100), .S(n8151), .Q(n11014) );
  MUX21X1 U15714 ( .IN1(\mem2[75][17] ), .IN2(n1078), .S(n8151), .Q(n11013) );
  MUX21X1 U15715 ( .IN1(\mem2[75][16] ), .IN2(n1056), .S(n8151), .Q(n11012) );
  AND2X1 U15716 ( .IN1(n8147), .IN2(n7108), .Q(n8151) );
  MUX21X1 U15717 ( .IN1(\mem2[74][23] ), .IN2(n1210), .S(n8152), .Q(n11011) );
  MUX21X1 U15718 ( .IN1(\mem2[74][22] ), .IN2(n1188), .S(n8152), .Q(n11010) );
  MUX21X1 U15719 ( .IN1(\mem2[74][21] ), .IN2(n1166), .S(n8152), .Q(n11009) );
  MUX21X1 U15720 ( .IN1(\mem2[74][20] ), .IN2(n1144), .S(n8152), .Q(n11008) );
  MUX21X1 U15721 ( .IN1(\mem2[74][19] ), .IN2(n1122), .S(n8152), .Q(n11007) );
  MUX21X1 U15722 ( .IN1(\mem2[74][18] ), .IN2(n1100), .S(n8152), .Q(n11006) );
  MUX21X1 U15723 ( .IN1(\mem2[74][17] ), .IN2(n1078), .S(n8152), .Q(n11005) );
  MUX21X1 U15724 ( .IN1(\mem2[74][16] ), .IN2(n1056), .S(n8152), .Q(n11004) );
  AND2X1 U15725 ( .IN1(n8147), .IN2(n7110), .Q(n8152) );
  MUX21X1 U15726 ( .IN1(\mem2[73][23] ), .IN2(n1210), .S(n8153), .Q(n11003) );
  MUX21X1 U15727 ( .IN1(\mem2[73][22] ), .IN2(n1188), .S(n8153), .Q(n11002) );
  MUX21X1 U15728 ( .IN1(\mem2[73][21] ), .IN2(n1166), .S(n8153), .Q(n11001) );
  MUX21X1 U15729 ( .IN1(\mem2[73][20] ), .IN2(n1144), .S(n8153), .Q(n11000) );
  MUX21X1 U15730 ( .IN1(\mem2[73][19] ), .IN2(n1122), .S(n8153), .Q(n10999) );
  MUX21X1 U15731 ( .IN1(\mem2[73][18] ), .IN2(n1100), .S(n8153), .Q(n10998) );
  MUX21X1 U15732 ( .IN1(\mem2[73][17] ), .IN2(n1078), .S(n8153), .Q(n10997) );
  MUX21X1 U15733 ( .IN1(\mem2[73][16] ), .IN2(n1056), .S(n8153), .Q(n10996) );
  AND2X1 U15734 ( .IN1(n8147), .IN2(n7112), .Q(n8153) );
  MUX21X1 U15735 ( .IN1(\mem2[72][23] ), .IN2(n1210), .S(n8154), .Q(n10995) );
  MUX21X1 U15736 ( .IN1(\mem2[72][22] ), .IN2(n1188), .S(n8154), .Q(n10994) );
  MUX21X1 U15737 ( .IN1(\mem2[72][21] ), .IN2(n1166), .S(n8154), .Q(n10993) );
  MUX21X1 U15738 ( .IN1(\mem2[72][20] ), .IN2(n1144), .S(n8154), .Q(n10992) );
  MUX21X1 U15739 ( .IN1(\mem2[72][19] ), .IN2(n1122), .S(n8154), .Q(n10991) );
  MUX21X1 U15740 ( .IN1(\mem2[72][18] ), .IN2(n1100), .S(n8154), .Q(n10990) );
  MUX21X1 U15741 ( .IN1(\mem2[72][17] ), .IN2(n1078), .S(n8154), .Q(n10989) );
  MUX21X1 U15742 ( .IN1(\mem2[72][16] ), .IN2(n1056), .S(n8154), .Q(n10988) );
  AND2X1 U15743 ( .IN1(n8147), .IN2(n7114), .Q(n8154) );
  MUX21X1 U15744 ( .IN1(\mem2[71][23] ), .IN2(n1210), .S(n8155), .Q(n10987) );
  MUX21X1 U15745 ( .IN1(\mem2[71][22] ), .IN2(n1188), .S(n8155), .Q(n10986) );
  MUX21X1 U15746 ( .IN1(\mem2[71][21] ), .IN2(n1166), .S(n8155), .Q(n10985) );
  MUX21X1 U15747 ( .IN1(\mem2[71][20] ), .IN2(n1144), .S(n8155), .Q(n10984) );
  MUX21X1 U15748 ( .IN1(\mem2[71][19] ), .IN2(n1122), .S(n8155), .Q(n10983) );
  MUX21X1 U15749 ( .IN1(\mem2[71][18] ), .IN2(n1100), .S(n8155), .Q(n10982) );
  MUX21X1 U15750 ( .IN1(\mem2[71][17] ), .IN2(n1078), .S(n8155), .Q(n10981) );
  MUX21X1 U15751 ( .IN1(\mem2[71][16] ), .IN2(n1056), .S(n8155), .Q(n10980) );
  AND2X1 U15752 ( .IN1(n8147), .IN2(n7116), .Q(n8155) );
  MUX21X1 U15753 ( .IN1(\mem2[70][23] ), .IN2(n1210), .S(n8156), .Q(n10979) );
  MUX21X1 U15754 ( .IN1(\mem2[70][22] ), .IN2(n1188), .S(n8156), .Q(n10978) );
  MUX21X1 U15755 ( .IN1(\mem2[70][21] ), .IN2(n1166), .S(n8156), .Q(n10977) );
  MUX21X1 U15756 ( .IN1(\mem2[70][20] ), .IN2(n1144), .S(n8156), .Q(n10976) );
  MUX21X1 U15757 ( .IN1(\mem2[70][19] ), .IN2(n1122), .S(n8156), .Q(n10975) );
  MUX21X1 U15758 ( .IN1(\mem2[70][18] ), .IN2(n1100), .S(n8156), .Q(n10974) );
  MUX21X1 U15759 ( .IN1(\mem2[70][17] ), .IN2(n1078), .S(n8156), .Q(n10973) );
  MUX21X1 U15760 ( .IN1(\mem2[70][16] ), .IN2(n1056), .S(n8156), .Q(n10972) );
  AND2X1 U15761 ( .IN1(n8147), .IN2(n7118), .Q(n8156) );
  MUX21X1 U15762 ( .IN1(\mem2[69][23] ), .IN2(n1210), .S(n8157), .Q(n10971) );
  MUX21X1 U15763 ( .IN1(\mem2[69][22] ), .IN2(n1188), .S(n8157), .Q(n10970) );
  MUX21X1 U15764 ( .IN1(\mem2[69][21] ), .IN2(n1166), .S(n8157), .Q(n10969) );
  MUX21X1 U15765 ( .IN1(\mem2[69][20] ), .IN2(n1144), .S(n8157), .Q(n10968) );
  MUX21X1 U15766 ( .IN1(\mem2[69][19] ), .IN2(n1122), .S(n8157), .Q(n10967) );
  MUX21X1 U15767 ( .IN1(\mem2[69][18] ), .IN2(n1100), .S(n8157), .Q(n10966) );
  MUX21X1 U15768 ( .IN1(\mem2[69][17] ), .IN2(n1078), .S(n8157), .Q(n10965) );
  MUX21X1 U15769 ( .IN1(\mem2[69][16] ), .IN2(n1056), .S(n8157), .Q(n10964) );
  AND2X1 U15770 ( .IN1(n8147), .IN2(n7120), .Q(n8157) );
  MUX21X1 U15771 ( .IN1(\mem2[68][23] ), .IN2(n1210), .S(n8158), .Q(n10963) );
  MUX21X1 U15772 ( .IN1(\mem2[68][22] ), .IN2(n1188), .S(n8158), .Q(n10962) );
  MUX21X1 U15773 ( .IN1(\mem2[68][21] ), .IN2(n1166), .S(n8158), .Q(n10961) );
  MUX21X1 U15774 ( .IN1(\mem2[68][20] ), .IN2(n1144), .S(n8158), .Q(n10960) );
  MUX21X1 U15775 ( .IN1(\mem2[68][19] ), .IN2(n1122), .S(n8158), .Q(n10959) );
  MUX21X1 U15776 ( .IN1(\mem2[68][18] ), .IN2(n1100), .S(n8158), .Q(n10958) );
  MUX21X1 U15777 ( .IN1(\mem2[68][17] ), .IN2(n1078), .S(n8158), .Q(n10957) );
  MUX21X1 U15778 ( .IN1(\mem2[68][16] ), .IN2(n1056), .S(n8158), .Q(n10956) );
  AND2X1 U15779 ( .IN1(n8147), .IN2(n7122), .Q(n8158) );
  MUX21X1 U15780 ( .IN1(\mem2[67][23] ), .IN2(n1210), .S(n8159), .Q(n10955) );
  MUX21X1 U15781 ( .IN1(\mem2[67][22] ), .IN2(n1188), .S(n8159), .Q(n10954) );
  MUX21X1 U15782 ( .IN1(\mem2[67][21] ), .IN2(n1166), .S(n8159), .Q(n10953) );
  MUX21X1 U15783 ( .IN1(\mem2[67][20] ), .IN2(n1144), .S(n8159), .Q(n10952) );
  MUX21X1 U15784 ( .IN1(\mem2[67][19] ), .IN2(n1122), .S(n8159), .Q(n10951) );
  MUX21X1 U15785 ( .IN1(\mem2[67][18] ), .IN2(n1100), .S(n8159), .Q(n10950) );
  MUX21X1 U15786 ( .IN1(\mem2[67][17] ), .IN2(n1078), .S(n8159), .Q(n10949) );
  MUX21X1 U15787 ( .IN1(\mem2[67][16] ), .IN2(n1056), .S(n8159), .Q(n10948) );
  AND2X1 U15788 ( .IN1(n8147), .IN2(n7124), .Q(n8159) );
  MUX21X1 U15789 ( .IN1(\mem2[66][23] ), .IN2(n1210), .S(n8160), .Q(n10947) );
  MUX21X1 U15790 ( .IN1(\mem2[66][22] ), .IN2(n1188), .S(n8160), .Q(n10946) );
  MUX21X1 U15791 ( .IN1(\mem2[66][21] ), .IN2(n1166), .S(n8160), .Q(n10945) );
  MUX21X1 U15792 ( .IN1(\mem2[66][20] ), .IN2(n1144), .S(n8160), .Q(n10944) );
  MUX21X1 U15793 ( .IN1(\mem2[66][19] ), .IN2(n1122), .S(n8160), .Q(n10943) );
  MUX21X1 U15794 ( .IN1(\mem2[66][18] ), .IN2(n1100), .S(n8160), .Q(n10942) );
  MUX21X1 U15795 ( .IN1(\mem2[66][17] ), .IN2(n1078), .S(n8160), .Q(n10941) );
  MUX21X1 U15796 ( .IN1(\mem2[66][16] ), .IN2(n1056), .S(n8160), .Q(n10940) );
  AND2X1 U15797 ( .IN1(n8147), .IN2(n7126), .Q(n8160) );
  MUX21X1 U15798 ( .IN1(\mem2[65][23] ), .IN2(n1210), .S(n8161), .Q(n10939) );
  MUX21X1 U15799 ( .IN1(\mem2[65][22] ), .IN2(n1188), .S(n8161), .Q(n10938) );
  MUX21X1 U15800 ( .IN1(\mem2[65][21] ), .IN2(n1166), .S(n8161), .Q(n10937) );
  MUX21X1 U15801 ( .IN1(\mem2[65][20] ), .IN2(n1144), .S(n8161), .Q(n10936) );
  MUX21X1 U15802 ( .IN1(\mem2[65][19] ), .IN2(n1122), .S(n8161), .Q(n10935) );
  MUX21X1 U15803 ( .IN1(\mem2[65][18] ), .IN2(n1100), .S(n8161), .Q(n10934) );
  MUX21X1 U15804 ( .IN1(\mem2[65][17] ), .IN2(n1078), .S(n8161), .Q(n10933) );
  MUX21X1 U15805 ( .IN1(\mem2[65][16] ), .IN2(n1056), .S(n8161), .Q(n10932) );
  AND2X1 U15806 ( .IN1(n8147), .IN2(n7128), .Q(n8161) );
  MUX21X1 U15807 ( .IN1(\mem2[64][23] ), .IN2(n1210), .S(n8162), .Q(n10931) );
  MUX21X1 U15808 ( .IN1(\mem2[64][22] ), .IN2(n1188), .S(n8162), .Q(n10930) );
  MUX21X1 U15809 ( .IN1(\mem2[64][21] ), .IN2(n1166), .S(n8162), .Q(n10929) );
  MUX21X1 U15810 ( .IN1(\mem2[64][20] ), .IN2(n1144), .S(n8162), .Q(n10928) );
  MUX21X1 U15811 ( .IN1(\mem2[64][19] ), .IN2(n1122), .S(n8162), .Q(n10927) );
  MUX21X1 U15812 ( .IN1(\mem2[64][18] ), .IN2(n1100), .S(n8162), .Q(n10926) );
  MUX21X1 U15813 ( .IN1(\mem2[64][17] ), .IN2(n1078), .S(n8162), .Q(n10925) );
  MUX21X1 U15814 ( .IN1(\mem2[64][16] ), .IN2(n1056), .S(n8162), .Q(n10924) );
  AND2X1 U15815 ( .IN1(n8147), .IN2(n7130), .Q(n8162) );
  AND2X1 U15816 ( .IN1(n7966), .IN2(n7330), .Q(n8147) );
  AND2X1 U15817 ( .IN1(n8111), .IN2(n8022), .Q(n7330) );
  NOR2X0 U15818 ( .IN1(n8024), .IN2(addr[7]), .QN(n8111) );
  INVX0 U15819 ( .INP(addr[6]), .ZN(n8024) );
  MUX21X1 U15820 ( .IN1(\mem2[63][23] ), .IN2(n1211), .S(n8163), .Q(n10923) );
  MUX21X1 U15821 ( .IN1(\mem2[63][22] ), .IN2(n1189), .S(n8163), .Q(n10922) );
  MUX21X1 U15822 ( .IN1(\mem2[63][21] ), .IN2(n1167), .S(n8163), .Q(n10921) );
  MUX21X1 U15823 ( .IN1(\mem2[63][20] ), .IN2(n1145), .S(n8163), .Q(n10920) );
  MUX21X1 U15824 ( .IN1(\mem2[63][19] ), .IN2(n1123), .S(n8163), .Q(n10919) );
  MUX21X1 U15825 ( .IN1(\mem2[63][18] ), .IN2(n1101), .S(n8163), .Q(n10918) );
  MUX21X1 U15826 ( .IN1(\mem2[63][17] ), .IN2(n1079), .S(n8163), .Q(n10917) );
  MUX21X1 U15827 ( .IN1(\mem2[63][16] ), .IN2(n1057), .S(n8163), .Q(n10916) );
  AND2X1 U15828 ( .IN1(n8164), .IN2(n7099), .Q(n8163) );
  MUX21X1 U15829 ( .IN1(\mem2[62][23] ), .IN2(n1211), .S(n8165), .Q(n10915) );
  MUX21X1 U15830 ( .IN1(\mem2[62][22] ), .IN2(n1189), .S(n8165), .Q(n10914) );
  MUX21X1 U15831 ( .IN1(\mem2[62][21] ), .IN2(n1167), .S(n8165), .Q(n10913) );
  MUX21X1 U15832 ( .IN1(\mem2[62][20] ), .IN2(n1145), .S(n8165), .Q(n10912) );
  MUX21X1 U15833 ( .IN1(\mem2[62][19] ), .IN2(n1123), .S(n8165), .Q(n10911) );
  MUX21X1 U15834 ( .IN1(\mem2[62][18] ), .IN2(n1101), .S(n8165), .Q(n10910) );
  MUX21X1 U15835 ( .IN1(\mem2[62][17] ), .IN2(n1079), .S(n8165), .Q(n10909) );
  MUX21X1 U15836 ( .IN1(\mem2[62][16] ), .IN2(n1057), .S(n8165), .Q(n10908) );
  AND2X1 U15837 ( .IN1(n8164), .IN2(n7102), .Q(n8165) );
  MUX21X1 U15838 ( .IN1(\mem2[61][23] ), .IN2(n1211), .S(n8166), .Q(n10907) );
  MUX21X1 U15839 ( .IN1(\mem2[61][22] ), .IN2(n1189), .S(n8166), .Q(n10906) );
  MUX21X1 U15840 ( .IN1(\mem2[61][21] ), .IN2(n1167), .S(n8166), .Q(n10905) );
  MUX21X1 U15841 ( .IN1(\mem2[61][20] ), .IN2(n1145), .S(n8166), .Q(n10904) );
  MUX21X1 U15842 ( .IN1(\mem2[61][19] ), .IN2(n1123), .S(n8166), .Q(n10903) );
  MUX21X1 U15843 ( .IN1(\mem2[61][18] ), .IN2(n1101), .S(n8166), .Q(n10902) );
  MUX21X1 U15844 ( .IN1(\mem2[61][17] ), .IN2(n1079), .S(n8166), .Q(n10901) );
  MUX21X1 U15845 ( .IN1(\mem2[61][16] ), .IN2(n1057), .S(n8166), .Q(n10900) );
  AND2X1 U15846 ( .IN1(n8164), .IN2(n7104), .Q(n8166) );
  MUX21X1 U15847 ( .IN1(\mem2[60][23] ), .IN2(n1211), .S(n8167), .Q(n10899) );
  MUX21X1 U15848 ( .IN1(\mem2[60][22] ), .IN2(n1189), .S(n8167), .Q(n10898) );
  MUX21X1 U15849 ( .IN1(\mem2[60][21] ), .IN2(n1167), .S(n8167), .Q(n10897) );
  MUX21X1 U15850 ( .IN1(\mem2[60][20] ), .IN2(n1145), .S(n8167), .Q(n10896) );
  MUX21X1 U15851 ( .IN1(\mem2[60][19] ), .IN2(n1123), .S(n8167), .Q(n10895) );
  MUX21X1 U15852 ( .IN1(\mem2[60][18] ), .IN2(n1101), .S(n8167), .Q(n10894) );
  MUX21X1 U15853 ( .IN1(\mem2[60][17] ), .IN2(n1079), .S(n8167), .Q(n10893) );
  MUX21X1 U15854 ( .IN1(\mem2[60][16] ), .IN2(n1057), .S(n8167), .Q(n10892) );
  AND2X1 U15855 ( .IN1(n8164), .IN2(n7106), .Q(n8167) );
  MUX21X1 U15856 ( .IN1(\mem2[59][23] ), .IN2(n1211), .S(n8168), .Q(n10891) );
  MUX21X1 U15857 ( .IN1(\mem2[59][22] ), .IN2(n1189), .S(n8168), .Q(n10890) );
  MUX21X1 U15858 ( .IN1(\mem2[59][21] ), .IN2(n1167), .S(n8168), .Q(n10889) );
  MUX21X1 U15859 ( .IN1(\mem2[59][20] ), .IN2(n1145), .S(n8168), .Q(n10888) );
  MUX21X1 U15860 ( .IN1(\mem2[59][19] ), .IN2(n1123), .S(n8168), .Q(n10887) );
  MUX21X1 U15861 ( .IN1(\mem2[59][18] ), .IN2(n1101), .S(n8168), .Q(n10886) );
  MUX21X1 U15862 ( .IN1(\mem2[59][17] ), .IN2(n1079), .S(n8168), .Q(n10885) );
  MUX21X1 U15863 ( .IN1(\mem2[59][16] ), .IN2(n1057), .S(n8168), .Q(n10884) );
  AND2X1 U15864 ( .IN1(n8164), .IN2(n7108), .Q(n8168) );
  MUX21X1 U15865 ( .IN1(\mem2[58][23] ), .IN2(n1211), .S(n8169), .Q(n10883) );
  MUX21X1 U15866 ( .IN1(\mem2[58][22] ), .IN2(n1189), .S(n8169), .Q(n10882) );
  MUX21X1 U15867 ( .IN1(\mem2[58][21] ), .IN2(n1167), .S(n8169), .Q(n10881) );
  MUX21X1 U15868 ( .IN1(\mem2[58][20] ), .IN2(n1145), .S(n8169), .Q(n10880) );
  MUX21X1 U15869 ( .IN1(\mem2[58][19] ), .IN2(n1123), .S(n8169), .Q(n10879) );
  MUX21X1 U15870 ( .IN1(\mem2[58][18] ), .IN2(n1101), .S(n8169), .Q(n10878) );
  MUX21X1 U15871 ( .IN1(\mem2[58][17] ), .IN2(n1079), .S(n8169), .Q(n10877) );
  MUX21X1 U15872 ( .IN1(\mem2[58][16] ), .IN2(n1057), .S(n8169), .Q(n10876) );
  AND2X1 U15873 ( .IN1(n8164), .IN2(n7110), .Q(n8169) );
  MUX21X1 U15874 ( .IN1(\mem2[57][23] ), .IN2(n1211), .S(n8170), .Q(n10875) );
  MUX21X1 U15875 ( .IN1(\mem2[57][22] ), .IN2(n1189), .S(n8170), .Q(n10874) );
  MUX21X1 U15876 ( .IN1(\mem2[57][21] ), .IN2(n1167), .S(n8170), .Q(n10873) );
  MUX21X1 U15877 ( .IN1(\mem2[57][20] ), .IN2(n1145), .S(n8170), .Q(n10872) );
  MUX21X1 U15878 ( .IN1(\mem2[57][19] ), .IN2(n1123), .S(n8170), .Q(n10871) );
  MUX21X1 U15879 ( .IN1(\mem2[57][18] ), .IN2(n1101), .S(n8170), .Q(n10870) );
  MUX21X1 U15880 ( .IN1(\mem2[57][17] ), .IN2(n1079), .S(n8170), .Q(n10869) );
  MUX21X1 U15881 ( .IN1(\mem2[57][16] ), .IN2(n1057), .S(n8170), .Q(n10868) );
  AND2X1 U15882 ( .IN1(n8164), .IN2(n7112), .Q(n8170) );
  MUX21X1 U15883 ( .IN1(\mem2[56][23] ), .IN2(n1211), .S(n8171), .Q(n10867) );
  MUX21X1 U15884 ( .IN1(\mem2[56][22] ), .IN2(n1189), .S(n8171), .Q(n10866) );
  MUX21X1 U15885 ( .IN1(\mem2[56][21] ), .IN2(n1167), .S(n8171), .Q(n10865) );
  MUX21X1 U15886 ( .IN1(\mem2[56][20] ), .IN2(n1145), .S(n8171), .Q(n10864) );
  MUX21X1 U15887 ( .IN1(\mem2[56][19] ), .IN2(n1123), .S(n8171), .Q(n10863) );
  MUX21X1 U15888 ( .IN1(\mem2[56][18] ), .IN2(n1101), .S(n8171), .Q(n10862) );
  MUX21X1 U15889 ( .IN1(\mem2[56][17] ), .IN2(n1079), .S(n8171), .Q(n10861) );
  MUX21X1 U15890 ( .IN1(\mem2[56][16] ), .IN2(n1057), .S(n8171), .Q(n10860) );
  AND2X1 U15891 ( .IN1(n8164), .IN2(n7114), .Q(n8171) );
  MUX21X1 U15892 ( .IN1(\mem2[55][23] ), .IN2(n1211), .S(n8172), .Q(n10859) );
  MUX21X1 U15893 ( .IN1(\mem2[55][22] ), .IN2(n1189), .S(n8172), .Q(n10858) );
  MUX21X1 U15894 ( .IN1(\mem2[55][21] ), .IN2(n1167), .S(n8172), .Q(n10857) );
  MUX21X1 U15895 ( .IN1(\mem2[55][20] ), .IN2(n1145), .S(n8172), .Q(n10856) );
  MUX21X1 U15896 ( .IN1(\mem2[55][19] ), .IN2(n1123), .S(n8172), .Q(n10855) );
  MUX21X1 U15897 ( .IN1(\mem2[55][18] ), .IN2(n1101), .S(n8172), .Q(n10854) );
  MUX21X1 U15898 ( .IN1(\mem2[55][17] ), .IN2(n1079), .S(n8172), .Q(n10853) );
  MUX21X1 U15899 ( .IN1(\mem2[55][16] ), .IN2(n1057), .S(n8172), .Q(n10852) );
  AND2X1 U15900 ( .IN1(n8164), .IN2(n7116), .Q(n8172) );
  MUX21X1 U15901 ( .IN1(\mem2[54][23] ), .IN2(n1211), .S(n8173), .Q(n10851) );
  MUX21X1 U15902 ( .IN1(\mem2[54][22] ), .IN2(n1189), .S(n8173), .Q(n10850) );
  MUX21X1 U15903 ( .IN1(\mem2[54][21] ), .IN2(n1167), .S(n8173), .Q(n10849) );
  MUX21X1 U15904 ( .IN1(\mem2[54][20] ), .IN2(n1145), .S(n8173), .Q(n10848) );
  MUX21X1 U15905 ( .IN1(\mem2[54][19] ), .IN2(n1123), .S(n8173), .Q(n10847) );
  MUX21X1 U15906 ( .IN1(\mem2[54][18] ), .IN2(n1101), .S(n8173), .Q(n10846) );
  MUX21X1 U15907 ( .IN1(\mem2[54][17] ), .IN2(n1079), .S(n8173), .Q(n10845) );
  MUX21X1 U15908 ( .IN1(\mem2[54][16] ), .IN2(n1057), .S(n8173), .Q(n10844) );
  AND2X1 U15909 ( .IN1(n8164), .IN2(n7118), .Q(n8173) );
  MUX21X1 U15910 ( .IN1(\mem2[53][23] ), .IN2(n1211), .S(n8174), .Q(n10843) );
  MUX21X1 U15911 ( .IN1(\mem2[53][22] ), .IN2(n1189), .S(n8174), .Q(n10842) );
  MUX21X1 U15912 ( .IN1(\mem2[53][21] ), .IN2(n1167), .S(n8174), .Q(n10841) );
  MUX21X1 U15913 ( .IN1(\mem2[53][20] ), .IN2(n1145), .S(n8174), .Q(n10840) );
  MUX21X1 U15914 ( .IN1(\mem2[53][19] ), .IN2(n1123), .S(n8174), .Q(n10839) );
  MUX21X1 U15915 ( .IN1(\mem2[53][18] ), .IN2(n1101), .S(n8174), .Q(n10838) );
  MUX21X1 U15916 ( .IN1(\mem2[53][17] ), .IN2(n1079), .S(n8174), .Q(n10837) );
  MUX21X1 U15917 ( .IN1(\mem2[53][16] ), .IN2(n1057), .S(n8174), .Q(n10836) );
  AND2X1 U15918 ( .IN1(n8164), .IN2(n7120), .Q(n8174) );
  MUX21X1 U15919 ( .IN1(\mem2[52][23] ), .IN2(n1211), .S(n8175), .Q(n10835) );
  MUX21X1 U15920 ( .IN1(\mem2[52][22] ), .IN2(n1189), .S(n8175), .Q(n10834) );
  MUX21X1 U15921 ( .IN1(\mem2[52][21] ), .IN2(n1167), .S(n8175), .Q(n10833) );
  MUX21X1 U15922 ( .IN1(\mem2[52][20] ), .IN2(n1145), .S(n8175), .Q(n10832) );
  MUX21X1 U15923 ( .IN1(\mem2[52][19] ), .IN2(n1123), .S(n8175), .Q(n10831) );
  MUX21X1 U15924 ( .IN1(\mem2[52][18] ), .IN2(n1101), .S(n8175), .Q(n10830) );
  MUX21X1 U15925 ( .IN1(\mem2[52][17] ), .IN2(n1079), .S(n8175), .Q(n10829) );
  MUX21X1 U15926 ( .IN1(\mem2[52][16] ), .IN2(n1057), .S(n8175), .Q(n10828) );
  AND2X1 U15927 ( .IN1(n8164), .IN2(n7122), .Q(n8175) );
  MUX21X1 U15928 ( .IN1(\mem2[51][23] ), .IN2(n1212), .S(n8176), .Q(n10827) );
  MUX21X1 U15929 ( .IN1(\mem2[51][22] ), .IN2(n1190), .S(n8176), .Q(n10826) );
  MUX21X1 U15930 ( .IN1(\mem2[51][21] ), .IN2(n1168), .S(n8176), .Q(n10825) );
  MUX21X1 U15931 ( .IN1(\mem2[51][20] ), .IN2(n1146), .S(n8176), .Q(n10824) );
  MUX21X1 U15932 ( .IN1(\mem2[51][19] ), .IN2(n1124), .S(n8176), .Q(n10823) );
  MUX21X1 U15933 ( .IN1(\mem2[51][18] ), .IN2(n1102), .S(n8176), .Q(n10822) );
  MUX21X1 U15934 ( .IN1(\mem2[51][17] ), .IN2(n1080), .S(n8176), .Q(n10821) );
  MUX21X1 U15935 ( .IN1(\mem2[51][16] ), .IN2(n1058), .S(n8176), .Q(n10820) );
  AND2X1 U15936 ( .IN1(n8164), .IN2(n7124), .Q(n8176) );
  MUX21X1 U15937 ( .IN1(\mem2[50][23] ), .IN2(n1212), .S(n8177), .Q(n10819) );
  MUX21X1 U15938 ( .IN1(\mem2[50][22] ), .IN2(n1190), .S(n8177), .Q(n10818) );
  MUX21X1 U15939 ( .IN1(\mem2[50][21] ), .IN2(n1168), .S(n8177), .Q(n10817) );
  MUX21X1 U15940 ( .IN1(\mem2[50][20] ), .IN2(n1146), .S(n8177), .Q(n10816) );
  MUX21X1 U15941 ( .IN1(\mem2[50][19] ), .IN2(n1124), .S(n8177), .Q(n10815) );
  MUX21X1 U15942 ( .IN1(\mem2[50][18] ), .IN2(n1102), .S(n8177), .Q(n10814) );
  MUX21X1 U15943 ( .IN1(\mem2[50][17] ), .IN2(n1080), .S(n8177), .Q(n10813) );
  MUX21X1 U15944 ( .IN1(\mem2[50][16] ), .IN2(n1058), .S(n8177), .Q(n10812) );
  AND2X1 U15945 ( .IN1(n8164), .IN2(n7126), .Q(n8177) );
  MUX21X1 U15946 ( .IN1(\mem2[49][23] ), .IN2(n1212), .S(n8178), .Q(n10811) );
  MUX21X1 U15947 ( .IN1(\mem2[49][22] ), .IN2(n1190), .S(n8178), .Q(n10810) );
  MUX21X1 U15948 ( .IN1(\mem2[49][21] ), .IN2(n1168), .S(n8178), .Q(n10809) );
  MUX21X1 U15949 ( .IN1(\mem2[49][20] ), .IN2(n1146), .S(n8178), .Q(n10808) );
  MUX21X1 U15950 ( .IN1(\mem2[49][19] ), .IN2(n1124), .S(n8178), .Q(n10807) );
  MUX21X1 U15951 ( .IN1(\mem2[49][18] ), .IN2(n1102), .S(n8178), .Q(n10806) );
  MUX21X1 U15952 ( .IN1(\mem2[49][17] ), .IN2(n1080), .S(n8178), .Q(n10805) );
  MUX21X1 U15953 ( .IN1(\mem2[49][16] ), .IN2(n1058), .S(n8178), .Q(n10804) );
  AND2X1 U15954 ( .IN1(n8164), .IN2(n7128), .Q(n8178) );
  MUX21X1 U15955 ( .IN1(\mem2[48][23] ), .IN2(n1212), .S(n8179), .Q(n10803) );
  MUX21X1 U15956 ( .IN1(\mem2[48][22] ), .IN2(n1190), .S(n8179), .Q(n10802) );
  MUX21X1 U15957 ( .IN1(\mem2[48][21] ), .IN2(n1168), .S(n8179), .Q(n10801) );
  MUX21X1 U15958 ( .IN1(\mem2[48][20] ), .IN2(n1146), .S(n8179), .Q(n10800) );
  MUX21X1 U15959 ( .IN1(\mem2[48][19] ), .IN2(n1124), .S(n8179), .Q(n10799) );
  MUX21X1 U15960 ( .IN1(\mem2[48][18] ), .IN2(n1102), .S(n8179), .Q(n10798) );
  MUX21X1 U15961 ( .IN1(\mem2[48][17] ), .IN2(n1080), .S(n8179), .Q(n10797) );
  MUX21X1 U15962 ( .IN1(\mem2[48][16] ), .IN2(n1058), .S(n8179), .Q(n10796) );
  AND2X1 U15963 ( .IN1(n8164), .IN2(n7130), .Q(n8179) );
  AND2X1 U15964 ( .IN1(n7966), .IN2(n7348), .Q(n8164) );
  AND2X1 U15965 ( .IN1(n8180), .IN2(n7968), .Q(n7348) );
  NOR2X0 U15966 ( .IN1(n8181), .IN2(n8182), .QN(n7968) );
  MUX21X1 U15967 ( .IN1(\mem2[47][23] ), .IN2(n1212), .S(n8183), .Q(n10795) );
  MUX21X1 U15968 ( .IN1(\mem2[47][22] ), .IN2(n1190), .S(n8183), .Q(n10794) );
  MUX21X1 U15969 ( .IN1(\mem2[47][21] ), .IN2(n1168), .S(n8183), .Q(n10793) );
  MUX21X1 U15970 ( .IN1(\mem2[47][20] ), .IN2(n1146), .S(n8183), .Q(n10792) );
  MUX21X1 U15971 ( .IN1(\mem2[47][19] ), .IN2(n1124), .S(n8183), .Q(n10791) );
  MUX21X1 U15972 ( .IN1(\mem2[47][18] ), .IN2(n1102), .S(n8183), .Q(n10790) );
  MUX21X1 U15973 ( .IN1(\mem2[47][17] ), .IN2(n1080), .S(n8183), .Q(n10789) );
  MUX21X1 U15974 ( .IN1(\mem2[47][16] ), .IN2(n1058), .S(n8183), .Q(n10788) );
  AND2X1 U15975 ( .IN1(n8184), .IN2(n7099), .Q(n8183) );
  MUX21X1 U15976 ( .IN1(\mem2[46][23] ), .IN2(n1212), .S(n8185), .Q(n10787) );
  MUX21X1 U15977 ( .IN1(\mem2[46][22] ), .IN2(n1190), .S(n8185), .Q(n10786) );
  MUX21X1 U15978 ( .IN1(\mem2[46][21] ), .IN2(n1168), .S(n8185), .Q(n10785) );
  MUX21X1 U15979 ( .IN1(\mem2[46][20] ), .IN2(n1146), .S(n8185), .Q(n10784) );
  MUX21X1 U15980 ( .IN1(\mem2[46][19] ), .IN2(n1124), .S(n8185), .Q(n10783) );
  MUX21X1 U15981 ( .IN1(\mem2[46][18] ), .IN2(n1102), .S(n8185), .Q(n10782) );
  MUX21X1 U15982 ( .IN1(\mem2[46][17] ), .IN2(n1080), .S(n8185), .Q(n10781) );
  MUX21X1 U15983 ( .IN1(\mem2[46][16] ), .IN2(n1058), .S(n8185), .Q(n10780) );
  AND2X1 U15984 ( .IN1(n8184), .IN2(n7102), .Q(n8185) );
  MUX21X1 U15985 ( .IN1(\mem2[45][23] ), .IN2(n1212), .S(n8186), .Q(n10779) );
  MUX21X1 U15986 ( .IN1(\mem2[45][22] ), .IN2(n1190), .S(n8186), .Q(n10778) );
  MUX21X1 U15987 ( .IN1(\mem2[45][21] ), .IN2(n1168), .S(n8186), .Q(n10777) );
  MUX21X1 U15988 ( .IN1(\mem2[45][20] ), .IN2(n1146), .S(n8186), .Q(n10776) );
  MUX21X1 U15989 ( .IN1(\mem2[45][19] ), .IN2(n1124), .S(n8186), .Q(n10775) );
  MUX21X1 U15990 ( .IN1(\mem2[45][18] ), .IN2(n1102), .S(n8186), .Q(n10774) );
  MUX21X1 U15991 ( .IN1(\mem2[45][17] ), .IN2(n1080), .S(n8186), .Q(n10773) );
  MUX21X1 U15992 ( .IN1(\mem2[45][16] ), .IN2(n1058), .S(n8186), .Q(n10772) );
  AND2X1 U15993 ( .IN1(n8184), .IN2(n7104), .Q(n8186) );
  MUX21X1 U15994 ( .IN1(\mem2[44][23] ), .IN2(n1212), .S(n8187), .Q(n10771) );
  MUX21X1 U15995 ( .IN1(\mem2[44][22] ), .IN2(n1190), .S(n8187), .Q(n10770) );
  MUX21X1 U15996 ( .IN1(\mem2[44][21] ), .IN2(n1168), .S(n8187), .Q(n10769) );
  MUX21X1 U15997 ( .IN1(\mem2[44][20] ), .IN2(n1146), .S(n8187), .Q(n10768) );
  MUX21X1 U15998 ( .IN1(\mem2[44][19] ), .IN2(n1124), .S(n8187), .Q(n10767) );
  MUX21X1 U15999 ( .IN1(\mem2[44][18] ), .IN2(n1102), .S(n8187), .Q(n10766) );
  MUX21X1 U16000 ( .IN1(\mem2[44][17] ), .IN2(n1080), .S(n8187), .Q(n10765) );
  MUX21X1 U16001 ( .IN1(\mem2[44][16] ), .IN2(n1058), .S(n8187), .Q(n10764) );
  AND2X1 U16002 ( .IN1(n8184), .IN2(n7106), .Q(n8187) );
  MUX21X1 U16003 ( .IN1(\mem2[43][23] ), .IN2(n1212), .S(n8188), .Q(n10763) );
  MUX21X1 U16004 ( .IN1(\mem2[43][22] ), .IN2(n1190), .S(n8188), .Q(n10762) );
  MUX21X1 U16005 ( .IN1(\mem2[43][21] ), .IN2(n1168), .S(n8188), .Q(n10761) );
  MUX21X1 U16006 ( .IN1(\mem2[43][20] ), .IN2(n1146), .S(n8188), .Q(n10760) );
  MUX21X1 U16007 ( .IN1(\mem2[43][19] ), .IN2(n1124), .S(n8188), .Q(n10759) );
  MUX21X1 U16008 ( .IN1(\mem2[43][18] ), .IN2(n1102), .S(n8188), .Q(n10758) );
  MUX21X1 U16009 ( .IN1(\mem2[43][17] ), .IN2(n1080), .S(n8188), .Q(n10757) );
  MUX21X1 U16010 ( .IN1(\mem2[43][16] ), .IN2(n1058), .S(n8188), .Q(n10756) );
  AND2X1 U16011 ( .IN1(n8184), .IN2(n7108), .Q(n8188) );
  MUX21X1 U16012 ( .IN1(\mem2[42][23] ), .IN2(n1212), .S(n8189), .Q(n10755) );
  MUX21X1 U16013 ( .IN1(\mem2[42][22] ), .IN2(n1190), .S(n8189), .Q(n10754) );
  MUX21X1 U16014 ( .IN1(\mem2[42][21] ), .IN2(n1168), .S(n8189), .Q(n10753) );
  MUX21X1 U16015 ( .IN1(\mem2[42][20] ), .IN2(n1146), .S(n8189), .Q(n10752) );
  MUX21X1 U16016 ( .IN1(\mem2[42][19] ), .IN2(n1124), .S(n8189), .Q(n10751) );
  MUX21X1 U16017 ( .IN1(\mem2[42][18] ), .IN2(n1102), .S(n8189), .Q(n10750) );
  MUX21X1 U16018 ( .IN1(\mem2[42][17] ), .IN2(n1080), .S(n8189), .Q(n10749) );
  MUX21X1 U16019 ( .IN1(\mem2[42][16] ), .IN2(n1058), .S(n8189), .Q(n10748) );
  AND2X1 U16020 ( .IN1(n8184), .IN2(n7110), .Q(n8189) );
  MUX21X1 U16021 ( .IN1(\mem2[41][23] ), .IN2(n1212), .S(n8190), .Q(n10747) );
  MUX21X1 U16022 ( .IN1(\mem2[41][22] ), .IN2(n1190), .S(n8190), .Q(n10746) );
  MUX21X1 U16023 ( .IN1(\mem2[41][21] ), .IN2(n1168), .S(n8190), .Q(n10745) );
  MUX21X1 U16024 ( .IN1(\mem2[41][20] ), .IN2(n1146), .S(n8190), .Q(n10744) );
  MUX21X1 U16025 ( .IN1(\mem2[41][19] ), .IN2(n1124), .S(n8190), .Q(n10743) );
  MUX21X1 U16026 ( .IN1(\mem2[41][18] ), .IN2(n1102), .S(n8190), .Q(n10742) );
  MUX21X1 U16027 ( .IN1(\mem2[41][17] ), .IN2(n1080), .S(n8190), .Q(n10741) );
  MUX21X1 U16028 ( .IN1(\mem2[41][16] ), .IN2(n1058), .S(n8190), .Q(n10740) );
  AND2X1 U16029 ( .IN1(n8184), .IN2(n7112), .Q(n8190) );
  MUX21X1 U16030 ( .IN1(\mem2[40][23] ), .IN2(n1212), .S(n8191), .Q(n10739) );
  MUX21X1 U16031 ( .IN1(\mem2[40][22] ), .IN2(n1190), .S(n8191), .Q(n10738) );
  MUX21X1 U16032 ( .IN1(\mem2[40][21] ), .IN2(n1168), .S(n8191), .Q(n10737) );
  MUX21X1 U16033 ( .IN1(\mem2[40][20] ), .IN2(n1146), .S(n8191), .Q(n10736) );
  MUX21X1 U16034 ( .IN1(\mem2[40][19] ), .IN2(n1124), .S(n8191), .Q(n10735) );
  MUX21X1 U16035 ( .IN1(\mem2[40][18] ), .IN2(n1102), .S(n8191), .Q(n10734) );
  MUX21X1 U16036 ( .IN1(\mem2[40][17] ), .IN2(n1080), .S(n8191), .Q(n10733) );
  MUX21X1 U16037 ( .IN1(\mem2[40][16] ), .IN2(n1058), .S(n8191), .Q(n10732) );
  AND2X1 U16038 ( .IN1(n8184), .IN2(n7114), .Q(n8191) );
  MUX21X1 U16039 ( .IN1(\mem2[39][23] ), .IN2(n1213), .S(n8192), .Q(n10731) );
  MUX21X1 U16040 ( .IN1(\mem2[39][22] ), .IN2(n1191), .S(n8192), .Q(n10730) );
  MUX21X1 U16041 ( .IN1(\mem2[39][21] ), .IN2(n1169), .S(n8192), .Q(n10729) );
  MUX21X1 U16042 ( .IN1(\mem2[39][20] ), .IN2(n1147), .S(n8192), .Q(n10728) );
  MUX21X1 U16043 ( .IN1(\mem2[39][19] ), .IN2(n1125), .S(n8192), .Q(n10727) );
  MUX21X1 U16044 ( .IN1(\mem2[39][18] ), .IN2(n1103), .S(n8192), .Q(n10726) );
  MUX21X1 U16045 ( .IN1(\mem2[39][17] ), .IN2(n1081), .S(n8192), .Q(n10725) );
  MUX21X1 U16046 ( .IN1(\mem2[39][16] ), .IN2(n1059), .S(n8192), .Q(n10724) );
  AND2X1 U16047 ( .IN1(n8184), .IN2(n7116), .Q(n8192) );
  MUX21X1 U16048 ( .IN1(\mem2[38][23] ), .IN2(n1213), .S(n8193), .Q(n10723) );
  MUX21X1 U16049 ( .IN1(\mem2[38][22] ), .IN2(n1191), .S(n8193), .Q(n10722) );
  MUX21X1 U16050 ( .IN1(\mem2[38][21] ), .IN2(n1169), .S(n8193), .Q(n10721) );
  MUX21X1 U16051 ( .IN1(\mem2[38][20] ), .IN2(n1147), .S(n8193), .Q(n10720) );
  MUX21X1 U16052 ( .IN1(\mem2[38][19] ), .IN2(n1125), .S(n8193), .Q(n10719) );
  MUX21X1 U16053 ( .IN1(\mem2[38][18] ), .IN2(n1103), .S(n8193), .Q(n10718) );
  MUX21X1 U16054 ( .IN1(\mem2[38][17] ), .IN2(n1081), .S(n8193), .Q(n10717) );
  MUX21X1 U16055 ( .IN1(\mem2[38][16] ), .IN2(n1059), .S(n8193), .Q(n10716) );
  AND2X1 U16056 ( .IN1(n8184), .IN2(n7118), .Q(n8193) );
  MUX21X1 U16057 ( .IN1(\mem2[37][23] ), .IN2(n1213), .S(n8194), .Q(n10715) );
  MUX21X1 U16058 ( .IN1(\mem2[37][22] ), .IN2(n1191), .S(n8194), .Q(n10714) );
  MUX21X1 U16059 ( .IN1(\mem2[37][21] ), .IN2(n1169), .S(n8194), .Q(n10713) );
  MUX21X1 U16060 ( .IN1(\mem2[37][20] ), .IN2(n1147), .S(n8194), .Q(n10712) );
  MUX21X1 U16061 ( .IN1(\mem2[37][19] ), .IN2(n1125), .S(n8194), .Q(n10711) );
  MUX21X1 U16062 ( .IN1(\mem2[37][18] ), .IN2(n1103), .S(n8194), .Q(n10710) );
  MUX21X1 U16063 ( .IN1(\mem2[37][17] ), .IN2(n1081), .S(n8194), .Q(n10709) );
  MUX21X1 U16064 ( .IN1(\mem2[37][16] ), .IN2(n1059), .S(n8194), .Q(n10708) );
  AND2X1 U16065 ( .IN1(n8184), .IN2(n7120), .Q(n8194) );
  MUX21X1 U16066 ( .IN1(\mem2[36][23] ), .IN2(n1213), .S(n8195), .Q(n10707) );
  MUX21X1 U16067 ( .IN1(\mem2[36][22] ), .IN2(n1191), .S(n8195), .Q(n10706) );
  MUX21X1 U16068 ( .IN1(\mem2[36][21] ), .IN2(n1169), .S(n8195), .Q(n10705) );
  MUX21X1 U16069 ( .IN1(\mem2[36][20] ), .IN2(n1147), .S(n8195), .Q(n10704) );
  MUX21X1 U16070 ( .IN1(\mem2[36][19] ), .IN2(n1125), .S(n8195), .Q(n10703) );
  MUX21X1 U16071 ( .IN1(\mem2[36][18] ), .IN2(n1103), .S(n8195), .Q(n10702) );
  MUX21X1 U16072 ( .IN1(\mem2[36][17] ), .IN2(n1081), .S(n8195), .Q(n10701) );
  MUX21X1 U16073 ( .IN1(\mem2[36][16] ), .IN2(n1059), .S(n8195), .Q(n10700) );
  AND2X1 U16074 ( .IN1(n8184), .IN2(n7122), .Q(n8195) );
  MUX21X1 U16075 ( .IN1(\mem2[35][23] ), .IN2(n1213), .S(n8196), .Q(n10699) );
  MUX21X1 U16076 ( .IN1(\mem2[35][22] ), .IN2(n1191), .S(n8196), .Q(n10698) );
  MUX21X1 U16077 ( .IN1(\mem2[35][21] ), .IN2(n1169), .S(n8196), .Q(n10697) );
  MUX21X1 U16078 ( .IN1(\mem2[35][20] ), .IN2(n1147), .S(n8196), .Q(n10696) );
  MUX21X1 U16079 ( .IN1(\mem2[35][19] ), .IN2(n1125), .S(n8196), .Q(n10695) );
  MUX21X1 U16080 ( .IN1(\mem2[35][18] ), .IN2(n1103), .S(n8196), .Q(n10694) );
  MUX21X1 U16081 ( .IN1(\mem2[35][17] ), .IN2(n1081), .S(n8196), .Q(n10693) );
  MUX21X1 U16082 ( .IN1(\mem2[35][16] ), .IN2(n1059), .S(n8196), .Q(n10692) );
  AND2X1 U16083 ( .IN1(n8184), .IN2(n7124), .Q(n8196) );
  MUX21X1 U16084 ( .IN1(\mem2[34][23] ), .IN2(n1213), .S(n8197), .Q(n10691) );
  MUX21X1 U16085 ( .IN1(\mem2[34][22] ), .IN2(n1191), .S(n8197), .Q(n10690) );
  MUX21X1 U16086 ( .IN1(\mem2[34][21] ), .IN2(n1169), .S(n8197), .Q(n10689) );
  MUX21X1 U16087 ( .IN1(\mem2[34][20] ), .IN2(n1147), .S(n8197), .Q(n10688) );
  MUX21X1 U16088 ( .IN1(\mem2[34][19] ), .IN2(n1125), .S(n8197), .Q(n10687) );
  MUX21X1 U16089 ( .IN1(\mem2[34][18] ), .IN2(n1103), .S(n8197), .Q(n10686) );
  MUX21X1 U16090 ( .IN1(\mem2[34][17] ), .IN2(n1081), .S(n8197), .Q(n10685) );
  MUX21X1 U16091 ( .IN1(\mem2[34][16] ), .IN2(n1059), .S(n8197), .Q(n10684) );
  AND2X1 U16092 ( .IN1(n8184), .IN2(n7126), .Q(n8197) );
  MUX21X1 U16093 ( .IN1(\mem2[33][23] ), .IN2(n1213), .S(n8198), .Q(n10683) );
  MUX21X1 U16094 ( .IN1(\mem2[33][22] ), .IN2(n1191), .S(n8198), .Q(n10682) );
  MUX21X1 U16095 ( .IN1(\mem2[33][21] ), .IN2(n1169), .S(n8198), .Q(n10681) );
  MUX21X1 U16096 ( .IN1(\mem2[33][20] ), .IN2(n1147), .S(n8198), .Q(n10680) );
  MUX21X1 U16097 ( .IN1(\mem2[33][19] ), .IN2(n1125), .S(n8198), .Q(n10679) );
  MUX21X1 U16098 ( .IN1(\mem2[33][18] ), .IN2(n1103), .S(n8198), .Q(n10678) );
  MUX21X1 U16099 ( .IN1(\mem2[33][17] ), .IN2(n1081), .S(n8198), .Q(n10677) );
  MUX21X1 U16100 ( .IN1(\mem2[33][16] ), .IN2(n1059), .S(n8198), .Q(n10676) );
  AND2X1 U16101 ( .IN1(n8184), .IN2(n7128), .Q(n8198) );
  MUX21X1 U16102 ( .IN1(\mem2[32][23] ), .IN2(n1213), .S(n8199), .Q(n10675) );
  MUX21X1 U16103 ( .IN1(\mem2[32][22] ), .IN2(n1191), .S(n8199), .Q(n10674) );
  MUX21X1 U16104 ( .IN1(\mem2[32][21] ), .IN2(n1169), .S(n8199), .Q(n10673) );
  MUX21X1 U16105 ( .IN1(\mem2[32][20] ), .IN2(n1147), .S(n8199), .Q(n10672) );
  MUX21X1 U16106 ( .IN1(\mem2[32][19] ), .IN2(n1125), .S(n8199), .Q(n10671) );
  MUX21X1 U16107 ( .IN1(\mem2[32][18] ), .IN2(n1103), .S(n8199), .Q(n10670) );
  MUX21X1 U16108 ( .IN1(\mem2[32][17] ), .IN2(n1081), .S(n8199), .Q(n10669) );
  MUX21X1 U16109 ( .IN1(\mem2[32][16] ), .IN2(n1059), .S(n8199), .Q(n10668) );
  AND2X1 U16110 ( .IN1(n8184), .IN2(n7130), .Q(n8199) );
  AND2X1 U16111 ( .IN1(n7966), .IN2(n7366), .Q(n8184) );
  AND2X1 U16112 ( .IN1(n8180), .IN2(n7986), .Q(n7366) );
  NOR2X0 U16113 ( .IN1(n8181), .IN2(addr[4]), .QN(n7986) );
  INVX0 U16114 ( .INP(addr[5]), .ZN(n8181) );
  MUX21X1 U16115 ( .IN1(\mem2[31][23] ), .IN2(n1213), .S(n8200), .Q(n10667) );
  MUX21X1 U16116 ( .IN1(\mem2[31][22] ), .IN2(n1191), .S(n8200), .Q(n10666) );
  MUX21X1 U16117 ( .IN1(\mem2[31][21] ), .IN2(n1169), .S(n8200), .Q(n10665) );
  MUX21X1 U16118 ( .IN1(\mem2[31][20] ), .IN2(n1147), .S(n8200), .Q(n10664) );
  MUX21X1 U16119 ( .IN1(\mem2[31][19] ), .IN2(n1125), .S(n8200), .Q(n10663) );
  MUX21X1 U16120 ( .IN1(\mem2[31][18] ), .IN2(n1103), .S(n8200), .Q(n10662) );
  MUX21X1 U16121 ( .IN1(\mem2[31][17] ), .IN2(n1081), .S(n8200), .Q(n10661) );
  MUX21X1 U16122 ( .IN1(\mem2[31][16] ), .IN2(n1059), .S(n8200), .Q(n10660) );
  AND2X1 U16123 ( .IN1(n8201), .IN2(n7099), .Q(n8200) );
  MUX21X1 U16124 ( .IN1(\mem2[30][23] ), .IN2(n1213), .S(n8202), .Q(n10659) );
  MUX21X1 U16125 ( .IN1(\mem2[30][22] ), .IN2(n1191), .S(n8202), .Q(n10658) );
  MUX21X1 U16126 ( .IN1(\mem2[30][21] ), .IN2(n1169), .S(n8202), .Q(n10657) );
  MUX21X1 U16127 ( .IN1(\mem2[30][20] ), .IN2(n1147), .S(n8202), .Q(n10656) );
  MUX21X1 U16128 ( .IN1(\mem2[30][19] ), .IN2(n1125), .S(n8202), .Q(n10655) );
  MUX21X1 U16129 ( .IN1(\mem2[30][18] ), .IN2(n1103), .S(n8202), .Q(n10654) );
  MUX21X1 U16130 ( .IN1(\mem2[30][17] ), .IN2(n1081), .S(n8202), .Q(n10653) );
  MUX21X1 U16131 ( .IN1(\mem2[30][16] ), .IN2(n1059), .S(n8202), .Q(n10652) );
  AND2X1 U16132 ( .IN1(n8201), .IN2(n7102), .Q(n8202) );
  MUX21X1 U16133 ( .IN1(\mem2[29][23] ), .IN2(n1213), .S(n8203), .Q(n10651) );
  MUX21X1 U16134 ( .IN1(\mem2[29][22] ), .IN2(n1191), .S(n8203), .Q(n10650) );
  MUX21X1 U16135 ( .IN1(\mem2[29][21] ), .IN2(n1169), .S(n8203), .Q(n10649) );
  MUX21X1 U16136 ( .IN1(\mem2[29][20] ), .IN2(n1147), .S(n8203), .Q(n10648) );
  MUX21X1 U16137 ( .IN1(\mem2[29][19] ), .IN2(n1125), .S(n8203), .Q(n10647) );
  MUX21X1 U16138 ( .IN1(\mem2[29][18] ), .IN2(n1103), .S(n8203), .Q(n10646) );
  MUX21X1 U16139 ( .IN1(\mem2[29][17] ), .IN2(n1081), .S(n8203), .Q(n10645) );
  MUX21X1 U16140 ( .IN1(\mem2[29][16] ), .IN2(n1059), .S(n8203), .Q(n10644) );
  AND2X1 U16141 ( .IN1(n8201), .IN2(n7104), .Q(n8203) );
  MUX21X1 U16142 ( .IN1(\mem2[28][23] ), .IN2(n1213), .S(n8204), .Q(n10643) );
  MUX21X1 U16143 ( .IN1(\mem2[28][22] ), .IN2(n1191), .S(n8204), .Q(n10642) );
  MUX21X1 U16144 ( .IN1(\mem2[28][21] ), .IN2(n1169), .S(n8204), .Q(n10641) );
  MUX21X1 U16145 ( .IN1(\mem2[28][20] ), .IN2(n1147), .S(n8204), .Q(n10640) );
  MUX21X1 U16146 ( .IN1(\mem2[28][19] ), .IN2(n1125), .S(n8204), .Q(n10639) );
  MUX21X1 U16147 ( .IN1(\mem2[28][18] ), .IN2(n1103), .S(n8204), .Q(n10638) );
  MUX21X1 U16148 ( .IN1(\mem2[28][17] ), .IN2(n1081), .S(n8204), .Q(n10637) );
  MUX21X1 U16149 ( .IN1(\mem2[28][16] ), .IN2(n1059), .S(n8204), .Q(n10636) );
  AND2X1 U16150 ( .IN1(n8201), .IN2(n7106), .Q(n8204) );
  MUX21X1 U16151 ( .IN1(\mem2[27][23] ), .IN2(n1214), .S(n8205), .Q(n10635) );
  MUX21X1 U16152 ( .IN1(\mem2[27][22] ), .IN2(n1192), .S(n8205), .Q(n10634) );
  MUX21X1 U16153 ( .IN1(\mem2[27][21] ), .IN2(n1170), .S(n8205), .Q(n10633) );
  MUX21X1 U16154 ( .IN1(\mem2[27][20] ), .IN2(n1148), .S(n8205), .Q(n10632) );
  MUX21X1 U16155 ( .IN1(\mem2[27][19] ), .IN2(n1126), .S(n8205), .Q(n10631) );
  MUX21X1 U16156 ( .IN1(\mem2[27][18] ), .IN2(n1104), .S(n8205), .Q(n10630) );
  MUX21X1 U16157 ( .IN1(\mem2[27][17] ), .IN2(n1082), .S(n8205), .Q(n10629) );
  MUX21X1 U16158 ( .IN1(\mem2[27][16] ), .IN2(n1060), .S(n8205), .Q(n10628) );
  AND2X1 U16159 ( .IN1(n8201), .IN2(n7108), .Q(n8205) );
  MUX21X1 U16160 ( .IN1(\mem2[26][23] ), .IN2(n1214), .S(n8206), .Q(n10627) );
  MUX21X1 U16161 ( .IN1(\mem2[26][22] ), .IN2(n1192), .S(n8206), .Q(n10626) );
  MUX21X1 U16162 ( .IN1(\mem2[26][21] ), .IN2(n1170), .S(n8206), .Q(n10625) );
  MUX21X1 U16163 ( .IN1(\mem2[26][20] ), .IN2(n1148), .S(n8206), .Q(n10624) );
  MUX21X1 U16164 ( .IN1(\mem2[26][19] ), .IN2(n1126), .S(n8206), .Q(n10623) );
  MUX21X1 U16165 ( .IN1(\mem2[26][18] ), .IN2(n1104), .S(n8206), .Q(n10622) );
  MUX21X1 U16166 ( .IN1(\mem2[26][17] ), .IN2(n1082), .S(n8206), .Q(n10621) );
  MUX21X1 U16167 ( .IN1(\mem2[26][16] ), .IN2(n1060), .S(n8206), .Q(n10620) );
  AND2X1 U16168 ( .IN1(n8201), .IN2(n7110), .Q(n8206) );
  MUX21X1 U16169 ( .IN1(\mem2[25][23] ), .IN2(n1214), .S(n8207), .Q(n10619) );
  MUX21X1 U16170 ( .IN1(\mem2[25][22] ), .IN2(n1192), .S(n8207), .Q(n10618) );
  MUX21X1 U16171 ( .IN1(\mem2[25][21] ), .IN2(n1170), .S(n8207), .Q(n10617) );
  MUX21X1 U16172 ( .IN1(\mem2[25][20] ), .IN2(n1148), .S(n8207), .Q(n10616) );
  MUX21X1 U16173 ( .IN1(\mem2[25][19] ), .IN2(n1126), .S(n8207), .Q(n10615) );
  MUX21X1 U16174 ( .IN1(\mem2[25][18] ), .IN2(n1104), .S(n8207), .Q(n10614) );
  MUX21X1 U16175 ( .IN1(\mem2[25][17] ), .IN2(n1082), .S(n8207), .Q(n10613) );
  MUX21X1 U16176 ( .IN1(\mem2[25][16] ), .IN2(n1060), .S(n8207), .Q(n10612) );
  AND2X1 U16177 ( .IN1(n8201), .IN2(n7112), .Q(n8207) );
  MUX21X1 U16178 ( .IN1(\mem2[24][23] ), .IN2(n1214), .S(n8208), .Q(n10611) );
  MUX21X1 U16179 ( .IN1(\mem2[24][22] ), .IN2(n1192), .S(n8208), .Q(n10610) );
  MUX21X1 U16180 ( .IN1(\mem2[24][21] ), .IN2(n1170), .S(n8208), .Q(n10609) );
  MUX21X1 U16181 ( .IN1(\mem2[24][20] ), .IN2(n1148), .S(n8208), .Q(n10608) );
  MUX21X1 U16182 ( .IN1(\mem2[24][19] ), .IN2(n1126), .S(n8208), .Q(n10607) );
  MUX21X1 U16183 ( .IN1(\mem2[24][18] ), .IN2(n1104), .S(n8208), .Q(n10606) );
  MUX21X1 U16184 ( .IN1(\mem2[24][17] ), .IN2(n1082), .S(n8208), .Q(n10605) );
  MUX21X1 U16185 ( .IN1(\mem2[24][16] ), .IN2(n1060), .S(n8208), .Q(n10604) );
  AND2X1 U16186 ( .IN1(n8201), .IN2(n7114), .Q(n8208) );
  MUX21X1 U16187 ( .IN1(\mem2[23][23] ), .IN2(n1214), .S(n8209), .Q(n10603) );
  MUX21X1 U16188 ( .IN1(\mem2[23][22] ), .IN2(n1192), .S(n8209), .Q(n10602) );
  MUX21X1 U16189 ( .IN1(\mem2[23][21] ), .IN2(n1170), .S(n8209), .Q(n10601) );
  MUX21X1 U16190 ( .IN1(\mem2[23][20] ), .IN2(n1148), .S(n8209), .Q(n10600) );
  MUX21X1 U16191 ( .IN1(\mem2[23][19] ), .IN2(n1126), .S(n8209), .Q(n10599) );
  MUX21X1 U16192 ( .IN1(\mem2[23][18] ), .IN2(n1104), .S(n8209), .Q(n10598) );
  MUX21X1 U16193 ( .IN1(\mem2[23][17] ), .IN2(n1082), .S(n8209), .Q(n10597) );
  MUX21X1 U16194 ( .IN1(\mem2[23][16] ), .IN2(n1060), .S(n8209), .Q(n10596) );
  AND2X1 U16195 ( .IN1(n8201), .IN2(n7116), .Q(n8209) );
  MUX21X1 U16196 ( .IN1(\mem2[22][23] ), .IN2(n1214), .S(n8210), .Q(n10595) );
  MUX21X1 U16197 ( .IN1(\mem2[22][22] ), .IN2(n1192), .S(n8210), .Q(n10594) );
  MUX21X1 U16198 ( .IN1(\mem2[22][21] ), .IN2(n1170), .S(n8210), .Q(n10593) );
  MUX21X1 U16199 ( .IN1(\mem2[22][20] ), .IN2(n1148), .S(n8210), .Q(n10592) );
  MUX21X1 U16200 ( .IN1(\mem2[22][19] ), .IN2(n1126), .S(n8210), .Q(n10591) );
  MUX21X1 U16201 ( .IN1(\mem2[22][18] ), .IN2(n1104), .S(n8210), .Q(n10590) );
  MUX21X1 U16202 ( .IN1(\mem2[22][17] ), .IN2(n1082), .S(n8210), .Q(n10589) );
  MUX21X1 U16203 ( .IN1(\mem2[22][16] ), .IN2(n1060), .S(n8210), .Q(n10588) );
  AND2X1 U16204 ( .IN1(n8201), .IN2(n7118), .Q(n8210) );
  MUX21X1 U16205 ( .IN1(\mem2[21][23] ), .IN2(n1214), .S(n8211), .Q(n10587) );
  MUX21X1 U16206 ( .IN1(\mem2[21][22] ), .IN2(n1192), .S(n8211), .Q(n10586) );
  MUX21X1 U16207 ( .IN1(\mem2[21][21] ), .IN2(n1170), .S(n8211), .Q(n10585) );
  MUX21X1 U16208 ( .IN1(\mem2[21][20] ), .IN2(n1148), .S(n8211), .Q(n10584) );
  MUX21X1 U16209 ( .IN1(\mem2[21][19] ), .IN2(n1126), .S(n8211), .Q(n10583) );
  MUX21X1 U16210 ( .IN1(\mem2[21][18] ), .IN2(n1104), .S(n8211), .Q(n10582) );
  MUX21X1 U16211 ( .IN1(\mem2[21][17] ), .IN2(n1082), .S(n8211), .Q(n10581) );
  MUX21X1 U16212 ( .IN1(\mem2[21][16] ), .IN2(n1060), .S(n8211), .Q(n10580) );
  AND2X1 U16213 ( .IN1(n8201), .IN2(n7120), .Q(n8211) );
  MUX21X1 U16214 ( .IN1(\mem2[20][23] ), .IN2(n1214), .S(n8212), .Q(n10579) );
  MUX21X1 U16215 ( .IN1(\mem2[20][22] ), .IN2(n1192), .S(n8212), .Q(n10578) );
  MUX21X1 U16216 ( .IN1(\mem2[20][21] ), .IN2(n1170), .S(n8212), .Q(n10577) );
  MUX21X1 U16217 ( .IN1(\mem2[20][20] ), .IN2(n1148), .S(n8212), .Q(n10576) );
  MUX21X1 U16218 ( .IN1(\mem2[20][19] ), .IN2(n1126), .S(n8212), .Q(n10575) );
  MUX21X1 U16219 ( .IN1(\mem2[20][18] ), .IN2(n1104), .S(n8212), .Q(n10574) );
  MUX21X1 U16220 ( .IN1(\mem2[20][17] ), .IN2(n1082), .S(n8212), .Q(n10573) );
  MUX21X1 U16221 ( .IN1(\mem2[20][16] ), .IN2(n1060), .S(n8212), .Q(n10572) );
  AND2X1 U16222 ( .IN1(n8201), .IN2(n7122), .Q(n8212) );
  MUX21X1 U16223 ( .IN1(\mem2[19][23] ), .IN2(n1214), .S(n8213), .Q(n10571) );
  MUX21X1 U16224 ( .IN1(\mem2[19][22] ), .IN2(n1192), .S(n8213), .Q(n10570) );
  MUX21X1 U16225 ( .IN1(\mem2[19][21] ), .IN2(n1170), .S(n8213), .Q(n10569) );
  MUX21X1 U16226 ( .IN1(\mem2[19][20] ), .IN2(n1148), .S(n8213), .Q(n10568) );
  MUX21X1 U16227 ( .IN1(\mem2[19][19] ), .IN2(n1126), .S(n8213), .Q(n10567) );
  MUX21X1 U16228 ( .IN1(\mem2[19][18] ), .IN2(n1104), .S(n8213), .Q(n10566) );
  MUX21X1 U16229 ( .IN1(\mem2[19][17] ), .IN2(n1082), .S(n8213), .Q(n10565) );
  MUX21X1 U16230 ( .IN1(\mem2[19][16] ), .IN2(n1060), .S(n8213), .Q(n10564) );
  AND2X1 U16231 ( .IN1(n8201), .IN2(n7124), .Q(n8213) );
  MUX21X1 U16232 ( .IN1(\mem2[18][23] ), .IN2(n1214), .S(n8214), .Q(n10563) );
  MUX21X1 U16233 ( .IN1(\mem2[18][22] ), .IN2(n1192), .S(n8214), .Q(n10562) );
  MUX21X1 U16234 ( .IN1(\mem2[18][21] ), .IN2(n1170), .S(n8214), .Q(n10561) );
  MUX21X1 U16235 ( .IN1(\mem2[18][20] ), .IN2(n1148), .S(n8214), .Q(n10560) );
  MUX21X1 U16236 ( .IN1(\mem2[18][19] ), .IN2(n1126), .S(n8214), .Q(n10559) );
  MUX21X1 U16237 ( .IN1(\mem2[18][18] ), .IN2(n1104), .S(n8214), .Q(n10558) );
  MUX21X1 U16238 ( .IN1(\mem2[18][17] ), .IN2(n1082), .S(n8214), .Q(n10557) );
  MUX21X1 U16239 ( .IN1(\mem2[18][16] ), .IN2(n1060), .S(n8214), .Q(n10556) );
  AND2X1 U16240 ( .IN1(n8201), .IN2(n7126), .Q(n8214) );
  MUX21X1 U16241 ( .IN1(\mem2[17][23] ), .IN2(n1214), .S(n8215), .Q(n10555) );
  MUX21X1 U16242 ( .IN1(\mem2[17][22] ), .IN2(n1192), .S(n8215), .Q(n10554) );
  MUX21X1 U16243 ( .IN1(\mem2[17][21] ), .IN2(n1170), .S(n8215), .Q(n10553) );
  MUX21X1 U16244 ( .IN1(\mem2[17][20] ), .IN2(n1148), .S(n8215), .Q(n10552) );
  MUX21X1 U16245 ( .IN1(\mem2[17][19] ), .IN2(n1126), .S(n8215), .Q(n10551) );
  MUX21X1 U16246 ( .IN1(\mem2[17][18] ), .IN2(n1104), .S(n8215), .Q(n10550) );
  MUX21X1 U16247 ( .IN1(\mem2[17][17] ), .IN2(n1082), .S(n8215), .Q(n10549) );
  MUX21X1 U16248 ( .IN1(\mem2[17][16] ), .IN2(n1060), .S(n8215), .Q(n10548) );
  AND2X1 U16249 ( .IN1(n8201), .IN2(n7128), .Q(n8215) );
  MUX21X1 U16250 ( .IN1(\mem2[16][23] ), .IN2(n1214), .S(n8216), .Q(n10547) );
  MUX21X1 U16251 ( .IN1(\mem2[16][22] ), .IN2(n1192), .S(n8216), .Q(n10546) );
  MUX21X1 U16252 ( .IN1(\mem2[16][21] ), .IN2(n1170), .S(n8216), .Q(n10545) );
  MUX21X1 U16253 ( .IN1(\mem2[16][20] ), .IN2(n1148), .S(n8216), .Q(n10544) );
  MUX21X1 U16254 ( .IN1(\mem2[16][19] ), .IN2(n1126), .S(n8216), .Q(n10543) );
  MUX21X1 U16255 ( .IN1(\mem2[16][18] ), .IN2(n1104), .S(n8216), .Q(n10542) );
  MUX21X1 U16256 ( .IN1(\mem2[16][17] ), .IN2(n1082), .S(n8216), .Q(n10541) );
  MUX21X1 U16257 ( .IN1(\mem2[16][16] ), .IN2(n1060), .S(n8216), .Q(n10540) );
  AND2X1 U16258 ( .IN1(n8201), .IN2(n7130), .Q(n8216) );
  AND2X1 U16259 ( .IN1(n7966), .IN2(n7384), .Q(n8201) );
  AND2X1 U16260 ( .IN1(n8180), .IN2(n8004), .Q(n7384) );
  NOR2X0 U16261 ( .IN1(n8182), .IN2(addr[5]), .QN(n8004) );
  INVX0 U16262 ( .INP(addr[4]), .ZN(n8182) );
  MUX21X1 U16263 ( .IN1(\mem2[15][23] ), .IN2(n1215), .S(n8217), .Q(n10539) );
  MUX21X1 U16264 ( .IN1(\mem2[15][22] ), .IN2(n1193), .S(n8217), .Q(n10538) );
  MUX21X1 U16265 ( .IN1(\mem2[15][21] ), .IN2(n1171), .S(n8217), .Q(n10537) );
  MUX21X1 U16266 ( .IN1(\mem2[15][20] ), .IN2(n1149), .S(n8217), .Q(n10536) );
  MUX21X1 U16267 ( .IN1(\mem2[15][19] ), .IN2(n1127), .S(n8217), .Q(n10535) );
  MUX21X1 U16268 ( .IN1(\mem2[15][18] ), .IN2(n1105), .S(n8217), .Q(n10534) );
  MUX21X1 U16269 ( .IN1(\mem2[15][17] ), .IN2(n1083), .S(n8217), .Q(n10533) );
  MUX21X1 U16270 ( .IN1(\mem2[15][16] ), .IN2(n1061), .S(n8217), .Q(n10532) );
  AND2X1 U16271 ( .IN1(n8218), .IN2(n7099), .Q(n8217) );
  AND2X1 U16272 ( .IN1(n8219), .IN2(n8220), .Q(n7099) );
  MUX21X1 U16273 ( .IN1(\mem2[14][23] ), .IN2(n1215), .S(n8221), .Q(n10531) );
  MUX21X1 U16274 ( .IN1(\mem2[14][22] ), .IN2(n1193), .S(n8221), .Q(n10530) );
  MUX21X1 U16275 ( .IN1(\mem2[14][21] ), .IN2(n1171), .S(n8221), .Q(n10529) );
  MUX21X1 U16276 ( .IN1(\mem2[14][20] ), .IN2(n1149), .S(n8221), .Q(n10528) );
  MUX21X1 U16277 ( .IN1(\mem2[14][19] ), .IN2(n1127), .S(n8221), .Q(n10527) );
  MUX21X1 U16278 ( .IN1(\mem2[14][18] ), .IN2(n1105), .S(n8221), .Q(n10526) );
  MUX21X1 U16279 ( .IN1(\mem2[14][17] ), .IN2(n1083), .S(n8221), .Q(n10525) );
  MUX21X1 U16280 ( .IN1(\mem2[14][16] ), .IN2(n1061), .S(n8221), .Q(n10524) );
  AND2X1 U16281 ( .IN1(n8218), .IN2(n7102), .Q(n8221) );
  AND2X1 U16282 ( .IN1(n8222), .IN2(n8219), .Q(n7102) );
  MUX21X1 U16283 ( .IN1(\mem2[13][23] ), .IN2(n1215), .S(n8223), .Q(n10523) );
  MUX21X1 U16284 ( .IN1(\mem2[13][22] ), .IN2(n1193), .S(n8223), .Q(n10522) );
  MUX21X1 U16285 ( .IN1(\mem2[13][21] ), .IN2(n1171), .S(n8223), .Q(n10521) );
  MUX21X1 U16286 ( .IN1(\mem2[13][20] ), .IN2(n1149), .S(n8223), .Q(n10520) );
  MUX21X1 U16287 ( .IN1(\mem2[13][19] ), .IN2(n1127), .S(n8223), .Q(n10519) );
  MUX21X1 U16288 ( .IN1(\mem2[13][18] ), .IN2(n1105), .S(n8223), .Q(n10518) );
  MUX21X1 U16289 ( .IN1(\mem2[13][17] ), .IN2(n1083), .S(n8223), .Q(n10517) );
  MUX21X1 U16290 ( .IN1(\mem2[13][16] ), .IN2(n1061), .S(n8223), .Q(n10516) );
  AND2X1 U16291 ( .IN1(n8218), .IN2(n7104), .Q(n8223) );
  AND2X1 U16292 ( .IN1(n8224), .IN2(n8219), .Q(n7104) );
  MUX21X1 U16293 ( .IN1(\mem2[12][23] ), .IN2(n1215), .S(n8225), .Q(n10515) );
  MUX21X1 U16294 ( .IN1(\mem2[12][22] ), .IN2(n1193), .S(n8225), .Q(n10514) );
  MUX21X1 U16295 ( .IN1(\mem2[12][21] ), .IN2(n1171), .S(n8225), .Q(n10513) );
  MUX21X1 U16296 ( .IN1(\mem2[12][20] ), .IN2(n1149), .S(n8225), .Q(n10512) );
  MUX21X1 U16297 ( .IN1(\mem2[12][19] ), .IN2(n1127), .S(n8225), .Q(n10511) );
  MUX21X1 U16298 ( .IN1(\mem2[12][18] ), .IN2(n1105), .S(n8225), .Q(n10510) );
  MUX21X1 U16299 ( .IN1(\mem2[12][17] ), .IN2(n1083), .S(n8225), .Q(n10509) );
  MUX21X1 U16300 ( .IN1(\mem2[12][16] ), .IN2(n1061), .S(n8225), .Q(n10508) );
  AND2X1 U16301 ( .IN1(n8218), .IN2(n7106), .Q(n8225) );
  AND2X1 U16302 ( .IN1(n8226), .IN2(n8219), .Q(n7106) );
  NOR2X0 U16303 ( .IN1(n8227), .IN2(n8228), .QN(n8219) );
  MUX21X1 U16304 ( .IN1(\mem2[11][23] ), .IN2(n1215), .S(n8229), .Q(n10507) );
  MUX21X1 U16305 ( .IN1(\mem2[11][22] ), .IN2(n1193), .S(n8229), .Q(n10506) );
  MUX21X1 U16306 ( .IN1(\mem2[11][21] ), .IN2(n1171), .S(n8229), .Q(n10505) );
  MUX21X1 U16307 ( .IN1(\mem2[11][20] ), .IN2(n1149), .S(n8229), .Q(n10504) );
  MUX21X1 U16308 ( .IN1(\mem2[11][19] ), .IN2(n1127), .S(n8229), .Q(n10503) );
  MUX21X1 U16309 ( .IN1(\mem2[11][18] ), .IN2(n1105), .S(n8229), .Q(n10502) );
  MUX21X1 U16310 ( .IN1(\mem2[11][17] ), .IN2(n1083), .S(n8229), .Q(n10501) );
  MUX21X1 U16311 ( .IN1(\mem2[11][16] ), .IN2(n1061), .S(n8229), .Q(n10500) );
  AND2X1 U16312 ( .IN1(n8218), .IN2(n7108), .Q(n8229) );
  AND2X1 U16313 ( .IN1(n8230), .IN2(n8220), .Q(n7108) );
  MUX21X1 U16314 ( .IN1(\mem2[10][23] ), .IN2(n1215), .S(n8231), .Q(n10499) );
  MUX21X1 U16315 ( .IN1(\mem2[10][22] ), .IN2(n1193), .S(n8231), .Q(n10498) );
  MUX21X1 U16316 ( .IN1(\mem2[10][21] ), .IN2(n1171), .S(n8231), .Q(n10497) );
  MUX21X1 U16317 ( .IN1(\mem2[10][20] ), .IN2(n1149), .S(n8231), .Q(n10496) );
  MUX21X1 U16318 ( .IN1(\mem2[10][19] ), .IN2(n1127), .S(n8231), .Q(n10495) );
  MUX21X1 U16319 ( .IN1(\mem2[10][18] ), .IN2(n1105), .S(n8231), .Q(n10494) );
  MUX21X1 U16320 ( .IN1(\mem2[10][17] ), .IN2(n1083), .S(n8231), .Q(n10493) );
  MUX21X1 U16321 ( .IN1(\mem2[10][16] ), .IN2(n1061), .S(n8231), .Q(n10492) );
  AND2X1 U16322 ( .IN1(n8218), .IN2(n7110), .Q(n8231) );
  AND2X1 U16323 ( .IN1(n8230), .IN2(n8222), .Q(n7110) );
  MUX21X1 U16324 ( .IN1(\mem2[9][23] ), .IN2(n1215), .S(n8232), .Q(n10491) );
  MUX21X1 U16325 ( .IN1(\mem2[9][22] ), .IN2(n1193), .S(n8232), .Q(n10490) );
  MUX21X1 U16326 ( .IN1(\mem2[9][21] ), .IN2(n1171), .S(n8232), .Q(n10489) );
  MUX21X1 U16327 ( .IN1(\mem2[9][20] ), .IN2(n1149), .S(n8232), .Q(n10488) );
  MUX21X1 U16328 ( .IN1(\mem2[9][19] ), .IN2(n1127), .S(n8232), .Q(n10487) );
  MUX21X1 U16329 ( .IN1(\mem2[9][18] ), .IN2(n1105), .S(n8232), .Q(n10486) );
  MUX21X1 U16330 ( .IN1(\mem2[9][17] ), .IN2(n1083), .S(n8232), .Q(n10485) );
  MUX21X1 U16331 ( .IN1(\mem2[9][16] ), .IN2(n1061), .S(n8232), .Q(n10484) );
  AND2X1 U16332 ( .IN1(n8218), .IN2(n7112), .Q(n8232) );
  AND2X1 U16333 ( .IN1(n8230), .IN2(n8224), .Q(n7112) );
  MUX21X1 U16334 ( .IN1(\mem2[8][23] ), .IN2(n1215), .S(n8233), .Q(n10483) );
  MUX21X1 U16335 ( .IN1(\mem2[8][22] ), .IN2(n1193), .S(n8233), .Q(n10482) );
  MUX21X1 U16336 ( .IN1(\mem2[8][21] ), .IN2(n1171), .S(n8233), .Q(n10481) );
  MUX21X1 U16337 ( .IN1(\mem2[8][20] ), .IN2(n1149), .S(n8233), .Q(n10480) );
  MUX21X1 U16338 ( .IN1(\mem2[8][19] ), .IN2(n1127), .S(n8233), .Q(n10479) );
  MUX21X1 U16339 ( .IN1(\mem2[8][18] ), .IN2(n1105), .S(n8233), .Q(n10478) );
  MUX21X1 U16340 ( .IN1(\mem2[8][17] ), .IN2(n1083), .S(n8233), .Q(n10477) );
  MUX21X1 U16341 ( .IN1(\mem2[8][16] ), .IN2(n1061), .S(n8233), .Q(n10476) );
  AND2X1 U16342 ( .IN1(n8218), .IN2(n7114), .Q(n8233) );
  AND2X1 U16343 ( .IN1(n8230), .IN2(n8226), .Q(n7114) );
  NOR2X0 U16344 ( .IN1(n8227), .IN2(addr[2]), .QN(n8230) );
  INVX0 U16345 ( .INP(addr[3]), .ZN(n8227) );
  MUX21X1 U16346 ( .IN1(\mem2[7][23] ), .IN2(n1215), .S(n8234), .Q(n10475) );
  MUX21X1 U16347 ( .IN1(\mem2[7][22] ), .IN2(n1193), .S(n8234), .Q(n10474) );
  MUX21X1 U16348 ( .IN1(\mem2[7][21] ), .IN2(n1171), .S(n8234), .Q(n10473) );
  MUX21X1 U16349 ( .IN1(\mem2[7][20] ), .IN2(n1149), .S(n8234), .Q(n10472) );
  MUX21X1 U16350 ( .IN1(\mem2[7][19] ), .IN2(n1127), .S(n8234), .Q(n10471) );
  MUX21X1 U16351 ( .IN1(\mem2[7][18] ), .IN2(n1105), .S(n8234), .Q(n10470) );
  MUX21X1 U16352 ( .IN1(\mem2[7][17] ), .IN2(n1083), .S(n8234), .Q(n10469) );
  MUX21X1 U16353 ( .IN1(\mem2[7][16] ), .IN2(n1061), .S(n8234), .Q(n10468) );
  AND2X1 U16354 ( .IN1(n8218), .IN2(n7116), .Q(n8234) );
  AND2X1 U16355 ( .IN1(n8235), .IN2(n8220), .Q(n7116) );
  MUX21X1 U16356 ( .IN1(\mem2[6][23] ), .IN2(n1215), .S(n8236), .Q(n10467) );
  MUX21X1 U16357 ( .IN1(\mem2[6][22] ), .IN2(n1193), .S(n8236), .Q(n10466) );
  MUX21X1 U16358 ( .IN1(\mem2[6][21] ), .IN2(n1171), .S(n8236), .Q(n10465) );
  MUX21X1 U16359 ( .IN1(\mem2[6][20] ), .IN2(n1149), .S(n8236), .Q(n10464) );
  MUX21X1 U16360 ( .IN1(\mem2[6][19] ), .IN2(n1127), .S(n8236), .Q(n10463) );
  MUX21X1 U16361 ( .IN1(\mem2[6][18] ), .IN2(n1105), .S(n8236), .Q(n10462) );
  MUX21X1 U16362 ( .IN1(\mem2[6][17] ), .IN2(n1083), .S(n8236), .Q(n10461) );
  MUX21X1 U16363 ( .IN1(\mem2[6][16] ), .IN2(n1061), .S(n8236), .Q(n10460) );
  AND2X1 U16364 ( .IN1(n8218), .IN2(n7118), .Q(n8236) );
  AND2X1 U16365 ( .IN1(n8235), .IN2(n8222), .Q(n7118) );
  MUX21X1 U16366 ( .IN1(\mem2[5][23] ), .IN2(n1215), .S(n8237), .Q(n10459) );
  MUX21X1 U16367 ( .IN1(\mem2[5][22] ), .IN2(n1193), .S(n8237), .Q(n10458) );
  MUX21X1 U16368 ( .IN1(\mem2[5][21] ), .IN2(n1171), .S(n8237), .Q(n10457) );
  MUX21X1 U16369 ( .IN1(\mem2[5][20] ), .IN2(n1149), .S(n8237), .Q(n10456) );
  MUX21X1 U16370 ( .IN1(\mem2[5][19] ), .IN2(n1127), .S(n8237), .Q(n10455) );
  MUX21X1 U16371 ( .IN1(\mem2[5][18] ), .IN2(n1105), .S(n8237), .Q(n10454) );
  MUX21X1 U16372 ( .IN1(\mem2[5][17] ), .IN2(n1083), .S(n8237), .Q(n10453) );
  MUX21X1 U16373 ( .IN1(\mem2[5][16] ), .IN2(n1061), .S(n8237), .Q(n10452) );
  AND2X1 U16374 ( .IN1(n8218), .IN2(n7120), .Q(n8237) );
  AND2X1 U16375 ( .IN1(n8235), .IN2(n8224), .Q(n7120) );
  MUX21X1 U16376 ( .IN1(\mem2[4][23] ), .IN2(n1215), .S(n8238), .Q(n10451) );
  MUX21X1 U16377 ( .IN1(\mem2[4][22] ), .IN2(n1193), .S(n8238), .Q(n10450) );
  MUX21X1 U16378 ( .IN1(\mem2[4][21] ), .IN2(n1171), .S(n8238), .Q(n10449) );
  MUX21X1 U16379 ( .IN1(\mem2[4][20] ), .IN2(n1149), .S(n8238), .Q(n10448) );
  MUX21X1 U16380 ( .IN1(\mem2[4][19] ), .IN2(n1127), .S(n8238), .Q(n10447) );
  MUX21X1 U16381 ( .IN1(\mem2[4][18] ), .IN2(n1105), .S(n8238), .Q(n10446) );
  MUX21X1 U16382 ( .IN1(\mem2[4][17] ), .IN2(n1083), .S(n8238), .Q(n10445) );
  MUX21X1 U16383 ( .IN1(\mem2[4][16] ), .IN2(n1061), .S(n8238), .Q(n10444) );
  AND2X1 U16384 ( .IN1(n8218), .IN2(n7122), .Q(n8238) );
  AND2X1 U16385 ( .IN1(n8235), .IN2(n8226), .Q(n7122) );
  NOR2X0 U16386 ( .IN1(n8228), .IN2(addr[3]), .QN(n8235) );
  INVX0 U16387 ( .INP(addr[2]), .ZN(n8228) );
  MUX21X1 U16388 ( .IN1(\mem2[3][23] ), .IN2(n1216), .S(n8239), .Q(n10443) );
  MUX21X1 U16389 ( .IN1(\mem2[3][22] ), .IN2(n1194), .S(n8239), .Q(n10442) );
  MUX21X1 U16390 ( .IN1(\mem2[3][21] ), .IN2(n1172), .S(n8239), .Q(n10441) );
  MUX21X1 U16391 ( .IN1(\mem2[3][20] ), .IN2(n1150), .S(n8239), .Q(n10440) );
  MUX21X1 U16392 ( .IN1(\mem2[3][19] ), .IN2(n1128), .S(n8239), .Q(n10439) );
  MUX21X1 U16393 ( .IN1(\mem2[3][18] ), .IN2(n1106), .S(n8239), .Q(n10438) );
  MUX21X1 U16394 ( .IN1(\mem2[3][17] ), .IN2(n1084), .S(n8239), .Q(n10437) );
  MUX21X1 U16395 ( .IN1(\mem2[3][16] ), .IN2(n1062), .S(n8239), .Q(n10436) );
  AND2X1 U16396 ( .IN1(n8218), .IN2(n7124), .Q(n8239) );
  AND2X1 U16397 ( .IN1(n8240), .IN2(n8220), .Q(n7124) );
  NOR2X0 U16398 ( .IN1(n8241), .IN2(n8242), .QN(n8220) );
  MUX21X1 U16399 ( .IN1(\mem2[2][23] ), .IN2(n1216), .S(n8243), .Q(n10435) );
  MUX21X1 U16400 ( .IN1(\mem2[2][22] ), .IN2(n1194), .S(n8243), .Q(n10434) );
  MUX21X1 U16401 ( .IN1(\mem2[2][21] ), .IN2(n1172), .S(n8243), .Q(n10433) );
  MUX21X1 U16402 ( .IN1(\mem2[2][20] ), .IN2(n1150), .S(n8243), .Q(n10432) );
  MUX21X1 U16403 ( .IN1(\mem2[2][19] ), .IN2(n1128), .S(n8243), .Q(n10431) );
  MUX21X1 U16404 ( .IN1(\mem2[2][18] ), .IN2(n1106), .S(n8243), .Q(n10430) );
  MUX21X1 U16405 ( .IN1(\mem2[2][17] ), .IN2(n1084), .S(n8243), .Q(n10429) );
  MUX21X1 U16406 ( .IN1(\mem2[2][16] ), .IN2(n1062), .S(n8243), .Q(n10428) );
  AND2X1 U16407 ( .IN1(n8218), .IN2(n7126), .Q(n8243) );
  AND2X1 U16408 ( .IN1(n8240), .IN2(n8222), .Q(n7126) );
  NOR2X0 U16409 ( .IN1(n8241), .IN2(addr[0]), .QN(n8222) );
  INVX0 U16410 ( .INP(addr[1]), .ZN(n8241) );
  MUX21X1 U16411 ( .IN1(\mem2[1][23] ), .IN2(n1216), .S(n8244), .Q(n10427) );
  MUX21X1 U16412 ( .IN1(\mem2[1][22] ), .IN2(n1194), .S(n8244), .Q(n10426) );
  MUX21X1 U16413 ( .IN1(\mem2[1][21] ), .IN2(n1172), .S(n8244), .Q(n10425) );
  MUX21X1 U16414 ( .IN1(\mem2[1][20] ), .IN2(n1150), .S(n8244), .Q(n10424) );
  MUX21X1 U16415 ( .IN1(\mem2[1][19] ), .IN2(n1128), .S(n8244), .Q(n10423) );
  MUX21X1 U16416 ( .IN1(\mem2[1][18] ), .IN2(n1106), .S(n8244), .Q(n10422) );
  MUX21X1 U16417 ( .IN1(\mem2[1][17] ), .IN2(n1084), .S(n8244), .Q(n10421) );
  MUX21X1 U16418 ( .IN1(\mem2[1][16] ), .IN2(n1062), .S(n8244), .Q(n10420) );
  AND2X1 U16419 ( .IN1(n8218), .IN2(n7128), .Q(n8244) );
  AND2X1 U16420 ( .IN1(n8240), .IN2(n8224), .Q(n7128) );
  NOR2X0 U16421 ( .IN1(n8242), .IN2(addr[1]), .QN(n8224) );
  INVX0 U16422 ( .INP(addr[0]), .ZN(n8242) );
  MUX21X1 U16423 ( .IN1(\mem2[0][23] ), .IN2(n1216), .S(n8245), .Q(n10419) );
  MUX21X1 U16424 ( .IN1(\mem2[0][22] ), .IN2(n1194), .S(n8245), .Q(n10418) );
  MUX21X1 U16425 ( .IN1(\mem2[0][21] ), .IN2(n1172), .S(n8245), .Q(n10417) );
  MUX21X1 U16426 ( .IN1(\mem2[0][20] ), .IN2(n1150), .S(n8245), .Q(n10416) );
  MUX21X1 U16427 ( .IN1(\mem2[0][19] ), .IN2(n1128), .S(n8245), .Q(n10415) );
  MUX21X1 U16428 ( .IN1(\mem2[0][18] ), .IN2(n1106), .S(n8245), .Q(n10414) );
  MUX21X1 U16429 ( .IN1(\mem2[0][17] ), .IN2(n1084), .S(n8245), .Q(n10413) );
  MUX21X1 U16430 ( .IN1(\mem2[0][16] ), .IN2(n1062), .S(n8245), .Q(n10412) );
  AND2X1 U16431 ( .IN1(n8218), .IN2(n7130), .Q(n8245) );
  AND2X1 U16432 ( .IN1(n8240), .IN2(n8226), .Q(n7130) );
  NOR2X0 U16433 ( .IN1(addr[0]), .IN2(addr[1]), .QN(n8226) );
  NOR2X0 U16434 ( .IN1(addr[2]), .IN2(addr[3]), .QN(n8240) );
  AND2X1 U16435 ( .IN1(n7966), .IN2(n7402), .Q(n8218) );
  AND2X1 U16436 ( .IN1(n8180), .IN2(n8022), .Q(n7402) );
  NOR2X0 U16437 ( .IN1(addr[4]), .IN2(addr[5]), .QN(n8022) );
  NOR2X0 U16438 ( .IN1(addr[6]), .IN2(addr[7]), .QN(n8180) );
  AND2X1 U16439 ( .IN1(we[2]), .IN2(ce), .Q(n7966) );
  MUX21X1 U16440 ( .IN1(N61), .IN2(addr[7]), .S(ce), .Q(n10411) );
  MUX21X1 U16441 ( .IN1(N60), .IN2(addr[6]), .S(ce), .Q(n10409) );
  MUX21X1 U16442 ( .IN1(N59), .IN2(addr[5]), .S(ce), .Q(n10407) );
  MUX21X1 U16443 ( .IN1(N58), .IN2(addr[4]), .S(ce), .Q(n10405) );
  MUX21X1 U16444 ( .IN1(N57), .IN2(addr[3]), .S(ce), .Q(n10403) );
  MUX21X1 U16445 ( .IN1(N56), .IN2(addr[2]), .S(ce), .Q(n10401) );
  MUX21X1 U16446 ( .IN1(N55), .IN2(addr[1]), .S(ce), .Q(n10399) );
  MUX21X1 U16447 ( .IN1(N54), .IN2(addr[0]), .S(ce), .Q(n10397) );
endmodule


module eth_fifo_DATA_WIDTH32_DEPTH16_CNT_WIDTH5_test_0 ( data_in, data_out, 
        clk, reset, write, read, clear, almost_full, full, almost_empty, empty, 
        cnt, eth_top_test_point_11887_in, test_si, test_so, test_se );
  input [31:0] data_in;
  output [31:0] data_out;
  output [4:0] cnt;
  input clk, reset, write, read, clear, eth_top_test_point_11887_in, test_si,
         test_se;
  output almost_full, full, almost_empty, empty, test_so;
  wire   N15, N16, N17, \fifo[0][31] , \fifo[0][30] , \fifo[0][29] ,
         \fifo[0][28] , \fifo[0][27] , \fifo[0][26] , \fifo[0][25] ,
         \fifo[0][24] , \fifo[0][23] , \fifo[0][22] , \fifo[0][21] ,
         \fifo[0][20] , \fifo[0][19] , \fifo[0][18] , \fifo[0][17] ,
         \fifo[0][16] , \fifo[0][15] , \fifo[0][14] , \fifo[0][13] ,
         \fifo[0][12] , \fifo[0][11] , \fifo[0][10] , \fifo[0][9] ,
         \fifo[0][8] , \fifo[0][7] , \fifo[0][6] , \fifo[0][5] , \fifo[0][4] ,
         \fifo[0][3] , \fifo[0][2] , \fifo[0][1] , \fifo[0][0] , \fifo[1][31] ,
         \fifo[1][30] , \fifo[1][29] , \fifo[1][28] , \fifo[1][27] ,
         \fifo[1][26] , \fifo[1][25] , \fifo[1][24] , \fifo[1][23] ,
         \fifo[1][22] , \fifo[1][21] , \fifo[1][20] , \fifo[1][19] ,
         \fifo[1][18] , \fifo[1][17] , \fifo[1][16] , \fifo[1][15] ,
         \fifo[1][14] , \fifo[1][13] , \fifo[1][12] , \fifo[1][11] ,
         \fifo[1][10] , \fifo[1][9] , \fifo[1][8] , \fifo[1][7] , \fifo[1][6] ,
         \fifo[1][5] , \fifo[1][4] , \fifo[1][3] , \fifo[1][2] , \fifo[1][1] ,
         \fifo[1][0] , \fifo[2][31] , \fifo[2][30] , \fifo[2][29] ,
         \fifo[2][28] , \fifo[2][27] , \fifo[2][26] , \fifo[2][25] ,
         \fifo[2][24] , \fifo[2][23] , \fifo[2][22] , \fifo[2][21] ,
         \fifo[2][20] , \fifo[2][19] , \fifo[2][18] , \fifo[2][17] ,
         \fifo[2][16] , \fifo[2][15] , \fifo[2][14] , \fifo[2][13] ,
         \fifo[2][12] , \fifo[2][11] , \fifo[2][10] , \fifo[2][9] ,
         \fifo[2][8] , \fifo[2][7] , \fifo[2][6] , \fifo[2][5] , \fifo[2][4] ,
         \fifo[2][3] , \fifo[2][2] , \fifo[2][1] , \fifo[2][0] , \fifo[3][31] ,
         \fifo[3][30] , \fifo[3][29] , \fifo[3][28] , \fifo[3][27] ,
         \fifo[3][26] , \fifo[3][25] , \fifo[3][24] , \fifo[3][23] ,
         \fifo[3][22] , \fifo[3][21] , \fifo[3][20] , \fifo[3][19] ,
         \fifo[3][18] , \fifo[3][17] , \fifo[3][16] , \fifo[3][15] ,
         \fifo[3][14] , \fifo[3][13] , \fifo[3][12] , \fifo[3][11] ,
         \fifo[3][10] , \fifo[3][9] , \fifo[3][8] , \fifo[3][7] , \fifo[3][6] ,
         \fifo[3][5] , \fifo[3][4] , \fifo[3][3] , \fifo[3][2] , \fifo[3][1] ,
         \fifo[3][0] , \fifo[4][31] , \fifo[4][30] , \fifo[4][29] ,
         \fifo[4][28] , \fifo[4][27] , \fifo[4][26] , \fifo[4][25] ,
         \fifo[4][24] , \fifo[4][23] , \fifo[4][22] , \fifo[4][21] ,
         \fifo[4][20] , \fifo[4][19] , \fifo[4][18] , \fifo[4][17] ,
         \fifo[4][16] , \fifo[4][15] , \fifo[4][14] , \fifo[4][13] ,
         \fifo[4][12] , \fifo[4][11] , \fifo[4][10] , \fifo[4][9] ,
         \fifo[4][8] , \fifo[4][7] , \fifo[4][6] , \fifo[4][5] , \fifo[4][4] ,
         \fifo[4][3] , \fifo[4][2] , \fifo[4][1] , \fifo[4][0] , \fifo[5][31] ,
         \fifo[5][30] , \fifo[5][29] , \fifo[5][28] , \fifo[5][27] ,
         \fifo[5][26] , \fifo[5][25] , \fifo[5][24] , \fifo[5][23] ,
         \fifo[5][22] , \fifo[5][21] , \fifo[5][20] , \fifo[5][19] ,
         \fifo[5][18] , \fifo[5][17] , \fifo[5][16] , \fifo[5][15] ,
         \fifo[5][14] , \fifo[5][13] , \fifo[5][12] , \fifo[5][11] ,
         \fifo[5][10] , \fifo[5][9] , \fifo[5][8] , \fifo[5][7] , \fifo[5][6] ,
         \fifo[5][5] , \fifo[5][4] , \fifo[5][3] , \fifo[5][2] , \fifo[5][1] ,
         \fifo[5][0] , \fifo[6][31] , \fifo[6][30] , \fifo[6][29] ,
         \fifo[6][28] , \fifo[6][27] , \fifo[6][26] , \fifo[6][25] ,
         \fifo[6][24] , \fifo[6][23] , \fifo[6][22] , \fifo[6][21] ,
         \fifo[6][20] , \fifo[6][19] , \fifo[6][18] , \fifo[6][17] ,
         \fifo[6][16] , \fifo[6][15] , \fifo[6][14] , \fifo[6][13] ,
         \fifo[6][12] , \fifo[6][11] , \fifo[6][10] , \fifo[6][9] ,
         \fifo[6][8] , \fifo[6][7] , \fifo[6][6] , \fifo[6][5] , \fifo[6][4] ,
         \fifo[6][3] , \fifo[6][2] , \fifo[6][1] , \fifo[6][0] , \fifo[7][31] ,
         \fifo[7][30] , \fifo[7][29] , \fifo[7][28] , \fifo[7][27] ,
         \fifo[7][26] , \fifo[7][25] , \fifo[7][24] , \fifo[7][23] ,
         \fifo[7][22] , \fifo[7][21] , \fifo[7][20] , \fifo[7][19] ,
         \fifo[7][18] , \fifo[7][17] , \fifo[7][16] , \fifo[7][15] ,
         \fifo[7][14] , \fifo[7][13] , \fifo[7][12] , \fifo[7][11] ,
         \fifo[7][10] , \fifo[7][9] , \fifo[7][8] , \fifo[7][7] , \fifo[7][6] ,
         \fifo[7][5] , \fifo[7][4] , \fifo[7][3] , \fifo[7][2] , \fifo[7][1] ,
         \fifo[7][0] , \fifo[8][31] , \fifo[8][30] , \fifo[8][29] ,
         \fifo[8][28] , \fifo[8][27] , \fifo[8][26] , \fifo[8][25] ,
         \fifo[8][24] , \fifo[8][23] , \fifo[8][22] , \fifo[8][21] ,
         \fifo[8][20] , \fifo[8][19] , \fifo[8][18] , \fifo[8][17] ,
         \fifo[8][16] , \fifo[8][15] , \fifo[8][14] , \fifo[8][13] ,
         \fifo[8][12] , \fifo[8][11] , \fifo[8][10] , \fifo[8][9] ,
         \fifo[8][8] , \fifo[8][7] , \fifo[8][6] , \fifo[8][5] , \fifo[8][4] ,
         \fifo[8][3] , \fifo[8][2] , \fifo[8][1] , \fifo[8][0] , \fifo[9][31] ,
         \fifo[9][30] , \fifo[9][29] , \fifo[9][28] , \fifo[9][27] ,
         \fifo[9][26] , \fifo[9][25] , \fifo[9][24] , \fifo[9][23] ,
         \fifo[9][22] , \fifo[9][21] , \fifo[9][20] , \fifo[9][19] ,
         \fifo[9][18] , \fifo[9][17] , \fifo[9][16] , \fifo[9][15] ,
         \fifo[9][14] , \fifo[9][13] , \fifo[9][12] , \fifo[9][11] ,
         \fifo[9][10] , \fifo[9][9] , \fifo[9][8] , \fifo[9][7] , \fifo[9][6] ,
         \fifo[9][5] , \fifo[9][4] , \fifo[9][3] , \fifo[9][2] , \fifo[9][1] ,
         \fifo[9][0] , \fifo[10][31] , \fifo[10][30] , \fifo[10][29] ,
         \fifo[10][28] , \fifo[10][27] , \fifo[10][26] , \fifo[10][25] ,
         \fifo[10][24] , \fifo[10][23] , \fifo[10][22] , \fifo[10][21] ,
         \fifo[10][20] , \fifo[10][19] , \fifo[10][18] , \fifo[10][17] ,
         \fifo[10][16] , \fifo[10][15] , \fifo[10][14] , \fifo[10][13] ,
         \fifo[10][12] , \fifo[10][11] , \fifo[10][10] , \fifo[10][9] ,
         \fifo[10][8] , \fifo[10][7] , \fifo[10][6] , \fifo[10][5] ,
         \fifo[10][4] , \fifo[10][3] , \fifo[10][2] , \fifo[10][1] ,
         \fifo[10][0] , \fifo[11][31] , \fifo[11][30] , \fifo[11][29] ,
         \fifo[11][28] , \fifo[11][27] , \fifo[11][26] , \fifo[11][25] ,
         \fifo[11][24] , \fifo[11][23] , \fifo[11][22] , \fifo[11][21] ,
         \fifo[11][20] , \fifo[11][19] , \fifo[11][18] , \fifo[11][17] ,
         \fifo[11][16] , \fifo[11][15] , \fifo[11][14] , \fifo[11][13] ,
         \fifo[11][12] , \fifo[11][11] , \fifo[11][10] , \fifo[11][9] ,
         \fifo[11][8] , \fifo[11][7] , \fifo[11][6] , \fifo[11][5] ,
         \fifo[11][4] , \fifo[11][3] , \fifo[11][2] , \fifo[11][1] ,
         \fifo[11][0] , \fifo[12][31] , \fifo[12][30] , \fifo[12][29] ,
         \fifo[12][28] , \fifo[12][27] , \fifo[12][26] , \fifo[12][25] ,
         \fifo[12][24] , \fifo[12][23] , \fifo[12][22] , \fifo[12][21] ,
         \fifo[12][20] , \fifo[12][19] , \fifo[12][18] , \fifo[12][17] ,
         \fifo[12][16] , \fifo[12][15] , \fifo[12][14] , \fifo[12][13] ,
         \fifo[12][12] , \fifo[12][11] , \fifo[12][10] , \fifo[12][9] ,
         \fifo[12][8] , \fifo[12][7] , \fifo[12][6] , \fifo[12][5] ,
         \fifo[12][4] , \fifo[12][3] , \fifo[12][2] , \fifo[12][1] ,
         \fifo[12][0] , \fifo[13][31] , \fifo[13][30] , \fifo[13][29] ,
         \fifo[13][28] , \fifo[13][27] , \fifo[13][26] , \fifo[13][25] ,
         \fifo[13][24] , \fifo[13][23] , \fifo[13][22] , \fifo[13][21] ,
         \fifo[13][20] , \fifo[13][19] , \fifo[13][18] , \fifo[13][17] ,
         \fifo[13][16] , \fifo[13][15] , \fifo[13][14] , \fifo[13][13] ,
         \fifo[13][12] , \fifo[13][11] , \fifo[13][10] , \fifo[13][9] ,
         \fifo[13][8] , \fifo[13][7] , \fifo[13][6] , \fifo[13][5] ,
         \fifo[13][4] , \fifo[13][3] , \fifo[13][2] , \fifo[13][1] ,
         \fifo[13][0] , \fifo[14][31] , \fifo[14][30] , \fifo[14][29] ,
         \fifo[14][28] , \fifo[14][27] , \fifo[14][26] , \fifo[14][25] ,
         \fifo[14][24] , \fifo[14][23] , \fifo[14][22] , \fifo[14][21] ,
         \fifo[14][20] , \fifo[14][19] , \fifo[14][18] , \fifo[14][17] ,
         \fifo[14][16] , \fifo[14][15] , \fifo[14][14] , \fifo[14][13] ,
         \fifo[14][12] , \fifo[14][11] , \fifo[14][10] , \fifo[14][9] ,
         \fifo[14][8] , \fifo[14][7] , \fifo[14][6] , \fifo[14][5] ,
         \fifo[14][4] , \fifo[14][3] , \fifo[14][2] , \fifo[14][1] ,
         \fifo[14][0] , \fifo[15][31] , \fifo[15][30] , \fifo[15][29] ,
         \fifo[15][28] , \fifo[15][27] , \fifo[15][26] , \fifo[15][25] ,
         \fifo[15][24] , \fifo[15][23] , \fifo[15][22] , \fifo[15][21] ,
         \fifo[15][20] , \fifo[15][19] , \fifo[15][18] , \fifo[15][17] ,
         \fifo[15][16] , \fifo[15][15] , \fifo[15][14] , \fifo[15][13] ,
         \fifo[15][12] , \fifo[15][11] , \fifo[15][10] , \fifo[15][9] ,
         \fifo[15][8] , \fifo[15][7] , \fifo[15][6] , \fifo[15][5] ,
         \fifo[15][4] , \fifo[15][3] , \fifo[15][2] , \fifo[15][1] ,
         \fifo[15][0] , N124, N125, N126, N127, N128, N129, N130, N131, N132,
         N133, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, \U3/U1/Z_0 , n564, n584, n585, n586, n587, n588, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n2, n1311, n1312, n1313, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n428;
  wire   [3:0] write_pointer;
  assign test_so = write_pointer[3];
  assign \U3/U1/Z_0  = read;

  SDFFARX1 \cnt_reg[0]  ( .D(n1162), .SI(test_si), .SE(test_se), .CLK(n6), 
        .RSTB(n428), .Q(cnt[0]), .QN(n1311) );
  SDFFARX1 \cnt_reg[1]  ( .D(n1161), .SI(cnt[0]), .SE(test_se), .CLK(n5), 
        .RSTB(n428), .Q(cnt[1]), .QN(n584) );
  SDFFARX1 \cnt_reg[2]  ( .D(n1160), .SI(cnt[1]), .SE(test_se), .CLK(n5), 
        .RSTB(n428), .Q(cnt[2]), .QN(n1312) );
  SDFFARX1 \cnt_reg[3]  ( .D(n1159), .SI(cnt[2]), .SE(test_se), .CLK(n5), 
        .RSTB(n428), .Q(cnt[3]), .QN(n1313) );
  SDFFARX1 \cnt_reg[4]  ( .D(n1158), .SI(cnt[3]), .SE(test_se), .CLK(n5), 
        .RSTB(n428), .Q(cnt[4]), .QN(n564) );
  SDFFARX1 \read_pointer_reg[0]  ( .D(n1157), .SI(\fifo[15][31] ), .SE(test_se), .CLK(n5), .RSTB(n428), .Q(n2), .QN(n588) );
  SDFFARX1 \read_pointer_reg[1]  ( .D(n1156), .SI(n2), .SE(test_se), .CLK(n5), 
        .RSTB(n428), .Q(N15), .QN(n587) );
  SDFFARX1 \read_pointer_reg[2]  ( .D(n1155), .SI(N15), .SE(test_se), .CLK(n5), 
        .RSTB(n428), .Q(N16), .QN(n586) );
  SDFFARX1 \read_pointer_reg[3]  ( .D(n1154), .SI(N16), .SE(test_se), .CLK(n5), 
        .RSTB(n428), .Q(N17), .QN(n585) );
  SDFFARX1 \write_pointer_reg[0]  ( .D(n1153), .SI(N17), .SE(test_se), .CLK(n5), .RSTB(n428), .Q(write_pointer[0]) );
  SDFFARX1 \write_pointer_reg[1]  ( .D(n1152), .SI(write_pointer[0]), .SE(
        test_se), .CLK(n5), .RSTB(n428), .Q(write_pointer[1]), .QN(n4) );
  SDFFARX1 \write_pointer_reg[2]  ( .D(n1151), .SI(write_pointer[1]), .SE(
        test_se), .CLK(n5), .RSTB(n428), .Q(write_pointer[2]), .QN(n1) );
  SDFFARX1 \write_pointer_reg[3]  ( .D(n1150), .SI(write_pointer[2]), .SE(
        test_se), .CLK(n5), .RSTB(n428), .Q(write_pointer[3]), .QN(n3) );
  SDFFX1 \fifo_reg[0][31]  ( .D(n1149), .SI(\fifo[0][30] ), .SE(test_se), 
        .CLK(n20), .Q(\fifo[0][31] ), .QN(n1939) );
  SDFFX1 \fifo_reg[0][30]  ( .D(n1148), .SI(\fifo[0][29] ), .SE(test_se), 
        .CLK(n20), .Q(\fifo[0][30] ), .QN(n1940) );
  SDFFX1 \fifo_reg[0][29]  ( .D(n1147), .SI(\fifo[0][28] ), .SE(test_se), 
        .CLK(n20), .Q(\fifo[0][29] ), .QN(n1941) );
  SDFFX1 \fifo_reg[0][28]  ( .D(n1146), .SI(\fifo[0][27] ), .SE(test_se), 
        .CLK(n19), .Q(\fifo[0][28] ), .QN(n1942) );
  SDFFX1 \fifo_reg[0][27]  ( .D(n1145), .SI(\fifo[0][26] ), .SE(test_se), 
        .CLK(n19), .Q(\fifo[0][27] ), .QN(n1943) );
  SDFFX1 \fifo_reg[0][26]  ( .D(n1144), .SI(\fifo[0][25] ), .SE(test_se), 
        .CLK(n19), .Q(\fifo[0][26] ), .QN(n1944) );
  SDFFX1 \fifo_reg[0][25]  ( .D(n1143), .SI(\fifo[0][24] ), .SE(test_se), 
        .CLK(n19), .Q(\fifo[0][25] ), .QN(n1945) );
  SDFFX1 \fifo_reg[0][24]  ( .D(n1142), .SI(\fifo[0][23] ), .SE(test_se), 
        .CLK(n19), .Q(\fifo[0][24] ), .QN(n1946) );
  SDFFX1 \fifo_reg[0][23]  ( .D(n1141), .SI(\fifo[0][22] ), .SE(test_se), 
        .CLK(n19), .Q(\fifo[0][23] ), .QN(n1947) );
  SDFFX1 \fifo_reg[0][22]  ( .D(n1140), .SI(\fifo[0][21] ), .SE(test_se), 
        .CLK(n19), .Q(\fifo[0][22] ), .QN(n1948) );
  SDFFX1 \fifo_reg[0][21]  ( .D(n1139), .SI(\fifo[0][20] ), .SE(test_se), 
        .CLK(n19), .Q(\fifo[0][21] ), .QN(n1949) );
  SDFFX1 \fifo_reg[0][20]  ( .D(n1138), .SI(\fifo[0][19] ), .SE(test_se), 
        .CLK(n19), .Q(\fifo[0][20] ), .QN(n1950) );
  SDFFX1 \fifo_reg[0][19]  ( .D(n1137), .SI(\fifo[0][18] ), .SE(test_se), 
        .CLK(n19), .Q(\fifo[0][19] ), .QN(n1951) );
  SDFFX1 \fifo_reg[0][18]  ( .D(n1136), .SI(\fifo[0][17] ), .SE(test_se), 
        .CLK(n19), .Q(\fifo[0][18] ), .QN(n1952) );
  SDFFX1 \fifo_reg[0][17]  ( .D(n1135), .SI(\fifo[0][16] ), .SE(test_se), 
        .CLK(n19), .Q(\fifo[0][17] ), .QN(n1953) );
  SDFFX1 \fifo_reg[0][16]  ( .D(n1134), .SI(\fifo[0][15] ), .SE(test_se), 
        .CLK(n19), .Q(\fifo[0][16] ), .QN(n1954) );
  SDFFX1 \fifo_reg[0][15]  ( .D(n1133), .SI(\fifo[0][14] ), .SE(test_se), 
        .CLK(n19), .Q(\fifo[0][15] ), .QN(n1955) );
  SDFFX1 \fifo_reg[0][14]  ( .D(n1132), .SI(\fifo[0][13] ), .SE(test_se), 
        .CLK(n18), .Q(\fifo[0][14] ), .QN(n1956) );
  SDFFX1 \fifo_reg[0][13]  ( .D(n1131), .SI(\fifo[0][12] ), .SE(test_se), 
        .CLK(n18), .Q(\fifo[0][13] ), .QN(n1957) );
  SDFFX1 \fifo_reg[0][12]  ( .D(n1130), .SI(\fifo[0][11] ), .SE(test_se), 
        .CLK(n18), .Q(\fifo[0][12] ), .QN(n1958) );
  SDFFX1 \fifo_reg[0][11]  ( .D(n1129), .SI(\fifo[0][10] ), .SE(test_se), 
        .CLK(n18), .Q(\fifo[0][11] ), .QN(n1959) );
  SDFFX1 \fifo_reg[0][10]  ( .D(n1128), .SI(\fifo[0][9] ), .SE(test_se), .CLK(
        n18), .Q(\fifo[0][10] ), .QN(n1960) );
  SDFFX1 \fifo_reg[0][9]  ( .D(n1127), .SI(\fifo[0][8] ), .SE(test_se), .CLK(
        n18), .Q(\fifo[0][9] ), .QN(n1961) );
  SDFFX1 \fifo_reg[0][8]  ( .D(n1126), .SI(\fifo[0][7] ), .SE(test_se), .CLK(
        n18), .Q(\fifo[0][8] ), .QN(n1962) );
  SDFFX1 \fifo_reg[0][7]  ( .D(n1125), .SI(\fifo[0][6] ), .SE(test_se), .CLK(
        n18), .Q(\fifo[0][7] ), .QN(n1963) );
  SDFFX1 \fifo_reg[0][6]  ( .D(n1124), .SI(\fifo[0][5] ), .SE(test_se), .CLK(
        n18), .Q(\fifo[0][6] ), .QN(n1964) );
  SDFFX1 \fifo_reg[0][5]  ( .D(n1123), .SI(\fifo[0][4] ), .SE(test_se), .CLK(
        n18), .Q(\fifo[0][5] ), .QN(n1965) );
  SDFFX1 \fifo_reg[0][4]  ( .D(n1122), .SI(\fifo[0][3] ), .SE(test_se), .CLK(
        n18), .Q(\fifo[0][4] ), .QN(n1966) );
  SDFFX1 \fifo_reg[0][3]  ( .D(n1121), .SI(\fifo[0][2] ), .SE(test_se), .CLK(
        n18), .Q(\fifo[0][3] ), .QN(n1967) );
  SDFFX1 \fifo_reg[0][2]  ( .D(n1120), .SI(\fifo[0][1] ), .SE(test_se), .CLK(
        n18), .Q(\fifo[0][2] ), .QN(n1968) );
  SDFFX1 \fifo_reg[0][1]  ( .D(n1119), .SI(\fifo[0][0] ), .SE(test_se), .CLK(
        n18), .Q(\fifo[0][1] ), .QN(n1969) );
  SDFFX1 \fifo_reg[0][0]  ( .D(n1118), .SI(data_out[31]), .SE(test_se), .CLK(
        n17), .Q(\fifo[0][0] ), .QN(n1970) );
  SDFFX1 \fifo_reg[1][31]  ( .D(n1117), .SI(\fifo[1][30] ), .SE(test_se), 
        .CLK(n22), .Q(\fifo[1][31] ), .QN(n1821) );
  SDFFX1 \fifo_reg[1][30]  ( .D(n1116), .SI(\fifo[1][29] ), .SE(test_se), 
        .CLK(n22), .Q(\fifo[1][30] ), .QN(n1822) );
  SDFFX1 \fifo_reg[1][29]  ( .D(n1115), .SI(\fifo[1][28] ), .SE(test_se), 
        .CLK(n22), .Q(\fifo[1][29] ), .QN(n1823) );
  SDFFX1 \fifo_reg[1][28]  ( .D(n1114), .SI(\fifo[1][27] ), .SE(test_se), 
        .CLK(n22), .Q(\fifo[1][28] ), .QN(n1824) );
  SDFFX1 \fifo_reg[1][27]  ( .D(n1113), .SI(\fifo[1][26] ), .SE(test_se), 
        .CLK(n22), .Q(\fifo[1][27] ), .QN(n1825) );
  SDFFX1 \fifo_reg[1][26]  ( .D(n1112), .SI(\fifo[1][25] ), .SE(test_se), 
        .CLK(n22), .Q(\fifo[1][26] ), .QN(n1826) );
  SDFFX1 \fifo_reg[1][25]  ( .D(n1111), .SI(\fifo[1][24] ), .SE(test_se), 
        .CLK(n22), .Q(\fifo[1][25] ), .QN(n1827) );
  SDFFX1 \fifo_reg[1][24]  ( .D(n1110), .SI(\fifo[1][23] ), .SE(test_se), 
        .CLK(n22), .Q(\fifo[1][24] ), .QN(n1828) );
  SDFFX1 \fifo_reg[1][23]  ( .D(n1109), .SI(\fifo[1][22] ), .SE(test_se), 
        .CLK(n21), .Q(\fifo[1][23] ), .QN(n1829) );
  SDFFX1 \fifo_reg[1][22]  ( .D(n1108), .SI(\fifo[1][21] ), .SE(test_se), 
        .CLK(n21), .Q(\fifo[1][22] ), .QN(n1830) );
  SDFFX1 \fifo_reg[1][21]  ( .D(n1107), .SI(\fifo[1][20] ), .SE(test_se), 
        .CLK(n21), .Q(\fifo[1][21] ), .QN(n1831) );
  SDFFX1 \fifo_reg[1][20]  ( .D(n1106), .SI(\fifo[1][19] ), .SE(test_se), 
        .CLK(n21), .Q(\fifo[1][20] ), .QN(n1832) );
  SDFFX1 \fifo_reg[1][19]  ( .D(n1105), .SI(\fifo[1][18] ), .SE(test_se), 
        .CLK(n21), .Q(\fifo[1][19] ), .QN(n1833) );
  SDFFX1 \fifo_reg[1][18]  ( .D(n1104), .SI(\fifo[1][17] ), .SE(test_se), 
        .CLK(n21), .Q(\fifo[1][18] ), .QN(n1834) );
  SDFFX1 \fifo_reg[1][17]  ( .D(n1103), .SI(\fifo[1][16] ), .SE(test_se), 
        .CLK(n21), .Q(\fifo[1][17] ), .QN(n1835) );
  SDFFX1 \fifo_reg[1][16]  ( .D(n1102), .SI(\fifo[1][15] ), .SE(test_se), 
        .CLK(n21), .Q(\fifo[1][16] ), .QN(n1836) );
  SDFFX1 \fifo_reg[1][15]  ( .D(n1101), .SI(\fifo[1][14] ), .SE(test_se), 
        .CLK(n21), .Q(\fifo[1][15] ), .QN(n1837) );
  SDFFX1 \fifo_reg[1][14]  ( .D(n1100), .SI(\fifo[1][13] ), .SE(test_se), 
        .CLK(n21), .Q(\fifo[1][14] ), .QN(n1838) );
  SDFFX1 \fifo_reg[1][13]  ( .D(n1099), .SI(\fifo[1][12] ), .SE(test_se), 
        .CLK(n21), .Q(\fifo[1][13] ), .QN(n1839) );
  SDFFX1 \fifo_reg[1][12]  ( .D(n1098), .SI(\fifo[1][11] ), .SE(test_se), 
        .CLK(n21), .Q(\fifo[1][12] ), .QN(n1840) );
  SDFFX1 \fifo_reg[1][11]  ( .D(n1097), .SI(\fifo[1][10] ), .SE(test_se), 
        .CLK(n21), .Q(\fifo[1][11] ), .QN(n1841) );
  SDFFX1 \fifo_reg[1][10]  ( .D(n1096), .SI(\fifo[1][9] ), .SE(test_se), .CLK(
        n21), .Q(\fifo[1][10] ), .QN(n1842) );
  SDFFX1 \fifo_reg[1][9]  ( .D(n1095), .SI(\fifo[1][8] ), .SE(test_se), .CLK(
        n20), .Q(\fifo[1][9] ), .QN(n1843) );
  SDFFX1 \fifo_reg[1][8]  ( .D(n1094), .SI(\fifo[1][7] ), .SE(test_se), .CLK(
        n20), .Q(\fifo[1][8] ), .QN(n1844) );
  SDFFX1 \fifo_reg[1][7]  ( .D(n1093), .SI(\fifo[1][6] ), .SE(test_se), .CLK(
        n20), .Q(\fifo[1][7] ), .QN(n1845) );
  SDFFX1 \fifo_reg[1][6]  ( .D(n1092), .SI(\fifo[1][5] ), .SE(test_se), .CLK(
        n20), .Q(\fifo[1][6] ), .QN(n1846) );
  SDFFX1 \fifo_reg[1][5]  ( .D(n1091), .SI(\fifo[1][4] ), .SE(test_se), .CLK(
        n20), .Q(\fifo[1][5] ), .QN(n1847) );
  SDFFX1 \fifo_reg[1][4]  ( .D(n1090), .SI(\fifo[1][3] ), .SE(test_se), .CLK(
        n20), .Q(\fifo[1][4] ), .QN(n1848) );
  SDFFX1 \fifo_reg[1][3]  ( .D(n1089), .SI(\fifo[1][2] ), .SE(test_se), .CLK(
        n20), .Q(\fifo[1][3] ), .QN(n1849) );
  SDFFX1 \fifo_reg[1][2]  ( .D(n1088), .SI(\fifo[1][1] ), .SE(test_se), .CLK(
        n20), .Q(\fifo[1][2] ), .QN(n1850) );
  SDFFX1 \fifo_reg[1][1]  ( .D(n1087), .SI(\fifo[1][0] ), .SE(test_se), .CLK(
        n20), .Q(\fifo[1][1] ), .QN(n1851) );
  SDFFX1 \fifo_reg[1][0]  ( .D(n1086), .SI(\fifo[0][31] ), .SE(test_se), .CLK(
        n20), .Q(\fifo[1][0] ), .QN(n1852) );
  SDFFX1 \fifo_reg[2][31]  ( .D(n1085), .SI(\fifo[2][30] ), .SE(test_se), 
        .CLK(n24), .Q(\fifo[2][31] ), .QN(n1853) );
  SDFFX1 \fifo_reg[2][30]  ( .D(n1084), .SI(\fifo[2][29] ), .SE(test_se), 
        .CLK(n24), .Q(\fifo[2][30] ), .QN(n1854) );
  SDFFX1 \fifo_reg[2][29]  ( .D(n1083), .SI(\fifo[2][28] ), .SE(test_se), 
        .CLK(n24), .Q(\fifo[2][29] ), .QN(n1855) );
  SDFFX1 \fifo_reg[2][28]  ( .D(n1082), .SI(\fifo[2][27] ), .SE(test_se), 
        .CLK(n24), .Q(\fifo[2][28] ), .QN(n1856) );
  SDFFX1 \fifo_reg[2][27]  ( .D(n1081), .SI(\fifo[2][26] ), .SE(test_se), 
        .CLK(n24), .Q(\fifo[2][27] ), .QN(n1857) );
  SDFFX1 \fifo_reg[2][26]  ( .D(n1080), .SI(\fifo[2][25] ), .SE(test_se), 
        .CLK(n24), .Q(\fifo[2][26] ), .QN(n1858) );
  SDFFX1 \fifo_reg[2][25]  ( .D(n1079), .SI(\fifo[2][24] ), .SE(test_se), 
        .CLK(n24), .Q(\fifo[2][25] ), .QN(n1859) );
  SDFFX1 \fifo_reg[2][24]  ( .D(n1078), .SI(\fifo[2][23] ), .SE(test_se), 
        .CLK(n24), .Q(\fifo[2][24] ), .QN(n1860) );
  SDFFX1 \fifo_reg[2][23]  ( .D(n1077), .SI(\fifo[2][22] ), .SE(test_se), 
        .CLK(n24), .Q(\fifo[2][23] ), .QN(n1861) );
  SDFFX1 \fifo_reg[2][22]  ( .D(n1076), .SI(\fifo[2][21] ), .SE(test_se), 
        .CLK(n24), .Q(\fifo[2][22] ), .QN(n1862) );
  SDFFX1 \fifo_reg[2][21]  ( .D(n1075), .SI(\fifo[2][20] ), .SE(test_se), 
        .CLK(n24), .Q(\fifo[2][21] ), .QN(n1863) );
  SDFFX1 \fifo_reg[2][20]  ( .D(n1074), .SI(\fifo[2][19] ), .SE(test_se), 
        .CLK(n24), .Q(\fifo[2][20] ), .QN(n1864) );
  SDFFX1 \fifo_reg[2][19]  ( .D(n1073), .SI(\fifo[2][18] ), .SE(test_se), 
        .CLK(n23), .Q(\fifo[2][19] ), .QN(n1865) );
  SDFFX1 \fifo_reg[2][18]  ( .D(n1072), .SI(\fifo[2][17] ), .SE(test_se), 
        .CLK(n23), .Q(\fifo[2][18] ), .QN(n1866) );
  SDFFX1 \fifo_reg[2][17]  ( .D(n1071), .SI(\fifo[2][16] ), .SE(test_se), 
        .CLK(n23), .Q(\fifo[2][17] ), .QN(n1867) );
  SDFFX1 \fifo_reg[2][16]  ( .D(n1070), .SI(\fifo[2][15] ), .SE(test_se), 
        .CLK(n23), .Q(\fifo[2][16] ), .QN(n1868) );
  SDFFX1 \fifo_reg[2][15]  ( .D(n1069), .SI(\fifo[2][14] ), .SE(test_se), 
        .CLK(n23), .Q(\fifo[2][15] ), .QN(n1869) );
  SDFFX1 \fifo_reg[2][14]  ( .D(n1068), .SI(\fifo[2][13] ), .SE(test_se), 
        .CLK(n23), .Q(\fifo[2][14] ), .QN(n1870) );
  SDFFX1 \fifo_reg[2][13]  ( .D(n1067), .SI(\fifo[2][12] ), .SE(test_se), 
        .CLK(n23), .Q(\fifo[2][13] ), .QN(n1871) );
  SDFFX1 \fifo_reg[2][12]  ( .D(n1066), .SI(\fifo[2][11] ), .SE(test_se), 
        .CLK(n23), .Q(\fifo[2][12] ), .QN(n1872) );
  SDFFX1 \fifo_reg[2][11]  ( .D(n1065), .SI(\fifo[2][10] ), .SE(test_se), 
        .CLK(n23), .Q(\fifo[2][11] ), .QN(n1873) );
  SDFFX1 \fifo_reg[2][10]  ( .D(n1064), .SI(\fifo[2][9] ), .SE(test_se), .CLK(
        n23), .Q(\fifo[2][10] ), .QN(n1874) );
  SDFFX1 \fifo_reg[2][9]  ( .D(n1063), .SI(\fifo[2][8] ), .SE(test_se), .CLK(
        n23), .Q(\fifo[2][9] ), .QN(n1875) );
  SDFFX1 \fifo_reg[2][8]  ( .D(n1062), .SI(\fifo[2][7] ), .SE(test_se), .CLK(
        n23), .Q(\fifo[2][8] ), .QN(n1876) );
  SDFFX1 \fifo_reg[2][7]  ( .D(n1061), .SI(\fifo[2][6] ), .SE(test_se), .CLK(
        n23), .Q(\fifo[2][7] ), .QN(n1877) );
  SDFFX1 \fifo_reg[2][6]  ( .D(n1060), .SI(\fifo[2][5] ), .SE(test_se), .CLK(
        n23), .Q(\fifo[2][6] ), .QN(n1878) );
  SDFFX1 \fifo_reg[2][5]  ( .D(n1059), .SI(\fifo[2][4] ), .SE(test_se), .CLK(
        n22), .Q(\fifo[2][5] ), .QN(n1879) );
  SDFFX1 \fifo_reg[2][4]  ( .D(n1058), .SI(\fifo[2][3] ), .SE(test_se), .CLK(
        n22), .Q(\fifo[2][4] ), .QN(n1880) );
  SDFFX1 \fifo_reg[2][3]  ( .D(n1057), .SI(\fifo[2][2] ), .SE(test_se), .CLK(
        n22), .Q(\fifo[2][3] ), .QN(n1881) );
  SDFFX1 \fifo_reg[2][2]  ( .D(n1056), .SI(\fifo[2][1] ), .SE(test_se), .CLK(
        n22), .Q(\fifo[2][2] ), .QN(n1882) );
  SDFFX1 \fifo_reg[2][1]  ( .D(n1055), .SI(\fifo[2][0] ), .SE(test_se), .CLK(
        n22), .Q(\fifo[2][1] ), .QN(n1883) );
  SDFFX1 \fifo_reg[2][0]  ( .D(n1054), .SI(\fifo[1][31] ), .SE(test_se), .CLK(
        n22), .Q(\fifo[2][0] ), .QN(n1884) );
  SDFFX1 \fifo_reg[3][31]  ( .D(n1053), .SI(\fifo[3][30] ), .SE(test_se), 
        .CLK(n7), .Q(\fifo[3][31] ), .QN(n1885) );
  SDFFX1 \fifo_reg[3][30]  ( .D(n1052), .SI(\fifo[3][29] ), .SE(test_se), 
        .CLK(n7), .Q(\fifo[3][30] ), .QN(n1886) );
  SDFFX1 \fifo_reg[3][29]  ( .D(n1051), .SI(\fifo[3][28] ), .SE(test_se), 
        .CLK(n7), .Q(\fifo[3][29] ), .QN(n1887) );
  SDFFX1 \fifo_reg[3][28]  ( .D(n1050), .SI(\fifo[3][27] ), .SE(test_se), 
        .CLK(n7), .Q(\fifo[3][28] ), .QN(n1888) );
  SDFFX1 \fifo_reg[3][27]  ( .D(n1049), .SI(\fifo[3][26] ), .SE(test_se), 
        .CLK(n8), .Q(\fifo[3][27] ), .QN(n1889) );
  SDFFX1 \fifo_reg[3][26]  ( .D(n1048), .SI(\fifo[3][25] ), .SE(test_se), 
        .CLK(n7), .Q(\fifo[3][26] ), .QN(n1890) );
  SDFFX1 \fifo_reg[3][25]  ( .D(n1047), .SI(\fifo[3][24] ), .SE(test_se), 
        .CLK(n7), .Q(\fifo[3][25] ), .QN(n1891) );
  SDFFX1 \fifo_reg[3][24]  ( .D(n1046), .SI(\fifo[3][23] ), .SE(test_se), 
        .CLK(n7), .Q(\fifo[3][24] ), .QN(n1892) );
  SDFFX1 \fifo_reg[3][23]  ( .D(n1045), .SI(\fifo[3][22] ), .SE(test_se), 
        .CLK(n7), .Q(\fifo[3][23] ), .QN(n1893) );
  SDFFX1 \fifo_reg[3][22]  ( .D(n1044), .SI(\fifo[3][21] ), .SE(test_se), 
        .CLK(n7), .Q(\fifo[3][22] ), .QN(n1894) );
  SDFFX1 \fifo_reg[3][21]  ( .D(n1043), .SI(\fifo[3][20] ), .SE(test_se), 
        .CLK(n7), .Q(\fifo[3][21] ), .QN(n1895) );
  SDFFX1 \fifo_reg[3][20]  ( .D(n1042), .SI(\fifo[3][19] ), .SE(test_se), 
        .CLK(n7), .Q(\fifo[3][20] ), .QN(n1896) );
  SDFFX1 \fifo_reg[3][19]  ( .D(n1041), .SI(\fifo[3][18] ), .SE(test_se), 
        .CLK(n6), .Q(\fifo[3][19] ), .QN(n1897) );
  SDFFX1 \fifo_reg[3][18]  ( .D(n1040), .SI(\fifo[3][17] ), .SE(test_se), 
        .CLK(n6), .Q(\fifo[3][18] ), .QN(n1898) );
  SDFFX1 \fifo_reg[3][17]  ( .D(n1039), .SI(\fifo[3][16] ), .SE(test_se), 
        .CLK(n6), .Q(\fifo[3][17] ), .QN(n1899) );
  SDFFX1 \fifo_reg[3][16]  ( .D(n1038), .SI(\fifo[3][15] ), .SE(test_se), 
        .CLK(n6), .Q(\fifo[3][16] ), .QN(n1900) );
  SDFFX1 \fifo_reg[3][15]  ( .D(n1037), .SI(\fifo[3][14] ), .SE(test_se), 
        .CLK(n6), .Q(\fifo[3][15] ), .QN(n1901) );
  SDFFX1 \fifo_reg[3][14]  ( .D(n1036), .SI(\fifo[3][13] ), .SE(test_se), 
        .CLK(n6), .Q(\fifo[3][14] ), .QN(n1902) );
  SDFFX1 \fifo_reg[3][13]  ( .D(n1035), .SI(\fifo[3][12] ), .SE(test_se), 
        .CLK(n6), .Q(\fifo[3][13] ), .QN(n1903) );
  SDFFX1 \fifo_reg[3][12]  ( .D(n1034), .SI(\fifo[3][11] ), .SE(test_se), 
        .CLK(n7), .Q(\fifo[3][12] ), .QN(n1904) );
  SDFFX1 \fifo_reg[3][11]  ( .D(n1033), .SI(\fifo[3][10] ), .SE(test_se), 
        .CLK(n6), .Q(\fifo[3][11] ), .QN(n1905) );
  SDFFX1 \fifo_reg[3][10]  ( .D(n1032), .SI(\fifo[3][9] ), .SE(test_se), .CLK(
        n6), .Q(\fifo[3][10] ), .QN(n1906) );
  SDFFX1 \fifo_reg[3][9]  ( .D(n1031), .SI(\fifo[3][8] ), .SE(test_se), .CLK(
        n6), .Q(\fifo[3][9] ), .QN(n1907) );
  SDFFX1 \fifo_reg[3][8]  ( .D(n1030), .SI(\fifo[3][7] ), .SE(test_se), .CLK(
        n6), .Q(\fifo[3][8] ), .QN(n1908) );
  SDFFX1 \fifo_reg[3][7]  ( .D(n1029), .SI(\fifo[3][6] ), .SE(test_se), .CLK(
        n6), .Q(\fifo[3][7] ), .QN(n1909) );
  SDFFX1 \fifo_reg[3][6]  ( .D(n1028), .SI(\fifo[3][5] ), .SE(test_se), .CLK(
        n25), .Q(\fifo[3][6] ), .QN(n1910) );
  SDFFX1 \fifo_reg[3][5]  ( .D(n1027), .SI(\fifo[3][4] ), .SE(test_se), .CLK(
        n25), .Q(\fifo[3][5] ), .QN(n1911) );
  SDFFX1 \fifo_reg[3][4]  ( .D(n1026), .SI(\fifo[3][3] ), .SE(test_se), .CLK(
        n25), .Q(\fifo[3][4] ), .QN(n1912) );
  SDFFX1 \fifo_reg[3][3]  ( .D(n1025), .SI(\fifo[3][2] ), .SE(test_se), .CLK(
        n25), .Q(\fifo[3][3] ), .QN(n1913) );
  SDFFX1 \fifo_reg[3][2]  ( .D(n1024), .SI(\fifo[3][1] ), .SE(test_se), .CLK(
        n25), .Q(\fifo[3][2] ), .QN(n1914) );
  SDFFX1 \fifo_reg[3][1]  ( .D(n1023), .SI(\fifo[3][0] ), .SE(test_se), .CLK(
        n24), .Q(\fifo[3][1] ), .QN(n1915) );
  SDFFX1 \fifo_reg[3][0]  ( .D(n1022), .SI(\fifo[2][31] ), .SE(test_se), .CLK(
        n24), .Q(\fifo[3][0] ), .QN(n1916) );
  SDFFX1 \fifo_reg[4][31]  ( .D(n1021), .SI(\fifo[4][30] ), .SE(test_se), 
        .CLK(n10), .Q(\fifo[4][31] ), .QN(n1917) );
  SDFFX1 \fifo_reg[4][30]  ( .D(n1020), .SI(\fifo[4][29] ), .SE(test_se), 
        .CLK(n10), .Q(\fifo[4][30] ), .QN(n1918) );
  SDFFX1 \fifo_reg[4][29]  ( .D(n1019), .SI(\fifo[4][28] ), .SE(test_se), 
        .CLK(n9), .Q(\fifo[4][29] ), .QN(n1919) );
  SDFFX1 \fifo_reg[4][28]  ( .D(n1018), .SI(\fifo[4][27] ), .SE(test_se), 
        .CLK(n9), .Q(\fifo[4][28] ), .QN(n1920) );
  SDFFX1 \fifo_reg[4][27]  ( .D(n1017), .SI(\fifo[4][26] ), .SE(test_se), 
        .CLK(n9), .Q(\fifo[4][27] ), .QN(n1921) );
  SDFFX1 \fifo_reg[4][26]  ( .D(n1016), .SI(\fifo[4][25] ), .SE(test_se), 
        .CLK(n9), .Q(\fifo[4][26] ), .QN(n1922) );
  SDFFX1 \fifo_reg[4][25]  ( .D(n1015), .SI(\fifo[4][24] ), .SE(test_se), 
        .CLK(n9), .Q(\fifo[4][25] ), .QN(n1923) );
  SDFFX1 \fifo_reg[4][24]  ( .D(n1014), .SI(\fifo[4][23] ), .SE(test_se), 
        .CLK(n9), .Q(\fifo[4][24] ), .QN(n1924) );
  SDFFX1 \fifo_reg[4][23]  ( .D(n1013), .SI(\fifo[4][22] ), .SE(test_se), 
        .CLK(n9), .Q(\fifo[4][23] ), .QN(n1925) );
  SDFFX1 \fifo_reg[4][22]  ( .D(n1012), .SI(\fifo[4][21] ), .SE(test_se), 
        .CLK(n9), .Q(\fifo[4][22] ), .QN(n1926) );
  SDFFX1 \fifo_reg[4][21]  ( .D(n1011), .SI(\fifo[4][20] ), .SE(test_se), 
        .CLK(n9), .Q(\fifo[4][21] ), .QN(n1927) );
  SDFFX1 \fifo_reg[4][20]  ( .D(n1010), .SI(\fifo[4][19] ), .SE(test_se), 
        .CLK(n9), .Q(\fifo[4][20] ), .QN(n1928) );
  SDFFX1 \fifo_reg[4][19]  ( .D(n1009), .SI(\fifo[4][18] ), .SE(test_se), 
        .CLK(n9), .Q(\fifo[4][19] ), .QN(n1929) );
  SDFFX1 \fifo_reg[4][18]  ( .D(n1008), .SI(\fifo[4][17] ), .SE(test_se), 
        .CLK(n9), .Q(\fifo[4][18] ), .QN(n1930) );
  SDFFX1 \fifo_reg[4][17]  ( .D(n1007), .SI(\fifo[4][16] ), .SE(test_se), 
        .CLK(n9), .Q(\fifo[4][17] ), .QN(n1931) );
  SDFFX1 \fifo_reg[4][16]  ( .D(n1006), .SI(\fifo[4][15] ), .SE(test_se), 
        .CLK(n9), .Q(\fifo[4][16] ), .QN(n1932) );
  SDFFX1 \fifo_reg[4][15]  ( .D(n1005), .SI(\fifo[4][14] ), .SE(test_se), 
        .CLK(n8), .Q(\fifo[4][15] ), .QN(n1933) );
  SDFFX1 \fifo_reg[4][14]  ( .D(n1004), .SI(\fifo[4][13] ), .SE(test_se), 
        .CLK(n8), .Q(\fifo[4][14] ), .QN(n1934) );
  SDFFX1 \fifo_reg[4][13]  ( .D(n1003), .SI(\fifo[4][12] ), .SE(test_se), 
        .CLK(n8), .Q(\fifo[4][13] ), .QN(n1935) );
  SDFFX1 \fifo_reg[4][12]  ( .D(n1002), .SI(\fifo[4][11] ), .SE(test_se), 
        .CLK(n8), .Q(\fifo[4][12] ), .QN(n1936) );
  SDFFX1 \fifo_reg[4][11]  ( .D(n1001), .SI(\fifo[4][10] ), .SE(test_se), 
        .CLK(n8), .Q(\fifo[4][11] ), .QN(n1937) );
  SDFFX1 \fifo_reg[4][10]  ( .D(n1000), .SI(\fifo[4][9] ), .SE(test_se), .CLK(
        n10), .Q(\fifo[4][10] ), .QN(n1938) );
  SDFFX1 \fifo_reg[4][9]  ( .D(n999), .SI(\fifo[4][8] ), .SE(test_se), .CLK(n8), .Q(\fifo[4][9] ), .QN(n1459) );
  SDFFX1 \fifo_reg[4][8]  ( .D(n998), .SI(\fifo[4][7] ), .SE(test_se), .CLK(n8), .Q(\fifo[4][8] ), .QN(n1460) );
  SDFFX1 \fifo_reg[4][7]  ( .D(n997), .SI(\fifo[4][6] ), .SE(test_se), .CLK(n8), .Q(\fifo[4][7] ), .QN(n1461) );
  SDFFX1 \fifo_reg[4][6]  ( .D(n996), .SI(\fifo[4][5] ), .SE(test_se), .CLK(n8), .Q(\fifo[4][6] ), .QN(n1462) );
  SDFFX1 \fifo_reg[4][5]  ( .D(n995), .SI(\fifo[4][4] ), .SE(test_se), .CLK(n8), .Q(\fifo[4][5] ), .QN(n1463) );
  SDFFX1 \fifo_reg[4][4]  ( .D(n994), .SI(\fifo[4][3] ), .SE(test_se), .CLK(n8), .Q(\fifo[4][4] ), .QN(n1464) );
  SDFFX1 \fifo_reg[4][3]  ( .D(n993), .SI(\fifo[4][2] ), .SE(test_se), .CLK(n8), .Q(\fifo[4][3] ), .QN(n1465) );
  SDFFX1 \fifo_reg[4][2]  ( .D(n992), .SI(\fifo[4][1] ), .SE(test_se), .CLK(n8), .Q(\fifo[4][2] ), .QN(n1466) );
  SDFFX1 \fifo_reg[4][1]  ( .D(n991), .SI(\fifo[4][0] ), .SE(test_se), .CLK(n7), .Q(\fifo[4][1] ), .QN(n1467) );
  SDFFX1 \fifo_reg[4][0]  ( .D(n990), .SI(\fifo[3][31] ), .SE(test_se), .CLK(
        n7), .Q(\fifo[4][0] ), .QN(n1468) );
  SDFFX1 \fifo_reg[5][31]  ( .D(n989), .SI(\fifo[5][30] ), .SE(test_se), .CLK(
        n12), .Q(\fifo[5][31] ), .QN(n1469) );
  SDFFX1 \fifo_reg[5][30]  ( .D(n988), .SI(\fifo[5][29] ), .SE(test_se), .CLK(
        n12), .Q(\fifo[5][30] ), .QN(n1470) );
  SDFFX1 \fifo_reg[5][29]  ( .D(n987), .SI(\fifo[5][28] ), .SE(test_se), .CLK(
        n12), .Q(\fifo[5][29] ), .QN(n1471) );
  SDFFX1 \fifo_reg[5][28]  ( .D(n986), .SI(\fifo[5][27] ), .SE(test_se), .CLK(
        n12), .Q(\fifo[5][28] ), .QN(n1472) );
  SDFFX1 \fifo_reg[5][27]  ( .D(n985), .SI(\fifo[5][26] ), .SE(test_se), .CLK(
        n12), .Q(\fifo[5][27] ), .QN(n1473) );
  SDFFX1 \fifo_reg[5][26]  ( .D(n984), .SI(\fifo[5][25] ), .SE(test_se), .CLK(
        n12), .Q(\fifo[5][26] ), .QN(n1474) );
  SDFFX1 \fifo_reg[5][25]  ( .D(n983), .SI(\fifo[5][24] ), .SE(test_se), .CLK(
        n12), .Q(\fifo[5][25] ), .QN(n1475) );
  SDFFX1 \fifo_reg[5][24]  ( .D(n982), .SI(\fifo[5][23] ), .SE(test_se), .CLK(
        n11), .Q(\fifo[5][24] ), .QN(n1476) );
  SDFFX1 \fifo_reg[5][23]  ( .D(n981), .SI(\fifo[5][22] ), .SE(test_se), .CLK(
        n11), .Q(\fifo[5][23] ), .QN(n1477) );
  SDFFX1 \fifo_reg[5][22]  ( .D(n980), .SI(\fifo[5][21] ), .SE(test_se), .CLK(
        n11), .Q(\fifo[5][22] ), .QN(n1478) );
  SDFFX1 \fifo_reg[5][21]  ( .D(n979), .SI(\fifo[5][20] ), .SE(test_se), .CLK(
        n11), .Q(\fifo[5][21] ), .QN(n1479) );
  SDFFX1 \fifo_reg[5][20]  ( .D(n978), .SI(\fifo[5][19] ), .SE(test_se), .CLK(
        n11), .Q(\fifo[5][20] ), .QN(n1480) );
  SDFFX1 \fifo_reg[5][19]  ( .D(n977), .SI(\fifo[5][18] ), .SE(test_se), .CLK(
        n11), .Q(\fifo[5][19] ), .QN(n1481) );
  SDFFX1 \fifo_reg[5][18]  ( .D(n976), .SI(\fifo[5][17] ), .SE(test_se), .CLK(
        n11), .Q(\fifo[5][18] ), .QN(n1482) );
  SDFFX1 \fifo_reg[5][17]  ( .D(n975), .SI(\fifo[5][16] ), .SE(test_se), .CLK(
        n11), .Q(\fifo[5][17] ), .QN(n1483) );
  SDFFX1 \fifo_reg[5][16]  ( .D(n974), .SI(\fifo[5][15] ), .SE(test_se), .CLK(
        n11), .Q(\fifo[5][16] ), .QN(n1484) );
  SDFFX1 \fifo_reg[5][15]  ( .D(n973), .SI(\fifo[5][14] ), .SE(test_se), .CLK(
        n11), .Q(\fifo[5][15] ), .QN(n1485) );
  SDFFX1 \fifo_reg[5][14]  ( .D(n972), .SI(\fifo[5][13] ), .SE(test_se), .CLK(
        n11), .Q(\fifo[5][14] ), .QN(n1486) );
  SDFFX1 \fifo_reg[5][13]  ( .D(n971), .SI(\fifo[5][12] ), .SE(test_se), .CLK(
        n11), .Q(\fifo[5][13] ), .QN(n1487) );
  SDFFX1 \fifo_reg[5][12]  ( .D(n970), .SI(\fifo[5][11] ), .SE(test_se), .CLK(
        n11), .Q(\fifo[5][12] ), .QN(n1488) );
  SDFFX1 \fifo_reg[5][11]  ( .D(n969), .SI(\fifo[5][10] ), .SE(test_se), .CLK(
        n11), .Q(\fifo[5][11] ), .QN(n1489) );
  SDFFX1 \fifo_reg[5][10]  ( .D(n968), .SI(\fifo[5][9] ), .SE(test_se), .CLK(
        n10), .Q(\fifo[5][10] ), .QN(n1490) );
  SDFFX1 \fifo_reg[5][9]  ( .D(n967), .SI(\fifo[5][8] ), .SE(test_se), .CLK(
        n10), .Q(\fifo[5][9] ), .QN(n1491) );
  SDFFX1 \fifo_reg[5][8]  ( .D(n966), .SI(\fifo[5][7] ), .SE(test_se), .CLK(
        n10), .Q(\fifo[5][8] ), .QN(n1492) );
  SDFFX1 \fifo_reg[5][7]  ( .D(n965), .SI(\fifo[5][6] ), .SE(test_se), .CLK(
        n10), .Q(\fifo[5][7] ), .QN(n1493) );
  SDFFX1 \fifo_reg[5][6]  ( .D(n964), .SI(\fifo[5][5] ), .SE(test_se), .CLK(
        n10), .Q(\fifo[5][6] ), .QN(n1494) );
  SDFFX1 \fifo_reg[5][5]  ( .D(n963), .SI(\fifo[5][4] ), .SE(test_se), .CLK(
        n10), .Q(\fifo[5][5] ), .QN(n1495) );
  SDFFX1 \fifo_reg[5][4]  ( .D(n962), .SI(\fifo[5][3] ), .SE(test_se), .CLK(
        n10), .Q(\fifo[5][4] ), .QN(n1496) );
  SDFFX1 \fifo_reg[5][3]  ( .D(n961), .SI(\fifo[5][2] ), .SE(test_se), .CLK(
        n10), .Q(\fifo[5][3] ), .QN(n1497) );
  SDFFX1 \fifo_reg[5][2]  ( .D(n960), .SI(\fifo[5][1] ), .SE(test_se), .CLK(
        n10), .Q(\fifo[5][2] ), .QN(n1498) );
  SDFFX1 \fifo_reg[5][1]  ( .D(n959), .SI(\fifo[5][0] ), .SE(test_se), .CLK(
        n10), .Q(\fifo[5][1] ), .QN(n1499) );
  SDFFX1 \fifo_reg[5][0]  ( .D(n958), .SI(\fifo[4][31] ), .SE(test_se), .CLK(
        n10), .Q(\fifo[5][0] ), .QN(n1500) );
  SDFFX1 \fifo_reg[6][31]  ( .D(n957), .SI(\fifo[6][30] ), .SE(test_se), .CLK(
        n14), .Q(\fifo[6][31] ), .QN(n1501) );
  SDFFX1 \fifo_reg[6][30]  ( .D(n956), .SI(\fifo[6][29] ), .SE(test_se), .CLK(
        n14), .Q(\fifo[6][30] ), .QN(n1502) );
  SDFFX1 \fifo_reg[6][29]  ( .D(n955), .SI(\fifo[6][28] ), .SE(test_se), .CLK(
        n14), .Q(\fifo[6][29] ), .QN(n1503) );
  SDFFX1 \fifo_reg[6][28]  ( .D(n954), .SI(\fifo[6][27] ), .SE(test_se), .CLK(
        n14), .Q(\fifo[6][28] ), .QN(n1504) );
  SDFFX1 \fifo_reg[6][27]  ( .D(n953), .SI(\fifo[6][26] ), .SE(test_se), .CLK(
        n14), .Q(\fifo[6][27] ), .QN(n1505) );
  SDFFX1 \fifo_reg[6][26]  ( .D(n952), .SI(\fifo[6][25] ), .SE(test_se), .CLK(
        n14), .Q(\fifo[6][26] ), .QN(n1506) );
  SDFFX1 \fifo_reg[6][25]  ( .D(n951), .SI(\fifo[6][24] ), .SE(test_se), .CLK(
        n14), .Q(\fifo[6][25] ), .QN(n1507) );
  SDFFX1 \fifo_reg[6][24]  ( .D(n950), .SI(\fifo[6][23] ), .SE(test_se), .CLK(
        n14), .Q(\fifo[6][24] ), .QN(n1508) );
  SDFFX1 \fifo_reg[6][23]  ( .D(n949), .SI(\fifo[6][22] ), .SE(test_se), .CLK(
        n14), .Q(\fifo[6][23] ), .QN(n1509) );
  SDFFX1 \fifo_reg[6][22]  ( .D(n948), .SI(\fifo[6][21] ), .SE(test_se), .CLK(
        n14), .Q(\fifo[6][22] ), .QN(n1510) );
  SDFFX1 \fifo_reg[6][21]  ( .D(n947), .SI(\fifo[6][20] ), .SE(test_se), .CLK(
        n14), .Q(\fifo[6][21] ), .QN(n1511) );
  SDFFX1 \fifo_reg[6][20]  ( .D(n946), .SI(\fifo[6][19] ), .SE(test_se), .CLK(
        n13), .Q(\fifo[6][20] ), .QN(n1512) );
  SDFFX1 \fifo_reg[6][19]  ( .D(n945), .SI(\fifo[6][18] ), .SE(test_se), .CLK(
        n13), .Q(\fifo[6][19] ), .QN(n1513) );
  SDFFX1 \fifo_reg[6][18]  ( .D(n944), .SI(\fifo[6][17] ), .SE(test_se), .CLK(
        n13), .Q(\fifo[6][18] ), .QN(n1514) );
  SDFFX1 \fifo_reg[6][17]  ( .D(n943), .SI(\fifo[6][16] ), .SE(test_se), .CLK(
        n13), .Q(\fifo[6][17] ), .QN(n1515) );
  SDFFX1 \fifo_reg[6][16]  ( .D(n942), .SI(\fifo[6][15] ), .SE(test_se), .CLK(
        n13), .Q(\fifo[6][16] ), .QN(n1516) );
  SDFFX1 \fifo_reg[6][15]  ( .D(n941), .SI(\fifo[6][14] ), .SE(test_se), .CLK(
        n13), .Q(\fifo[6][15] ), .QN(n1517) );
  SDFFX1 \fifo_reg[6][14]  ( .D(n940), .SI(\fifo[6][13] ), .SE(test_se), .CLK(
        n13), .Q(\fifo[6][14] ), .QN(n1518) );
  SDFFX1 \fifo_reg[6][13]  ( .D(n939), .SI(\fifo[6][12] ), .SE(test_se), .CLK(
        n13), .Q(\fifo[6][13] ), .QN(n1519) );
  SDFFX1 \fifo_reg[6][12]  ( .D(n938), .SI(\fifo[6][11] ), .SE(test_se), .CLK(
        n13), .Q(\fifo[6][12] ), .QN(n1520) );
  SDFFX1 \fifo_reg[6][11]  ( .D(n937), .SI(\fifo[6][10] ), .SE(test_se), .CLK(
        n13), .Q(\fifo[6][11] ), .QN(n1521) );
  SDFFX1 \fifo_reg[6][10]  ( .D(n936), .SI(\fifo[6][9] ), .SE(test_se), .CLK(
        n13), .Q(\fifo[6][10] ), .QN(n1522) );
  SDFFX1 \fifo_reg[6][9]  ( .D(n935), .SI(\fifo[6][8] ), .SE(test_se), .CLK(
        n13), .Q(\fifo[6][9] ), .QN(n1523) );
  SDFFX1 \fifo_reg[6][8]  ( .D(n934), .SI(\fifo[6][7] ), .SE(test_se), .CLK(
        n13), .Q(\fifo[6][8] ), .QN(n1524) );
  SDFFX1 \fifo_reg[6][7]  ( .D(n933), .SI(\fifo[6][6] ), .SE(test_se), .CLK(
        n13), .Q(\fifo[6][7] ), .QN(n1525) );
  SDFFX1 \fifo_reg[6][6]  ( .D(n932), .SI(\fifo[6][5] ), .SE(test_se), .CLK(
        n12), .Q(\fifo[6][6] ), .QN(n1526) );
  SDFFX1 \fifo_reg[6][5]  ( .D(n931), .SI(\fifo[6][4] ), .SE(test_se), .CLK(
        n12), .Q(\fifo[6][5] ), .QN(n1527) );
  SDFFX1 \fifo_reg[6][4]  ( .D(n930), .SI(\fifo[6][3] ), .SE(test_se), .CLK(
        n12), .Q(\fifo[6][4] ), .QN(n1528) );
  SDFFX1 \fifo_reg[6][3]  ( .D(n929), .SI(\fifo[6][2] ), .SE(test_se), .CLK(
        n12), .Q(\fifo[6][3] ), .QN(n1529) );
  SDFFX1 \fifo_reg[6][2]  ( .D(n928), .SI(\fifo[6][1] ), .SE(test_se), .CLK(
        n12), .Q(\fifo[6][2] ), .QN(n1530) );
  SDFFX1 \fifo_reg[6][1]  ( .D(n927), .SI(\fifo[6][0] ), .SE(test_se), .CLK(
        n12), .Q(\fifo[6][1] ), .QN(n1531) );
  SDFFX1 \fifo_reg[6][0]  ( .D(n926), .SI(\fifo[5][31] ), .SE(test_se), .CLK(
        n12), .Q(\fifo[6][0] ), .QN(n1532) );
  SDFFX1 \fifo_reg[7][31]  ( .D(n925), .SI(\fifo[7][30] ), .SE(test_se), .CLK(
        n36), .Q(\fifo[7][31] ), .QN(n1533) );
  SDFFX1 \fifo_reg[7][30]  ( .D(n924), .SI(\fifo[7][29] ), .SE(test_se), .CLK(
        n36), .Q(\fifo[7][30] ), .QN(n1534) );
  SDFFX1 \fifo_reg[7][29]  ( .D(n923), .SI(\fifo[7][28] ), .SE(test_se), .CLK(
        n36), .Q(\fifo[7][29] ), .QN(n1535) );
  SDFFX1 \fifo_reg[7][28]  ( .D(n922), .SI(\fifo[7][27] ), .SE(test_se), .CLK(
        n36), .Q(\fifo[7][28] ), .QN(n1536) );
  SDFFX1 \fifo_reg[7][27]  ( .D(n921), .SI(\fifo[7][26] ), .SE(test_se), .CLK(
        n36), .Q(\fifo[7][27] ), .QN(n1537) );
  SDFFX1 \fifo_reg[7][26]  ( .D(n920), .SI(\fifo[7][25] ), .SE(test_se), .CLK(
        n36), .Q(\fifo[7][26] ), .QN(n1538) );
  SDFFX1 \fifo_reg[7][25]  ( .D(n919), .SI(\fifo[7][24] ), .SE(test_se), .CLK(
        n35), .Q(\fifo[7][25] ), .QN(n1539) );
  SDFFX1 \fifo_reg[7][24]  ( .D(n918), .SI(\fifo[7][23] ), .SE(test_se), .CLK(
        n35), .Q(\fifo[7][24] ), .QN(n1540) );
  SDFFX1 \fifo_reg[7][23]  ( .D(n917), .SI(\fifo[7][22] ), .SE(test_se), .CLK(
        n35), .Q(\fifo[7][23] ), .QN(n1541) );
  SDFFX1 \fifo_reg[7][22]  ( .D(n916), .SI(\fifo[7][21] ), .SE(test_se), .CLK(
        n35), .Q(\fifo[7][22] ), .QN(n1542) );
  SDFFX1 \fifo_reg[7][21]  ( .D(n915), .SI(\fifo[7][20] ), .SE(test_se), .CLK(
        n35), .Q(\fifo[7][21] ), .QN(n1543) );
  SDFFX1 \fifo_reg[7][20]  ( .D(n914), .SI(\fifo[7][19] ), .SE(test_se), .CLK(
        n35), .Q(\fifo[7][20] ), .QN(n1544) );
  SDFFX1 \fifo_reg[7][19]  ( .D(n913), .SI(\fifo[7][18] ), .SE(test_se), .CLK(
        n35), .Q(\fifo[7][19] ), .QN(n1545) );
  SDFFX1 \fifo_reg[7][18]  ( .D(n912), .SI(\fifo[7][17] ), .SE(test_se), .CLK(
        n35), .Q(\fifo[7][18] ), .QN(n1546) );
  SDFFX1 \fifo_reg[7][17]  ( .D(n911), .SI(\fifo[7][16] ), .SE(test_se), .CLK(
        n35), .Q(\fifo[7][17] ), .QN(n1547) );
  SDFFX1 \fifo_reg[7][16]  ( .D(n910), .SI(\fifo[7][15] ), .SE(test_se), .CLK(
        n35), .Q(\fifo[7][16] ), .QN(n1548) );
  SDFFX1 \fifo_reg[7][15]  ( .D(n909), .SI(\fifo[7][14] ), .SE(test_se), .CLK(
        n35), .Q(\fifo[7][15] ), .QN(n1549) );
  SDFFX1 \fifo_reg[7][14]  ( .D(n908), .SI(\fifo[7][13] ), .SE(test_se), .CLK(
        n35), .Q(\fifo[7][14] ), .QN(n1550) );
  SDFFX1 \fifo_reg[7][13]  ( .D(n907), .SI(\fifo[7][12] ), .SE(test_se), .CLK(
        n40), .Q(\fifo[7][13] ), .QN(n1551) );
  SDFFX1 \fifo_reg[7][12]  ( .D(n906), .SI(\fifo[7][11] ), .SE(test_se), .CLK(
        n15), .Q(\fifo[7][12] ), .QN(n1552) );
  SDFFX1 \fifo_reg[7][11]  ( .D(n905), .SI(\fifo[7][10] ), .SE(test_se), .CLK(
        n15), .Q(\fifo[7][11] ), .QN(n1553) );
  SDFFX1 \fifo_reg[7][10]  ( .D(n904), .SI(\fifo[7][9] ), .SE(test_se), .CLK(
        n15), .Q(\fifo[7][10] ), .QN(n1554) );
  SDFFX1 \fifo_reg[7][9]  ( .D(n903), .SI(\fifo[7][8] ), .SE(test_se), .CLK(
        n15), .Q(\fifo[7][9] ), .QN(n1555) );
  SDFFX1 \fifo_reg[7][8]  ( .D(n902), .SI(\fifo[7][7] ), .SE(test_se), .CLK(
        n15), .Q(\fifo[7][8] ), .QN(n1556) );
  SDFFX1 \fifo_reg[7][7]  ( .D(n901), .SI(\fifo[7][6] ), .SE(test_se), .CLK(
        n15), .Q(\fifo[7][7] ), .QN(n1557) );
  SDFFX1 \fifo_reg[7][6]  ( .D(n900), .SI(\fifo[7][5] ), .SE(test_se), .CLK(
        n15), .Q(\fifo[7][6] ), .QN(n1558) );
  SDFFX1 \fifo_reg[7][5]  ( .D(n899), .SI(\fifo[7][4] ), .SE(test_se), .CLK(
        n15), .Q(\fifo[7][5] ), .QN(n1559) );
  SDFFX1 \fifo_reg[7][4]  ( .D(n898), .SI(\fifo[7][3] ), .SE(test_se), .CLK(
        n15), .Q(\fifo[7][4] ), .QN(n1560) );
  SDFFX1 \fifo_reg[7][3]  ( .D(n897), .SI(\fifo[7][2] ), .SE(test_se), .CLK(
        n15), .Q(\fifo[7][3] ), .QN(n1561) );
  SDFFX1 \fifo_reg[7][2]  ( .D(n896), .SI(\fifo[7][1] ), .SE(test_se), .CLK(
        n14), .Q(\fifo[7][2] ), .QN(n1562) );
  SDFFX1 \fifo_reg[7][1]  ( .D(n895), .SI(\fifo[7][0] ), .SE(test_se), .CLK(
        n14), .Q(\fifo[7][1] ), .QN(n1563) );
  SDFFX1 \fifo_reg[7][0]  ( .D(n894), .SI(\fifo[6][31] ), .SE(test_se), .CLK(
        n14), .Q(\fifo[7][0] ), .QN(n1564) );
  SDFFX1 \fifo_reg[8][31]  ( .D(n893), .SI(\fifo[8][30] ), .SE(test_se), .CLK(
        n38), .Q(\fifo[8][31] ), .QN(n1565) );
  SDFFX1 \fifo_reg[8][30]  ( .D(n892), .SI(\fifo[8][29] ), .SE(test_se), .CLK(
        n38), .Q(\fifo[8][30] ), .QN(n1566) );
  SDFFX1 \fifo_reg[8][29]  ( .D(n891), .SI(\fifo[8][28] ), .SE(test_se), .CLK(
        n38), .Q(\fifo[8][29] ), .QN(n1567) );
  SDFFX1 \fifo_reg[8][28]  ( .D(n890), .SI(\fifo[8][27] ), .SE(test_se), .CLK(
        n38), .Q(\fifo[8][28] ), .QN(n1568) );
  SDFFX1 \fifo_reg[8][27]  ( .D(n889), .SI(\fifo[8][26] ), .SE(test_se), .CLK(
        n38), .Q(\fifo[8][27] ), .QN(n1569) );
  SDFFX1 \fifo_reg[8][26]  ( .D(n888), .SI(\fifo[8][25] ), .SE(test_se), .CLK(
        n38), .Q(\fifo[8][26] ), .QN(n1570) );
  SDFFX1 \fifo_reg[8][25]  ( .D(n887), .SI(\fifo[8][24] ), .SE(test_se), .CLK(
        n38), .Q(\fifo[8][25] ), .QN(n1571) );
  SDFFX1 \fifo_reg[8][24]  ( .D(n886), .SI(\fifo[8][23] ), .SE(test_se), .CLK(
        n38), .Q(\fifo[8][24] ), .QN(n1572) );
  SDFFX1 \fifo_reg[8][23]  ( .D(n885), .SI(\fifo[8][22] ), .SE(test_se), .CLK(
        n38), .Q(\fifo[8][23] ), .QN(n1573) );
  SDFFX1 \fifo_reg[8][22]  ( .D(n884), .SI(\fifo[8][21] ), .SE(test_se), .CLK(
        n38), .Q(\fifo[8][22] ), .QN(n1574) );
  SDFFX1 \fifo_reg[8][21]  ( .D(n883), .SI(\fifo[8][20] ), .SE(test_se), .CLK(
        n37), .Q(\fifo[8][21] ), .QN(n1575) );
  SDFFX1 \fifo_reg[8][20]  ( .D(n882), .SI(\fifo[8][19] ), .SE(test_se), .CLK(
        n37), .Q(\fifo[8][20] ), .QN(n1576) );
  SDFFX1 \fifo_reg[8][19]  ( .D(n881), .SI(\fifo[8][18] ), .SE(test_se), .CLK(
        n37), .Q(\fifo[8][19] ), .QN(n1577) );
  SDFFX1 \fifo_reg[8][18]  ( .D(n880), .SI(\fifo[8][17] ), .SE(test_se), .CLK(
        n37), .Q(\fifo[8][18] ), .QN(n1578) );
  SDFFX1 \fifo_reg[8][17]  ( .D(n879), .SI(\fifo[8][16] ), .SE(test_se), .CLK(
        n37), .Q(\fifo[8][17] ), .QN(n1579) );
  SDFFX1 \fifo_reg[8][16]  ( .D(n878), .SI(\fifo[8][15] ), .SE(test_se), .CLK(
        n37), .Q(\fifo[8][16] ), .QN(n1580) );
  SDFFX1 \fifo_reg[8][15]  ( .D(n877), .SI(\fifo[8][14] ), .SE(test_se), .CLK(
        n37), .Q(\fifo[8][15] ), .QN(n1581) );
  SDFFX1 \fifo_reg[8][14]  ( .D(n876), .SI(\fifo[8][13] ), .SE(test_se), .CLK(
        n37), .Q(\fifo[8][14] ), .QN(n1582) );
  SDFFX1 \fifo_reg[8][13]  ( .D(n875), .SI(\fifo[8][12] ), .SE(test_se), .CLK(
        n37), .Q(\fifo[8][13] ), .QN(n1583) );
  SDFFX1 \fifo_reg[8][12]  ( .D(n874), .SI(\fifo[8][11] ), .SE(test_se), .CLK(
        n37), .Q(\fifo[8][12] ), .QN(n1584) );
  SDFFX1 \fifo_reg[8][11]  ( .D(n873), .SI(\fifo[8][10] ), .SE(test_se), .CLK(
        n37), .Q(\fifo[8][11] ), .QN(n1585) );
  SDFFX1 \fifo_reg[8][10]  ( .D(n872), .SI(\fifo[8][9] ), .SE(test_se), .CLK(
        n37), .Q(\fifo[8][10] ), .QN(n1586) );
  SDFFX1 \fifo_reg[8][9]  ( .D(n871), .SI(\fifo[8][8] ), .SE(test_se), .CLK(
        n37), .Q(\fifo[8][9] ), .QN(n1587) );
  SDFFX1 \fifo_reg[8][8]  ( .D(n870), .SI(\fifo[8][7] ), .SE(test_se), .CLK(
        n37), .Q(\fifo[8][8] ), .QN(n1588) );
  SDFFX1 \fifo_reg[8][7]  ( .D(n869), .SI(\fifo[8][6] ), .SE(test_se), .CLK(
        n36), .Q(\fifo[8][7] ), .QN(n1589) );
  SDFFX1 \fifo_reg[8][6]  ( .D(n868), .SI(\fifo[8][5] ), .SE(test_se), .CLK(
        n36), .Q(\fifo[8][6] ), .QN(n1590) );
  SDFFX1 \fifo_reg[8][5]  ( .D(n867), .SI(\fifo[8][4] ), .SE(test_se), .CLK(
        n36), .Q(\fifo[8][5] ), .QN(n1591) );
  SDFFX1 \fifo_reg[8][4]  ( .D(n866), .SI(\fifo[8][3] ), .SE(test_se), .CLK(
        n36), .Q(\fifo[8][4] ), .QN(n1592) );
  SDFFX1 \fifo_reg[8][3]  ( .D(n865), .SI(\fifo[8][2] ), .SE(test_se), .CLK(
        n36), .Q(\fifo[8][3] ), .QN(n1593) );
  SDFFX1 \fifo_reg[8][2]  ( .D(n864), .SI(\fifo[8][1] ), .SE(test_se), .CLK(
        n36), .Q(\fifo[8][2] ), .QN(n1594) );
  SDFFX1 \fifo_reg[8][1]  ( .D(n863), .SI(\fifo[8][0] ), .SE(test_se), .CLK(
        n36), .Q(\fifo[8][1] ), .QN(n1595) );
  SDFFX1 \fifo_reg[8][0]  ( .D(n862), .SI(\fifo[7][31] ), .SE(test_se), .CLK(
        n36), .Q(\fifo[8][0] ), .QN(n1596) );
  SDFFX1 \fifo_reg[9][31]  ( .D(n861), .SI(\fifo[9][30] ), .SE(test_se), .CLK(
        n41), .Q(\fifo[9][31] ), .QN(n1597) );
  SDFFX1 \fifo_reg[9][30]  ( .D(n860), .SI(\fifo[9][29] ), .SE(test_se), .CLK(
        n40), .Q(\fifo[9][30] ), .QN(n1598) );
  SDFFX1 \fifo_reg[9][29]  ( .D(n859), .SI(\fifo[9][28] ), .SE(test_se), .CLK(
        n40), .Q(\fifo[9][29] ), .QN(n1599) );
  SDFFX1 \fifo_reg[9][28]  ( .D(n858), .SI(\fifo[9][27] ), .SE(test_se), .CLK(
        n40), .Q(\fifo[9][28] ), .QN(n1600) );
  SDFFX1 \fifo_reg[9][27]  ( .D(n857), .SI(\fifo[9][26] ), .SE(test_se), .CLK(
        n40), .Q(\fifo[9][27] ), .QN(n1601) );
  SDFFX1 \fifo_reg[9][26]  ( .D(n856), .SI(\fifo[9][25] ), .SE(test_se), .CLK(
        n40), .Q(\fifo[9][26] ), .QN(n1602) );
  SDFFX1 \fifo_reg[9][25]  ( .D(n855), .SI(\fifo[9][24] ), .SE(test_se), .CLK(
        n40), .Q(\fifo[9][25] ), .QN(n1603) );
  SDFFX1 \fifo_reg[9][24]  ( .D(n854), .SI(\fifo[9][23] ), .SE(test_se), .CLK(
        n40), .Q(\fifo[9][24] ), .QN(n1604) );
  SDFFX1 \fifo_reg[9][23]  ( .D(n853), .SI(\fifo[9][22] ), .SE(test_se), .CLK(
        n40), .Q(\fifo[9][23] ), .QN(n1605) );
  SDFFX1 \fifo_reg[9][22]  ( .D(n852), .SI(\fifo[9][21] ), .SE(test_se), .CLK(
        n40), .Q(\fifo[9][22] ), .QN(n1606) );
  SDFFX1 \fifo_reg[9][21]  ( .D(n851), .SI(\fifo[9][20] ), .SE(test_se), .CLK(
        n40), .Q(\fifo[9][21] ), .QN(n1607) );
  SDFFX1 \fifo_reg[9][20]  ( .D(n850), .SI(\fifo[9][19] ), .SE(test_se), .CLK(
        n40), .Q(\fifo[9][20] ), .QN(n1608) );
  SDFFX1 \fifo_reg[9][19]  ( .D(n849), .SI(\fifo[9][18] ), .SE(test_se), .CLK(
        n40), .Q(\fifo[9][19] ), .QN(n1609) );
  SDFFX1 \fifo_reg[9][18]  ( .D(n848), .SI(\fifo[9][17] ), .SE(test_se), .CLK(
        n40), .Q(\fifo[9][18] ), .QN(n1610) );
  SDFFX1 \fifo_reg[9][17]  ( .D(n847), .SI(\fifo[9][16] ), .SE(test_se), .CLK(
        n39), .Q(\fifo[9][17] ), .QN(n1611) );
  SDFFX1 \fifo_reg[9][16]  ( .D(n846), .SI(\fifo[9][15] ), .SE(test_se), .CLK(
        n39), .Q(\fifo[9][16] ), .QN(n1612) );
  SDFFX1 \fifo_reg[9][15]  ( .D(n845), .SI(\fifo[9][14] ), .SE(test_se), .CLK(
        n39), .Q(\fifo[9][15] ), .QN(n1613) );
  SDFFX1 \fifo_reg[9][14]  ( .D(n844), .SI(\fifo[9][13] ), .SE(test_se), .CLK(
        n39), .Q(\fifo[9][14] ), .QN(n1614) );
  SDFFX1 \fifo_reg[9][13]  ( .D(n843), .SI(\fifo[9][12] ), .SE(test_se), .CLK(
        n39), .Q(\fifo[9][13] ), .QN(n1615) );
  SDFFX1 \fifo_reg[9][12]  ( .D(n842), .SI(\fifo[9][11] ), .SE(test_se), .CLK(
        n39), .Q(\fifo[9][12] ), .QN(n1616) );
  SDFFX1 \fifo_reg[9][11]  ( .D(n841), .SI(\fifo[9][10] ), .SE(test_se), .CLK(
        n39), .Q(\fifo[9][11] ), .QN(n1617) );
  SDFFX1 \fifo_reg[9][10]  ( .D(n840), .SI(\fifo[9][9] ), .SE(test_se), .CLK(
        n39), .Q(\fifo[9][10] ), .QN(n1618) );
  SDFFX1 \fifo_reg[9][9]  ( .D(n839), .SI(\fifo[9][8] ), .SE(test_se), .CLK(
        n39), .Q(\fifo[9][9] ), .QN(n1619) );
  SDFFX1 \fifo_reg[9][8]  ( .D(n838), .SI(\fifo[9][7] ), .SE(test_se), .CLK(
        n39), .Q(\fifo[9][8] ), .QN(n1620) );
  SDFFX1 \fifo_reg[9][7]  ( .D(n837), .SI(\fifo[9][6] ), .SE(test_se), .CLK(
        n39), .Q(\fifo[9][7] ), .QN(n1621) );
  SDFFX1 \fifo_reg[9][6]  ( .D(n836), .SI(\fifo[9][5] ), .SE(test_se), .CLK(
        n39), .Q(\fifo[9][6] ), .QN(n1622) );
  SDFFX1 \fifo_reg[9][5]  ( .D(n835), .SI(\fifo[9][4] ), .SE(test_se), .CLK(
        n39), .Q(\fifo[9][5] ), .QN(n1623) );
  SDFFX1 \fifo_reg[9][4]  ( .D(n834), .SI(\fifo[9][3] ), .SE(test_se), .CLK(
        n39), .Q(\fifo[9][4] ), .QN(n1624) );
  SDFFX1 \fifo_reg[9][3]  ( .D(n833), .SI(\fifo[9][2] ), .SE(test_se), .CLK(
        n38), .Q(\fifo[9][3] ), .QN(n1625) );
  SDFFX1 \fifo_reg[9][2]  ( .D(n832), .SI(\fifo[9][1] ), .SE(test_se), .CLK(
        n38), .Q(\fifo[9][2] ), .QN(n1626) );
  SDFFX1 \fifo_reg[9][1]  ( .D(n831), .SI(\fifo[9][0] ), .SE(test_se), .CLK(
        n38), .Q(\fifo[9][1] ), .QN(n1627) );
  SDFFX1 \fifo_reg[9][0]  ( .D(n830), .SI(\fifo[8][31] ), .SE(test_se), .CLK(
        n38), .Q(\fifo[9][0] ), .QN(n1628) );
  SDFFX1 \fifo_reg[10][31]  ( .D(n829), .SI(\fifo[10][30] ), .SE(test_se), 
        .CLK(n43), .Q(\fifo[10][31] ), .QN(n1629) );
  SDFFX1 \fifo_reg[10][30]  ( .D(n828), .SI(\fifo[10][29] ), .SE(test_se), 
        .CLK(n43), .Q(\fifo[10][30] ), .QN(n1630) );
  SDFFX1 \fifo_reg[10][29]  ( .D(n827), .SI(\fifo[10][28] ), .SE(test_se), 
        .CLK(n43), .Q(\fifo[10][29] ), .QN(n1631) );
  SDFFX1 \fifo_reg[10][28]  ( .D(n826), .SI(\fifo[10][27] ), .SE(test_se), 
        .CLK(n43), .Q(\fifo[10][28] ), .QN(n1632) );
  SDFFX1 \fifo_reg[10][27]  ( .D(n825), .SI(\fifo[10][26] ), .SE(test_se), 
        .CLK(n43), .Q(\fifo[10][27] ), .QN(n1633) );
  SDFFX1 \fifo_reg[10][26]  ( .D(n824), .SI(\fifo[10][25] ), .SE(test_se), 
        .CLK(n42), .Q(\fifo[10][26] ), .QN(n1634) );
  SDFFX1 \fifo_reg[10][25]  ( .D(n823), .SI(\fifo[10][24] ), .SE(test_se), 
        .CLK(n42), .Q(\fifo[10][25] ), .QN(n1635) );
  SDFFX1 \fifo_reg[10][24]  ( .D(n822), .SI(\fifo[10][23] ), .SE(test_se), 
        .CLK(n42), .Q(\fifo[10][24] ), .QN(n1636) );
  SDFFX1 \fifo_reg[10][23]  ( .D(n821), .SI(\fifo[10][22] ), .SE(test_se), 
        .CLK(n42), .Q(\fifo[10][23] ), .QN(n1637) );
  SDFFX1 \fifo_reg[10][22]  ( .D(n820), .SI(\fifo[10][21] ), .SE(test_se), 
        .CLK(n42), .Q(\fifo[10][22] ), .QN(n1638) );
  SDFFX1 \fifo_reg[10][21]  ( .D(n819), .SI(\fifo[10][20] ), .SE(test_se), 
        .CLK(n42), .Q(\fifo[10][21] ), .QN(n1639) );
  SDFFX1 \fifo_reg[10][20]  ( .D(n818), .SI(\fifo[10][19] ), .SE(test_se), 
        .CLK(n42), .Q(\fifo[10][20] ), .QN(n1640) );
  SDFFX1 \fifo_reg[10][19]  ( .D(n817), .SI(\fifo[10][18] ), .SE(test_se), 
        .CLK(n42), .Q(\fifo[10][19] ), .QN(n1641) );
  SDFFX1 \fifo_reg[10][18]  ( .D(n816), .SI(\fifo[10][17] ), .SE(test_se), 
        .CLK(n42), .Q(\fifo[10][18] ), .QN(n1642) );
  SDFFX1 \fifo_reg[10][17]  ( .D(n815), .SI(\fifo[10][16] ), .SE(test_se), 
        .CLK(n42), .Q(\fifo[10][17] ), .QN(n1643) );
  SDFFX1 \fifo_reg[10][16]  ( .D(n814), .SI(\fifo[10][15] ), .SE(test_se), 
        .CLK(n42), .Q(\fifo[10][16] ), .QN(n1644) );
  SDFFX1 \fifo_reg[10][15]  ( .D(n813), .SI(\fifo[10][14] ), .SE(test_se), 
        .CLK(n42), .Q(\fifo[10][15] ), .QN(n1645) );
  SDFFX1 \fifo_reg[10][14]  ( .D(n812), .SI(\fifo[10][13] ), .SE(test_se), 
        .CLK(n42), .Q(\fifo[10][14] ), .QN(n1646) );
  SDFFX1 \fifo_reg[10][13]  ( .D(n811), .SI(\fifo[10][12] ), .SE(test_se), 
        .CLK(n42), .Q(\fifo[10][13] ), .QN(n1647) );
  SDFFX1 \fifo_reg[10][12]  ( .D(n810), .SI(\fifo[10][11] ), .SE(test_se), 
        .CLK(n41), .Q(\fifo[10][12] ), .QN(n1648) );
  SDFFX1 \fifo_reg[10][11]  ( .D(n809), .SI(\fifo[10][10] ), .SE(test_se), 
        .CLK(n41), .Q(\fifo[10][11] ), .QN(n1649) );
  SDFFX1 \fifo_reg[10][10]  ( .D(n808), .SI(\fifo[10][9] ), .SE(test_se), 
        .CLK(n41), .Q(\fifo[10][10] ), .QN(n1650) );
  SDFFX1 \fifo_reg[10][9]  ( .D(n807), .SI(\fifo[10][8] ), .SE(test_se), .CLK(
        n41), .Q(\fifo[10][9] ), .QN(n1651) );
  SDFFX1 \fifo_reg[10][8]  ( .D(n806), .SI(\fifo[10][7] ), .SE(test_se), .CLK(
        n41), .Q(\fifo[10][8] ), .QN(n1652) );
  SDFFX1 \fifo_reg[10][7]  ( .D(n805), .SI(\fifo[10][6] ), .SE(test_se), .CLK(
        n41), .Q(\fifo[10][7] ), .QN(n1653) );
  SDFFX1 \fifo_reg[10][6]  ( .D(n804), .SI(\fifo[10][5] ), .SE(test_se), .CLK(
        n41), .Q(\fifo[10][6] ), .QN(n1654) );
  SDFFX1 \fifo_reg[10][5]  ( .D(n803), .SI(\fifo[10][4] ), .SE(test_se), .CLK(
        n41), .Q(\fifo[10][5] ), .QN(n1655) );
  SDFFX1 \fifo_reg[10][4]  ( .D(n802), .SI(\fifo[10][3] ), .SE(test_se), .CLK(
        n41), .Q(\fifo[10][4] ), .QN(n1656) );
  SDFFX1 \fifo_reg[10][3]  ( .D(n801), .SI(\fifo[10][2] ), .SE(test_se), .CLK(
        n41), .Q(\fifo[10][3] ), .QN(n1657) );
  SDFFX1 \fifo_reg[10][2]  ( .D(n800), .SI(\fifo[10][1] ), .SE(test_se), .CLK(
        n41), .Q(\fifo[10][2] ), .QN(n1658) );
  SDFFX1 \fifo_reg[10][1]  ( .D(n799), .SI(\fifo[10][0] ), .SE(test_se), .CLK(
        n41), .Q(\fifo[10][1] ), .QN(n1659) );
  SDFFX1 \fifo_reg[10][0]  ( .D(n798), .SI(\fifo[9][31] ), .SE(test_se), .CLK(
        n41), .Q(\fifo[10][0] ), .QN(n1660) );
  SDFFX1 \fifo_reg[11][31]  ( .D(n797), .SI(\fifo[11][30] ), .SE(test_se), 
        .CLK(n25), .Q(\fifo[11][31] ), .QN(n1661) );
  SDFFX1 \fifo_reg[11][30]  ( .D(n796), .SI(\fifo[11][29] ), .SE(test_se), 
        .CLK(n25), .Q(\fifo[11][30] ), .QN(n1662) );
  SDFFX1 \fifo_reg[11][29]  ( .D(n795), .SI(\fifo[11][28] ), .SE(test_se), 
        .CLK(n25), .Q(\fifo[11][29] ), .QN(n1663) );
  SDFFX1 \fifo_reg[11][28]  ( .D(n794), .SI(\fifo[11][27] ), .SE(test_se), 
        .CLK(n25), .Q(\fifo[11][28] ), .QN(n1664) );
  SDFFX1 \fifo_reg[11][27]  ( .D(n793), .SI(\fifo[11][26] ), .SE(test_se), 
        .CLK(n25), .Q(\fifo[11][27] ), .QN(n1665) );
  SDFFX1 \fifo_reg[11][26]  ( .D(n792), .SI(\fifo[11][25] ), .SE(test_se), 
        .CLK(n25), .Q(\fifo[11][26] ), .QN(n1666) );
  SDFFX1 \fifo_reg[11][25]  ( .D(n791), .SI(\fifo[11][24] ), .SE(test_se), 
        .CLK(n25), .Q(\fifo[11][25] ), .QN(n1667) );
  SDFFX1 \fifo_reg[11][24]  ( .D(n790), .SI(\fifo[11][23] ), .SE(test_se), 
        .CLK(n25), .Q(\fifo[11][24] ), .QN(n1668) );
  SDFFX1 \fifo_reg[11][23]  ( .D(n789), .SI(\fifo[11][22] ), .SE(test_se), 
        .CLK(n25), .Q(\fifo[11][23] ), .QN(n1669) );
  SDFFX1 \fifo_reg[11][22]  ( .D(n788), .SI(\fifo[11][21] ), .SE(test_se), 
        .CLK(n30), .Q(\fifo[11][22] ), .QN(n1670) );
  SDFFX1 \fifo_reg[11][21]  ( .D(n787), .SI(\fifo[11][20] ), .SE(test_se), 
        .CLK(n44), .Q(\fifo[11][21] ), .QN(n1671) );
  SDFFX1 \fifo_reg[11][20]  ( .D(n786), .SI(\fifo[11][19] ), .SE(test_se), 
        .CLK(n44), .Q(\fifo[11][20] ), .QN(n1672) );
  SDFFX1 \fifo_reg[11][19]  ( .D(n785), .SI(\fifo[11][18] ), .SE(test_se), 
        .CLK(n44), .Q(\fifo[11][19] ), .QN(n1673) );
  SDFFX1 \fifo_reg[11][18]  ( .D(n784), .SI(\fifo[11][17] ), .SE(test_se), 
        .CLK(n44), .Q(\fifo[11][18] ), .QN(n1674) );
  SDFFX1 \fifo_reg[11][17]  ( .D(n783), .SI(\fifo[11][16] ), .SE(test_se), 
        .CLK(n44), .Q(\fifo[11][17] ), .QN(n1675) );
  SDFFX1 \fifo_reg[11][16]  ( .D(n782), .SI(\fifo[11][15] ), .SE(test_se), 
        .CLK(n44), .Q(\fifo[11][16] ), .QN(n1676) );
  SDFFX1 \fifo_reg[11][15]  ( .D(n781), .SI(\fifo[11][14] ), .SE(test_se), 
        .CLK(n44), .Q(\fifo[11][15] ), .QN(n1677) );
  SDFFX1 \fifo_reg[11][14]  ( .D(n780), .SI(\fifo[11][13] ), .SE(test_se), 
        .CLK(n44), .Q(\fifo[11][14] ), .QN(n1678) );
  SDFFX1 \fifo_reg[11][13]  ( .D(n779), .SI(\fifo[11][12] ), .SE(test_se), 
        .CLK(n44), .Q(\fifo[11][13] ), .QN(n1679) );
  SDFFX1 \fifo_reg[11][12]  ( .D(n778), .SI(\fifo[11][11] ), .SE(test_se), 
        .CLK(n44), .Q(\fifo[11][12] ), .QN(n1680) );
  SDFFX1 \fifo_reg[11][11]  ( .D(n777), .SI(\fifo[11][10] ), .SE(test_se), 
        .CLK(n44), .Q(\fifo[11][11] ), .QN(n1681) );
  SDFFX1 \fifo_reg[11][10]  ( .D(n776), .SI(\fifo[11][9] ), .SE(test_se), 
        .CLK(n44), .Q(\fifo[11][10] ), .QN(n1682) );
  SDFFX1 \fifo_reg[11][9]  ( .D(n775), .SI(\fifo[11][8] ), .SE(test_se), .CLK(
        n44), .Q(\fifo[11][9] ), .QN(n1683) );
  SDFFX1 \fifo_reg[11][8]  ( .D(n774), .SI(\fifo[11][7] ), .SE(test_se), .CLK(
        n43), .Q(\fifo[11][8] ), .QN(n1684) );
  SDFFX1 \fifo_reg[11][7]  ( .D(n773), .SI(\fifo[11][6] ), .SE(test_se), .CLK(
        n43), .Q(\fifo[11][7] ), .QN(n1685) );
  SDFFX1 \fifo_reg[11][6]  ( .D(n772), .SI(\fifo[11][5] ), .SE(test_se), .CLK(
        n43), .Q(\fifo[11][6] ), .QN(n1686) );
  SDFFX1 \fifo_reg[11][5]  ( .D(n771), .SI(\fifo[11][4] ), .SE(test_se), .CLK(
        n43), .Q(\fifo[11][5] ), .QN(n1687) );
  SDFFX1 \fifo_reg[11][4]  ( .D(n770), .SI(\fifo[11][3] ), .SE(test_se), .CLK(
        n43), .Q(\fifo[11][4] ), .QN(n1688) );
  SDFFX1 \fifo_reg[11][3]  ( .D(n769), .SI(\fifo[11][2] ), .SE(test_se), .CLK(
        n43), .Q(\fifo[11][3] ), .QN(n1689) );
  SDFFX1 \fifo_reg[11][2]  ( .D(n768), .SI(\fifo[11][1] ), .SE(test_se), .CLK(
        n43), .Q(\fifo[11][2] ), .QN(n1690) );
  SDFFX1 \fifo_reg[11][1]  ( .D(n767), .SI(\fifo[11][0] ), .SE(test_se), .CLK(
        n43), .Q(\fifo[11][1] ), .QN(n1691) );
  SDFFX1 \fifo_reg[11][0]  ( .D(n766), .SI(\fifo[10][31] ), .SE(test_se), 
        .CLK(n43), .Q(\fifo[11][0] ), .QN(n1692) );
  SDFFX1 \fifo_reg[12][31]  ( .D(n765), .SI(\fifo[12][30] ), .SE(test_se), 
        .CLK(n28), .Q(\fifo[12][31] ), .QN(n1693) );
  SDFFX1 \fifo_reg[12][30]  ( .D(n764), .SI(\fifo[12][29] ), .SE(test_se), 
        .CLK(n28), .Q(\fifo[12][30] ), .QN(n1694) );
  SDFFX1 \fifo_reg[12][29]  ( .D(n763), .SI(\fifo[12][28] ), .SE(test_se), 
        .CLK(n28), .Q(\fifo[12][29] ), .QN(n1695) );
  SDFFX1 \fifo_reg[12][28]  ( .D(n762), .SI(\fifo[12][27] ), .SE(test_se), 
        .CLK(n28), .Q(\fifo[12][28] ), .QN(n1696) );
  SDFFX1 \fifo_reg[12][27]  ( .D(n761), .SI(\fifo[12][26] ), .SE(test_se), 
        .CLK(n27), .Q(\fifo[12][27] ), .QN(n1697) );
  SDFFX1 \fifo_reg[12][26]  ( .D(n760), .SI(\fifo[12][25] ), .SE(test_se), 
        .CLK(n27), .Q(\fifo[12][26] ), .QN(n1698) );
  SDFFX1 \fifo_reg[12][25]  ( .D(n759), .SI(\fifo[12][24] ), .SE(test_se), 
        .CLK(n27), .Q(\fifo[12][25] ), .QN(n1699) );
  SDFFX1 \fifo_reg[12][24]  ( .D(n758), .SI(\fifo[12][23] ), .SE(test_se), 
        .CLK(n27), .Q(\fifo[12][24] ), .QN(n1700) );
  SDFFX1 \fifo_reg[12][23]  ( .D(n757), .SI(\fifo[12][22] ), .SE(test_se), 
        .CLK(n27), .Q(\fifo[12][23] ), .QN(n1701) );
  SDFFX1 \fifo_reg[12][22]  ( .D(n756), .SI(\fifo[12][21] ), .SE(test_se), 
        .CLK(n27), .Q(\fifo[12][22] ), .QN(n1702) );
  SDFFX1 \fifo_reg[12][21]  ( .D(n755), .SI(\fifo[12][20] ), .SE(test_se), 
        .CLK(n27), .Q(\fifo[12][21] ), .QN(n1703) );
  SDFFX1 \fifo_reg[12][20]  ( .D(n754), .SI(\fifo[12][19] ), .SE(test_se), 
        .CLK(n27), .Q(\fifo[12][20] ), .QN(n1704) );
  SDFFX1 \fifo_reg[12][19]  ( .D(n753), .SI(\fifo[12][18] ), .SE(test_se), 
        .CLK(n27), .Q(\fifo[12][19] ), .QN(n1705) );
  SDFFX1 \fifo_reg[12][18]  ( .D(n752), .SI(\fifo[12][17] ), .SE(test_se), 
        .CLK(n27), .Q(\fifo[12][18] ), .QN(n1706) );
  SDFFX1 \fifo_reg[12][17]  ( .D(n751), .SI(\fifo[12][16] ), .SE(test_se), 
        .CLK(n27), .Q(\fifo[12][17] ), .QN(n1707) );
  SDFFX1 \fifo_reg[12][16]  ( .D(n750), .SI(\fifo[12][15] ), .SE(test_se), 
        .CLK(n27), .Q(\fifo[12][16] ), .QN(n1708) );
  SDFFX1 \fifo_reg[12][15]  ( .D(n749), .SI(\fifo[12][14] ), .SE(test_se), 
        .CLK(n27), .Q(\fifo[12][15] ), .QN(n1709) );
  SDFFX1 \fifo_reg[12][14]  ( .D(n748), .SI(\fifo[12][13] ), .SE(test_se), 
        .CLK(n27), .Q(\fifo[12][14] ), .QN(n1710) );
  SDFFX1 \fifo_reg[12][13]  ( .D(n747), .SI(\fifo[12][12] ), .SE(test_se), 
        .CLK(n26), .Q(\fifo[12][13] ), .QN(n1711) );
  SDFFX1 \fifo_reg[12][12]  ( .D(n746), .SI(\fifo[12][11] ), .SE(test_se), 
        .CLK(n26), .Q(\fifo[12][12] ), .QN(n1712) );
  SDFFX1 \fifo_reg[12][11]  ( .D(n745), .SI(\fifo[12][10] ), .SE(test_se), 
        .CLK(n26), .Q(\fifo[12][11] ), .QN(n1713) );
  SDFFX1 \fifo_reg[12][10]  ( .D(n744), .SI(\fifo[12][9] ), .SE(test_se), 
        .CLK(n26), .Q(\fifo[12][10] ), .QN(n1714) );
  SDFFX1 \fifo_reg[12][9]  ( .D(n743), .SI(\fifo[12][8] ), .SE(test_se), .CLK(
        n26), .Q(\fifo[12][9] ), .QN(n1715) );
  SDFFX1 \fifo_reg[12][8]  ( .D(n742), .SI(\fifo[12][7] ), .SE(test_se), .CLK(
        n26), .Q(\fifo[12][8] ), .QN(n1716) );
  SDFFX1 \fifo_reg[12][7]  ( .D(n741), .SI(\fifo[12][6] ), .SE(test_se), .CLK(
        n26), .Q(\fifo[12][7] ), .QN(n1717) );
  SDFFX1 \fifo_reg[12][6]  ( .D(n740), .SI(\fifo[12][5] ), .SE(test_se), .CLK(
        n26), .Q(\fifo[12][6] ), .QN(n1718) );
  SDFFX1 \fifo_reg[12][5]  ( .D(n739), .SI(\fifo[12][4] ), .SE(test_se), .CLK(
        n26), .Q(\fifo[12][5] ), .QN(n1719) );
  SDFFX1 \fifo_reg[12][4]  ( .D(n738), .SI(\fifo[12][3] ), .SE(test_se), .CLK(
        n26), .Q(\fifo[12][4] ), .QN(n1720) );
  SDFFX1 \fifo_reg[12][3]  ( .D(n737), .SI(\fifo[12][2] ), .SE(test_se), .CLK(
        n26), .Q(\fifo[12][3] ), .QN(n1721) );
  SDFFX1 \fifo_reg[12][2]  ( .D(n736), .SI(\fifo[12][1] ), .SE(test_se), .CLK(
        n26), .Q(\fifo[12][2] ), .QN(n1722) );
  SDFFX1 \fifo_reg[12][1]  ( .D(n735), .SI(\fifo[12][0] ), .SE(test_se), .CLK(
        n26), .Q(\fifo[12][1] ), .QN(n1723) );
  SDFFX1 \fifo_reg[12][0]  ( .D(n734), .SI(\fifo[11][31] ), .SE(test_se), 
        .CLK(n26), .Q(\fifo[12][0] ), .QN(n1724) );
  SDFFX1 \fifo_reg[13][31]  ( .D(n733), .SI(\fifo[13][30] ), .SE(test_se), 
        .CLK(n30), .Q(\fifo[13][31] ), .QN(n1725) );
  SDFFX1 \fifo_reg[13][30]  ( .D(n732), .SI(\fifo[13][29] ), .SE(test_se), 
        .CLK(n30), .Q(\fifo[13][30] ), .QN(n1726) );
  SDFFX1 \fifo_reg[13][29]  ( .D(n731), .SI(\fifo[13][28] ), .SE(test_se), 
        .CLK(n30), .Q(\fifo[13][29] ), .QN(n1727) );
  SDFFX1 \fifo_reg[13][28]  ( .D(n730), .SI(\fifo[13][27] ), .SE(test_se), 
        .CLK(n30), .Q(\fifo[13][28] ), .QN(n1728) );
  SDFFX1 \fifo_reg[13][27]  ( .D(n729), .SI(\fifo[13][26] ), .SE(test_se), 
        .CLK(n30), .Q(\fifo[13][27] ), .QN(n1729) );
  SDFFX1 \fifo_reg[13][26]  ( .D(n728), .SI(\fifo[13][25] ), .SE(test_se), 
        .CLK(n30), .Q(\fifo[13][26] ), .QN(n1730) );
  SDFFX1 \fifo_reg[13][25]  ( .D(n727), .SI(\fifo[13][24] ), .SE(test_se), 
        .CLK(n30), .Q(\fifo[13][25] ), .QN(n1731) );
  SDFFX1 \fifo_reg[13][24]  ( .D(n726), .SI(\fifo[13][23] ), .SE(test_se), 
        .CLK(n30), .Q(\fifo[13][24] ), .QN(n1732) );
  SDFFX1 \fifo_reg[13][23]  ( .D(n725), .SI(\fifo[13][22] ), .SE(test_se), 
        .CLK(n29), .Q(\fifo[13][23] ), .QN(n1733) );
  SDFFX1 \fifo_reg[13][22]  ( .D(n724), .SI(\fifo[13][21] ), .SE(test_se), 
        .CLK(n29), .Q(\fifo[13][22] ), .QN(n1734) );
  SDFFX1 \fifo_reg[13][21]  ( .D(n723), .SI(\fifo[13][20] ), .SE(test_se), 
        .CLK(n29), .Q(\fifo[13][21] ), .QN(n1735) );
  SDFFX1 \fifo_reg[13][20]  ( .D(n722), .SI(\fifo[13][19] ), .SE(test_se), 
        .CLK(n29), .Q(\fifo[13][20] ), .QN(n1736) );
  SDFFX1 \fifo_reg[13][19]  ( .D(n721), .SI(\fifo[13][18] ), .SE(test_se), 
        .CLK(n29), .Q(\fifo[13][19] ), .QN(n1737) );
  SDFFX1 \fifo_reg[13][18]  ( .D(n720), .SI(\fifo[13][17] ), .SE(test_se), 
        .CLK(n29), .Q(\fifo[13][18] ), .QN(n1738) );
  SDFFX1 \fifo_reg[13][17]  ( .D(n719), .SI(\fifo[13][16] ), .SE(test_se), 
        .CLK(n29), .Q(\fifo[13][17] ), .QN(n1739) );
  SDFFX1 \fifo_reg[13][16]  ( .D(n718), .SI(\fifo[13][15] ), .SE(test_se), 
        .CLK(n29), .Q(\fifo[13][16] ), .QN(n1740) );
  SDFFX1 \fifo_reg[13][15]  ( .D(n717), .SI(\fifo[13][14] ), .SE(test_se), 
        .CLK(n29), .Q(\fifo[13][15] ), .QN(n1741) );
  SDFFX1 \fifo_reg[13][14]  ( .D(n716), .SI(\fifo[13][13] ), .SE(test_se), 
        .CLK(n29), .Q(\fifo[13][14] ), .QN(n1742) );
  SDFFX1 \fifo_reg[13][13]  ( .D(n715), .SI(\fifo[13][12] ), .SE(test_se), 
        .CLK(n29), .Q(\fifo[13][13] ), .QN(n1743) );
  SDFFX1 \fifo_reg[13][12]  ( .D(n714), .SI(\fifo[13][11] ), .SE(test_se), 
        .CLK(n29), .Q(\fifo[13][12] ), .QN(n1744) );
  SDFFX1 \fifo_reg[13][11]  ( .D(n713), .SI(\fifo[13][10] ), .SE(test_se), 
        .CLK(n29), .Q(\fifo[13][11] ), .QN(n1745) );
  SDFFX1 \fifo_reg[13][10]  ( .D(n712), .SI(\fifo[13][9] ), .SE(test_se), 
        .CLK(n29), .Q(\fifo[13][10] ), .QN(n1746) );
  SDFFX1 \fifo_reg[13][9]  ( .D(n711), .SI(\fifo[13][8] ), .SE(test_se), .CLK(
        n28), .Q(\fifo[13][9] ), .QN(n1747) );
  SDFFX1 \fifo_reg[13][8]  ( .D(n710), .SI(\fifo[13][7] ), .SE(test_se), .CLK(
        n28), .Q(\fifo[13][8] ), .QN(n1748) );
  SDFFX1 \fifo_reg[13][7]  ( .D(n709), .SI(\fifo[13][6] ), .SE(test_se), .CLK(
        n28), .Q(\fifo[13][7] ), .QN(n1749) );
  SDFFX1 \fifo_reg[13][6]  ( .D(n708), .SI(\fifo[13][5] ), .SE(test_se), .CLK(
        n28), .Q(\fifo[13][6] ), .QN(n1750) );
  SDFFX1 \fifo_reg[13][5]  ( .D(n707), .SI(\fifo[13][4] ), .SE(test_se), .CLK(
        n28), .Q(\fifo[13][5] ), .QN(n1751) );
  SDFFX1 \fifo_reg[13][4]  ( .D(n706), .SI(\fifo[13][3] ), .SE(test_se), .CLK(
        n28), .Q(\fifo[13][4] ), .QN(n1752) );
  SDFFX1 \fifo_reg[13][3]  ( .D(n705), .SI(\fifo[13][2] ), .SE(test_se), .CLK(
        n28), .Q(\fifo[13][3] ), .QN(n1753) );
  SDFFX1 \fifo_reg[13][2]  ( .D(n704), .SI(\fifo[13][1] ), .SE(test_se), .CLK(
        n28), .Q(\fifo[13][2] ), .QN(n1754) );
  SDFFX1 \fifo_reg[13][1]  ( .D(n703), .SI(\fifo[13][0] ), .SE(test_se), .CLK(
        n28), .Q(\fifo[13][1] ), .QN(n1755) );
  SDFFX1 \fifo_reg[13][0]  ( .D(n702), .SI(\fifo[12][31] ), .SE(test_se), 
        .CLK(n28), .Q(\fifo[13][0] ), .QN(n1756) );
  SDFFX1 \fifo_reg[14][31]  ( .D(n701), .SI(\fifo[14][30] ), .SE(test_se), 
        .CLK(n32), .Q(\fifo[14][31] ), .QN(n1757) );
  SDFFX1 \fifo_reg[14][30]  ( .D(n700), .SI(\fifo[14][29] ), .SE(test_se), 
        .CLK(n32), .Q(\fifo[14][30] ), .QN(n1758) );
  SDFFX1 \fifo_reg[14][29]  ( .D(n699), .SI(\fifo[14][28] ), .SE(test_se), 
        .CLK(n32), .Q(\fifo[14][29] ), .QN(n1759) );
  SDFFX1 \fifo_reg[14][28]  ( .D(n698), .SI(\fifo[14][27] ), .SE(test_se), 
        .CLK(n32), .Q(\fifo[14][28] ), .QN(n1760) );
  SDFFX1 \fifo_reg[14][27]  ( .D(n697), .SI(\fifo[14][26] ), .SE(test_se), 
        .CLK(n32), .Q(\fifo[14][27] ), .QN(n1761) );
  SDFFX1 \fifo_reg[14][26]  ( .D(n696), .SI(\fifo[14][25] ), .SE(test_se), 
        .CLK(n32), .Q(\fifo[14][26] ), .QN(n1762) );
  SDFFX1 \fifo_reg[14][25]  ( .D(n695), .SI(\fifo[14][24] ), .SE(test_se), 
        .CLK(n32), .Q(\fifo[14][25] ), .QN(n1763) );
  SDFFX1 \fifo_reg[14][24]  ( .D(n694), .SI(\fifo[14][23] ), .SE(test_se), 
        .CLK(n32), .Q(\fifo[14][24] ), .QN(n1764) );
  SDFFX1 \fifo_reg[14][23]  ( .D(n693), .SI(\fifo[14][22] ), .SE(test_se), 
        .CLK(n32), .Q(\fifo[14][23] ), .QN(n1765) );
  SDFFX1 \fifo_reg[14][22]  ( .D(n692), .SI(\fifo[14][21] ), .SE(test_se), 
        .CLK(n32), .Q(\fifo[14][22] ), .QN(n1766) );
  SDFFX1 \fifo_reg[14][21]  ( .D(n691), .SI(\fifo[14][20] ), .SE(test_se), 
        .CLK(n32), .Q(\fifo[14][21] ), .QN(n1767) );
  SDFFX1 \fifo_reg[14][20]  ( .D(n690), .SI(\fifo[14][19] ), .SE(test_se), 
        .CLK(n32), .Q(\fifo[14][20] ), .QN(n1768) );
  SDFFX1 \fifo_reg[14][19]  ( .D(n689), .SI(\fifo[14][18] ), .SE(test_se), 
        .CLK(n32), .Q(\fifo[14][19] ), .QN(n1769) );
  SDFFX1 \fifo_reg[14][18]  ( .D(n688), .SI(\fifo[14][17] ), .SE(test_se), 
        .CLK(n31), .Q(\fifo[14][18] ), .QN(n1770) );
  SDFFX1 \fifo_reg[14][17]  ( .D(n687), .SI(\fifo[14][16] ), .SE(test_se), 
        .CLK(n31), .Q(\fifo[14][17] ), .QN(n1771) );
  SDFFX1 \fifo_reg[14][16]  ( .D(n686), .SI(\fifo[14][15] ), .SE(test_se), 
        .CLK(n31), .Q(\fifo[14][16] ), .QN(n1772) );
  SDFFX1 \fifo_reg[14][15]  ( .D(n685), .SI(\fifo[14][14] ), .SE(test_se), 
        .CLK(n31), .Q(\fifo[14][15] ), .QN(n1773) );
  SDFFX1 \fifo_reg[14][14]  ( .D(n684), .SI(\fifo[14][13] ), .SE(test_se), 
        .CLK(n31), .Q(\fifo[14][14] ), .QN(n1774) );
  SDFFX1 \fifo_reg[14][13]  ( .D(n683), .SI(\fifo[14][12] ), .SE(test_se), 
        .CLK(n31), .Q(\fifo[14][13] ), .QN(n1775) );
  SDFFX1 \fifo_reg[14][12]  ( .D(n682), .SI(\fifo[14][11] ), .SE(test_se), 
        .CLK(n31), .Q(\fifo[14][12] ), .QN(n1776) );
  SDFFX1 \fifo_reg[14][11]  ( .D(n681), .SI(\fifo[14][10] ), .SE(test_se), 
        .CLK(n31), .Q(\fifo[14][11] ), .QN(n1777) );
  SDFFX1 \fifo_reg[14][10]  ( .D(n680), .SI(\fifo[14][9] ), .SE(test_se), 
        .CLK(n31), .Q(\fifo[14][10] ), .QN(n1778) );
  SDFFX1 \fifo_reg[14][9]  ( .D(n679), .SI(\fifo[14][8] ), .SE(test_se), .CLK(
        n31), .Q(\fifo[14][9] ), .QN(n1779) );
  SDFFX1 \fifo_reg[14][8]  ( .D(n678), .SI(\fifo[14][7] ), .SE(test_se), .CLK(
        n31), .Q(\fifo[14][8] ), .QN(n1780) );
  SDFFX1 \fifo_reg[14][7]  ( .D(n677), .SI(\fifo[14][6] ), .SE(test_se), .CLK(
        n31), .Q(\fifo[14][7] ), .QN(n1781) );
  SDFFX1 \fifo_reg[14][6]  ( .D(n676), .SI(\fifo[14][5] ), .SE(test_se), .CLK(
        n31), .Q(\fifo[14][6] ), .QN(n1782) );
  SDFFX1 \fifo_reg[14][5]  ( .D(n675), .SI(\fifo[14][4] ), .SE(test_se), .CLK(
        n31), .Q(\fifo[14][5] ), .QN(n1783) );
  SDFFX1 \fifo_reg[14][4]  ( .D(n674), .SI(\fifo[14][3] ), .SE(test_se), .CLK(
        n30), .Q(\fifo[14][4] ), .QN(n1784) );
  SDFFX1 \fifo_reg[14][3]  ( .D(n673), .SI(\fifo[14][2] ), .SE(test_se), .CLK(
        n30), .Q(\fifo[14][3] ), .QN(n1785) );
  SDFFX1 \fifo_reg[14][2]  ( .D(n672), .SI(\fifo[14][1] ), .SE(test_se), .CLK(
        n30), .Q(\fifo[14][2] ), .QN(n1786) );
  SDFFX1 \fifo_reg[14][1]  ( .D(n671), .SI(\fifo[14][0] ), .SE(test_se), .CLK(
        n30), .Q(\fifo[14][1] ), .QN(n1787) );
  SDFFX1 \fifo_reg[14][0]  ( .D(n670), .SI(\fifo[13][31] ), .SE(test_se), 
        .CLK(n30), .Q(\fifo[14][0] ), .QN(n1788) );
  SDFFX1 \fifo_reg[15][31]  ( .D(n669), .SI(\fifo[15][30] ), .SE(test_se), 
        .CLK(n6), .Q(\fifo[15][31] ), .QN(n1789) );
  SDFFX1 \fifo_reg[15][30]  ( .D(n668), .SI(\fifo[15][29] ), .SE(test_se), 
        .CLK(n35), .Q(\fifo[15][30] ), .QN(n1790) );
  SDFFX1 \fifo_reg[15][29]  ( .D(n667), .SI(\fifo[15][28] ), .SE(test_se), 
        .CLK(n35), .Q(\fifo[15][29] ), .QN(n1791) );
  SDFFX1 \fifo_reg[15][28]  ( .D(n666), .SI(\fifo[15][27] ), .SE(test_se), 
        .CLK(n34), .Q(\fifo[15][28] ), .QN(n1792) );
  SDFFX1 \fifo_reg[15][27]  ( .D(n665), .SI(\fifo[15][26] ), .SE(test_se), 
        .CLK(n34), .Q(\fifo[15][27] ), .QN(n1793) );
  SDFFX1 \fifo_reg[15][26]  ( .D(n664), .SI(\fifo[15][25] ), .SE(test_se), 
        .CLK(n34), .Q(\fifo[15][26] ), .QN(n1794) );
  SDFFX1 \fifo_reg[15][25]  ( .D(n663), .SI(\fifo[15][24] ), .SE(test_se), 
        .CLK(n34), .Q(\fifo[15][25] ), .QN(n1795) );
  SDFFX1 \fifo_reg[15][24]  ( .D(n662), .SI(\fifo[15][23] ), .SE(test_se), 
        .CLK(n34), .Q(\fifo[15][24] ), .QN(n1796) );
  SDFFX1 \fifo_reg[15][23]  ( .D(n661), .SI(\fifo[15][22] ), .SE(test_se), 
        .CLK(n34), .Q(\fifo[15][23] ), .QN(n1797) );
  SDFFX1 \fifo_reg[15][22]  ( .D(n660), .SI(\fifo[15][21] ), .SE(test_se), 
        .CLK(n34), .Q(\fifo[15][22] ), .QN(n1798) );
  SDFFX1 \fifo_reg[15][21]  ( .D(n659), .SI(\fifo[15][20] ), .SE(test_se), 
        .CLK(n34), .Q(\fifo[15][21] ), .QN(n1799) );
  SDFFX1 \fifo_reg[15][20]  ( .D(n658), .SI(\fifo[15][19] ), .SE(test_se), 
        .CLK(n34), .Q(\fifo[15][20] ), .QN(n1800) );
  SDFFX1 \fifo_reg[15][19]  ( .D(n657), .SI(\fifo[15][18] ), .SE(test_se), 
        .CLK(n34), .Q(\fifo[15][19] ), .QN(n1801) );
  SDFFX1 \fifo_reg[15][18]  ( .D(n656), .SI(\fifo[15][17] ), .SE(test_se), 
        .CLK(n34), .Q(\fifo[15][18] ), .QN(n1802) );
  SDFFX1 \fifo_reg[15][17]  ( .D(n655), .SI(\fifo[15][16] ), .SE(test_se), 
        .CLK(n34), .Q(\fifo[15][17] ), .QN(n1803) );
  SDFFX1 \fifo_reg[15][16]  ( .D(n654), .SI(\fifo[15][15] ), .SE(test_se), 
        .CLK(n34), .Q(\fifo[15][16] ), .QN(n1804) );
  SDFFX1 \fifo_reg[15][15]  ( .D(n653), .SI(\fifo[15][14] ), .SE(test_se), 
        .CLK(n34), .Q(\fifo[15][15] ), .QN(n1805) );
  SDFFX1 \fifo_reg[15][14]  ( .D(n652), .SI(\fifo[15][13] ), .SE(test_se), 
        .CLK(n33), .Q(\fifo[15][14] ), .QN(n1806) );
  SDFFX1 \fifo_reg[15][13]  ( .D(n651), .SI(\fifo[15][12] ), .SE(test_se), 
        .CLK(n33), .Q(\fifo[15][13] ), .QN(n1807) );
  SDFFX1 \fifo_reg[15][12]  ( .D(n650), .SI(\fifo[15][11] ), .SE(test_se), 
        .CLK(n33), .Q(\fifo[15][12] ), .QN(n1808) );
  SDFFX1 \fifo_reg[15][11]  ( .D(n649), .SI(\fifo[15][10] ), .SE(test_se), 
        .CLK(n33), .Q(\fifo[15][11] ), .QN(n1809) );
  SDFFX1 \fifo_reg[15][10]  ( .D(n648), .SI(\fifo[15][9] ), .SE(test_se), 
        .CLK(n33), .Q(\fifo[15][10] ), .QN(n1810) );
  SDFFX1 \fifo_reg[15][9]  ( .D(n647), .SI(\fifo[15][8] ), .SE(test_se), .CLK(
        n33), .Q(\fifo[15][9] ), .QN(n1811) );
  SDFFX1 \fifo_reg[15][8]  ( .D(n646), .SI(\fifo[15][7] ), .SE(test_se), .CLK(
        n33), .Q(\fifo[15][8] ), .QN(n1812) );
  SDFFX1 \fifo_reg[15][7]  ( .D(n645), .SI(\fifo[15][6] ), .SE(test_se), .CLK(
        n33), .Q(\fifo[15][7] ), .QN(n1813) );
  SDFFX1 \fifo_reg[15][6]  ( .D(n644), .SI(\fifo[15][5] ), .SE(test_se), .CLK(
        n33), .Q(\fifo[15][6] ), .QN(n1814) );
  SDFFX1 \fifo_reg[15][5]  ( .D(n643), .SI(\fifo[15][4] ), .SE(test_se), .CLK(
        n33), .Q(\fifo[15][5] ), .QN(n1815) );
  SDFFX1 \fifo_reg[15][4]  ( .D(n642), .SI(\fifo[15][3] ), .SE(test_se), .CLK(
        n33), .Q(\fifo[15][4] ), .QN(n1816) );
  SDFFX1 \fifo_reg[15][3]  ( .D(n641), .SI(\fifo[15][2] ), .SE(test_se), .CLK(
        n33), .Q(\fifo[15][3] ), .QN(n1817) );
  SDFFX1 \fifo_reg[15][2]  ( .D(n640), .SI(\fifo[15][1] ), .SE(test_se), .CLK(
        n33), .Q(\fifo[15][2] ), .QN(n1818) );
  SDFFX1 \fifo_reg[15][1]  ( .D(n639), .SI(\fifo[15][0] ), .SE(test_se), .CLK(
        n33), .Q(\fifo[15][1] ), .QN(n1819) );
  SDFFX1 \fifo_reg[15][0]  ( .D(n638), .SI(\fifo[14][31] ), .SE(test_se), 
        .CLK(n32), .Q(\fifo[15][0] ), .QN(n1820) );
  SDFFX1 \data_out_reg[31]  ( .D(N155), .SI(data_out[30]), .SE(test_se), .CLK(
        n17), .Q(data_out[31]) );
  SDFFX1 \data_out_reg[30]  ( .D(N154), .SI(data_out[29]), .SE(test_se), .CLK(
        n17), .Q(data_out[30]) );
  SDFFX1 \data_out_reg[29]  ( .D(N153), .SI(data_out[28]), .SE(test_se), .CLK(
        n17), .Q(data_out[29]) );
  SDFFX1 \data_out_reg[28]  ( .D(N152), .SI(data_out[27]), .SE(test_se), .CLK(
        n17), .Q(data_out[28]) );
  SDFFX1 \data_out_reg[27]  ( .D(N151), .SI(data_out[26]), .SE(test_se), .CLK(
        n17), .Q(data_out[27]) );
  SDFFX1 \data_out_reg[26]  ( .D(N150), .SI(data_out[25]), .SE(test_se), .CLK(
        n17), .Q(data_out[26]) );
  SDFFX1 \data_out_reg[25]  ( .D(N149), .SI(data_out[24]), .SE(test_se), .CLK(
        n17), .Q(data_out[25]) );
  SDFFX1 \data_out_reg[24]  ( .D(N148), .SI(data_out[23]), .SE(test_se), .CLK(
        n17), .Q(data_out[24]) );
  SDFFX1 \data_out_reg[23]  ( .D(N147), .SI(data_out[22]), .SE(test_se), .CLK(
        n17), .Q(data_out[23]) );
  SDFFX1 \data_out_reg[22]  ( .D(N146), .SI(data_out[21]), .SE(test_se), .CLK(
        n17), .Q(data_out[22]) );
  SDFFX1 \data_out_reg[21]  ( .D(N145), .SI(data_out[20]), .SE(test_se), .CLK(
        n17), .Q(data_out[21]) );
  SDFFX1 \data_out_reg[20]  ( .D(N144), .SI(data_out[19]), .SE(test_se), .CLK(
        n17), .Q(data_out[20]) );
  SDFFX1 \data_out_reg[19]  ( .D(N143), .SI(data_out[18]), .SE(test_se), .CLK(
        n17), .Q(data_out[19]) );
  SDFFX1 \data_out_reg[18]  ( .D(N142), .SI(data_out[17]), .SE(test_se), .CLK(
        n16), .Q(data_out[18]) );
  SDFFX1 \data_out_reg[17]  ( .D(N141), .SI(data_out[16]), .SE(test_se), .CLK(
        n16), .Q(data_out[17]) );
  SDFFX1 \data_out_reg[16]  ( .D(N140), .SI(data_out[15]), .SE(test_se), .CLK(
        n16), .Q(data_out[16]) );
  SDFFX1 \data_out_reg[15]  ( .D(N139), .SI(data_out[14]), .SE(test_se), .CLK(
        n16), .Q(data_out[15]) );
  SDFFX1 \data_out_reg[14]  ( .D(N138), .SI(data_out[13]), .SE(test_se), .CLK(
        n16), .Q(data_out[14]) );
  SDFFX1 \data_out_reg[13]  ( .D(N137), .SI(data_out[12]), .SE(test_se), .CLK(
        n16), .Q(data_out[13]) );
  SDFFX1 \data_out_reg[12]  ( .D(N136), .SI(data_out[11]), .SE(test_se), .CLK(
        n16), .Q(data_out[12]) );
  SDFFX1 \data_out_reg[11]  ( .D(N135), .SI(data_out[10]), .SE(test_se), .CLK(
        n16), .Q(data_out[11]) );
  SDFFX1 \data_out_reg[10]  ( .D(N134), .SI(data_out[9]), .SE(test_se), .CLK(
        n16), .Q(data_out[10]) );
  SDFFX1 \data_out_reg[9]  ( .D(N133), .SI(data_out[8]), .SE(test_se), .CLK(
        n16), .Q(data_out[9]) );
  SDFFX1 \data_out_reg[8]  ( .D(N132), .SI(data_out[7]), .SE(test_se), .CLK(
        n16), .Q(data_out[8]) );
  SDFFX1 \data_out_reg[7]  ( .D(N131), .SI(data_out[6]), .SE(test_se), .CLK(
        n16), .Q(data_out[7]) );
  SDFFX1 \data_out_reg[6]  ( .D(N130), .SI(data_out[5]), .SE(test_se), .CLK(
        n16), .Q(data_out[6]) );
  SDFFX1 \data_out_reg[5]  ( .D(N129), .SI(data_out[4]), .SE(test_se), .CLK(
        n16), .Q(data_out[5]) );
  SDFFX1 \data_out_reg[4]  ( .D(N128), .SI(data_out[3]), .SE(test_se), .CLK(
        n15), .Q(data_out[4]) );
  SDFFX1 \data_out_reg[3]  ( .D(N127), .SI(data_out[2]), .SE(test_se), .CLK(
        n15), .Q(data_out[3]) );
  SDFFX1 \data_out_reg[2]  ( .D(N126), .SI(data_out[1]), .SE(test_se), .CLK(
        n15), .Q(data_out[2]) );
  SDFFX1 \data_out_reg[1]  ( .D(N125), .SI(data_out[0]), .SE(test_se), .CLK(
        n15), .Q(data_out[1]) );
  SDFFX1 \data_out_reg[0]  ( .D(N124), .SI(cnt[4]), .SE(test_se), .CLK(n20), 
        .Q(data_out[0]) );
  NBUFFX2 U3 ( .INP(clk), .Z(n6) );
  NBUFFX2 U4 ( .INP(clk), .Z(n16) );
  NBUFFX2 U5 ( .INP(clk), .Z(n33) );
  NBUFFX2 U6 ( .INP(clk), .Z(n34) );
  NBUFFX2 U7 ( .INP(clk), .Z(n31) );
  NBUFFX2 U8 ( .INP(clk), .Z(n32) );
  NBUFFX2 U9 ( .INP(clk), .Z(n29) );
  NBUFFX2 U10 ( .INP(clk), .Z(n26) );
  NBUFFX2 U11 ( .INP(clk), .Z(n27) );
  NBUFFX2 U12 ( .INP(clk), .Z(n28) );
  NBUFFX2 U13 ( .INP(clk), .Z(n30) );
  NBUFFX2 U14 ( .INP(clk), .Z(n42) );
  NBUFFX2 U15 ( .INP(clk), .Z(n43) );
  NBUFFX2 U16 ( .INP(clk), .Z(n39) );
  NBUFFX2 U17 ( .INP(clk), .Z(n41) );
  NBUFFX2 U18 ( .INP(clk), .Z(n37) );
  NBUFFX2 U19 ( .INP(clk), .Z(n38) );
  NBUFFX2 U20 ( .INP(clk), .Z(n15) );
  NBUFFX2 U21 ( .INP(clk), .Z(n40) );
  NBUFFX2 U22 ( .INP(clk), .Z(n35) );
  NBUFFX2 U23 ( .INP(clk), .Z(n36) );
  NBUFFX2 U24 ( .INP(clk), .Z(n13) );
  NBUFFX2 U25 ( .INP(clk), .Z(n14) );
  NBUFFX2 U26 ( .INP(clk), .Z(n11) );
  NBUFFX2 U27 ( .INP(clk), .Z(n12) );
  NBUFFX2 U28 ( .INP(clk), .Z(n9) );
  NBUFFX2 U29 ( .INP(clk), .Z(n10) );
  NBUFFX2 U30 ( .INP(clk), .Z(n25) );
  NBUFFX2 U31 ( .INP(clk), .Z(n8) );
  NBUFFX2 U32 ( .INP(clk), .Z(n7) );
  NBUFFX2 U33 ( .INP(clk), .Z(n23) );
  NBUFFX2 U34 ( .INP(clk), .Z(n24) );
  NBUFFX2 U35 ( .INP(clk), .Z(n21) );
  NBUFFX2 U36 ( .INP(clk), .Z(n22) );
  NBUFFX2 U37 ( .INP(clk), .Z(n17) );
  NBUFFX2 U38 ( .INP(clk), .Z(n18) );
  NBUFFX2 U39 ( .INP(clk), .Z(n19) );
  NBUFFX2 U40 ( .INP(clk), .Z(n20) );
  NBUFFX2 U41 ( .INP(clk), .Z(n5) );
  NBUFFX2 U42 ( .INP(clk), .Z(n44) );
  INVX0 U43 ( .INP(n45), .ZN(empty) );
  INVX0 U44 ( .INP(n46), .ZN(full) );
  INVX0 U45 ( .INP(eth_top_test_point_11887_in), .ZN(n428) );
  MUX21X1 U46 ( .IN1(\fifo[4][9] ), .IN2(data_in[9]), .S(n47), .Q(n999) );
  MUX21X1 U47 ( .IN1(\fifo[4][8] ), .IN2(data_in[8]), .S(n47), .Q(n998) );
  MUX21X1 U48 ( .IN1(\fifo[4][7] ), .IN2(data_in[7]), .S(n47), .Q(n997) );
  MUX21X1 U49 ( .IN1(\fifo[4][6] ), .IN2(data_in[6]), .S(n47), .Q(n996) );
  MUX21X1 U50 ( .IN1(\fifo[4][5] ), .IN2(data_in[5]), .S(n47), .Q(n995) );
  MUX21X1 U51 ( .IN1(\fifo[4][4] ), .IN2(data_in[4]), .S(n47), .Q(n994) );
  MUX21X1 U52 ( .IN1(\fifo[4][3] ), .IN2(data_in[3]), .S(n47), .Q(n993) );
  MUX21X1 U53 ( .IN1(\fifo[4][2] ), .IN2(data_in[2]), .S(n47), .Q(n992) );
  MUX21X1 U54 ( .IN1(\fifo[4][1] ), .IN2(data_in[1]), .S(n47), .Q(n991) );
  MUX21X1 U55 ( .IN1(\fifo[4][0] ), .IN2(data_in[0]), .S(n47), .Q(n990) );
  MUX21X1 U56 ( .IN1(\fifo[5][31] ), .IN2(data_in[31]), .S(n48), .Q(n989) );
  MUX21X1 U57 ( .IN1(\fifo[5][30] ), .IN2(data_in[30]), .S(n48), .Q(n988) );
  MUX21X1 U58 ( .IN1(\fifo[5][29] ), .IN2(data_in[29]), .S(n48), .Q(n987) );
  MUX21X1 U59 ( .IN1(\fifo[5][28] ), .IN2(data_in[28]), .S(n48), .Q(n986) );
  MUX21X1 U60 ( .IN1(\fifo[5][27] ), .IN2(data_in[27]), .S(n48), .Q(n985) );
  MUX21X1 U61 ( .IN1(\fifo[5][26] ), .IN2(data_in[26]), .S(n48), .Q(n984) );
  MUX21X1 U62 ( .IN1(\fifo[5][25] ), .IN2(data_in[25]), .S(n48), .Q(n983) );
  MUX21X1 U63 ( .IN1(\fifo[5][24] ), .IN2(data_in[24]), .S(n48), .Q(n982) );
  MUX21X1 U64 ( .IN1(\fifo[5][23] ), .IN2(data_in[23]), .S(n48), .Q(n981) );
  MUX21X1 U65 ( .IN1(\fifo[5][22] ), .IN2(data_in[22]), .S(n48), .Q(n980) );
  MUX21X1 U66 ( .IN1(\fifo[5][21] ), .IN2(data_in[21]), .S(n48), .Q(n979) );
  MUX21X1 U67 ( .IN1(\fifo[5][20] ), .IN2(data_in[20]), .S(n48), .Q(n978) );
  MUX21X1 U68 ( .IN1(\fifo[5][19] ), .IN2(data_in[19]), .S(n48), .Q(n977) );
  MUX21X1 U69 ( .IN1(\fifo[5][18] ), .IN2(data_in[18]), .S(n48), .Q(n976) );
  MUX21X1 U70 ( .IN1(\fifo[5][17] ), .IN2(data_in[17]), .S(n48), .Q(n975) );
  MUX21X1 U71 ( .IN1(\fifo[5][16] ), .IN2(data_in[16]), .S(n48), .Q(n974) );
  MUX21X1 U72 ( .IN1(\fifo[5][15] ), .IN2(data_in[15]), .S(n48), .Q(n973) );
  MUX21X1 U73 ( .IN1(\fifo[5][14] ), .IN2(data_in[14]), .S(n48), .Q(n972) );
  MUX21X1 U74 ( .IN1(\fifo[5][13] ), .IN2(data_in[13]), .S(n48), .Q(n971) );
  MUX21X1 U75 ( .IN1(\fifo[5][12] ), .IN2(data_in[12]), .S(n48), .Q(n970) );
  MUX21X1 U76 ( .IN1(\fifo[5][11] ), .IN2(data_in[11]), .S(n48), .Q(n969) );
  MUX21X1 U77 ( .IN1(\fifo[5][10] ), .IN2(data_in[10]), .S(n48), .Q(n968) );
  MUX21X1 U78 ( .IN1(\fifo[5][9] ), .IN2(data_in[9]), .S(n48), .Q(n967) );
  MUX21X1 U79 ( .IN1(\fifo[5][8] ), .IN2(data_in[8]), .S(n48), .Q(n966) );
  MUX21X1 U80 ( .IN1(\fifo[5][7] ), .IN2(data_in[7]), .S(n48), .Q(n965) );
  MUX21X1 U81 ( .IN1(\fifo[5][6] ), .IN2(data_in[6]), .S(n48), .Q(n964) );
  MUX21X1 U82 ( .IN1(\fifo[5][5] ), .IN2(data_in[5]), .S(n48), .Q(n963) );
  MUX21X1 U83 ( .IN1(\fifo[5][4] ), .IN2(data_in[4]), .S(n48), .Q(n962) );
  MUX21X1 U84 ( .IN1(\fifo[5][3] ), .IN2(data_in[3]), .S(n48), .Q(n961) );
  MUX21X1 U85 ( .IN1(\fifo[5][2] ), .IN2(data_in[2]), .S(n48), .Q(n960) );
  MUX21X1 U86 ( .IN1(\fifo[5][1] ), .IN2(data_in[1]), .S(n48), .Q(n959) );
  MUX21X1 U87 ( .IN1(\fifo[5][0] ), .IN2(data_in[0]), .S(n48), .Q(n958) );
  AND2X1 U88 ( .IN1(n49), .IN2(n50), .Q(n48) );
  MUX21X1 U89 ( .IN1(\fifo[6][31] ), .IN2(data_in[31]), .S(n51), .Q(n957) );
  MUX21X1 U90 ( .IN1(\fifo[6][30] ), .IN2(data_in[30]), .S(n51), .Q(n956) );
  MUX21X1 U91 ( .IN1(\fifo[6][29] ), .IN2(data_in[29]), .S(n51), .Q(n955) );
  MUX21X1 U92 ( .IN1(\fifo[6][28] ), .IN2(data_in[28]), .S(n51), .Q(n954) );
  MUX21X1 U93 ( .IN1(\fifo[6][27] ), .IN2(data_in[27]), .S(n51), .Q(n953) );
  MUX21X1 U94 ( .IN1(\fifo[6][26] ), .IN2(data_in[26]), .S(n51), .Q(n952) );
  MUX21X1 U95 ( .IN1(\fifo[6][25] ), .IN2(data_in[25]), .S(n51), .Q(n951) );
  MUX21X1 U96 ( .IN1(\fifo[6][24] ), .IN2(data_in[24]), .S(n51), .Q(n950) );
  MUX21X1 U97 ( .IN1(\fifo[6][23] ), .IN2(data_in[23]), .S(n51), .Q(n949) );
  MUX21X1 U98 ( .IN1(\fifo[6][22] ), .IN2(data_in[22]), .S(n51), .Q(n948) );
  MUX21X1 U99 ( .IN1(\fifo[6][21] ), .IN2(data_in[21]), .S(n51), .Q(n947) );
  MUX21X1 U100 ( .IN1(\fifo[6][20] ), .IN2(data_in[20]), .S(n51), .Q(n946) );
  MUX21X1 U101 ( .IN1(\fifo[6][19] ), .IN2(data_in[19]), .S(n51), .Q(n945) );
  MUX21X1 U102 ( .IN1(\fifo[6][18] ), .IN2(data_in[18]), .S(n51), .Q(n944) );
  MUX21X1 U103 ( .IN1(\fifo[6][17] ), .IN2(data_in[17]), .S(n51), .Q(n943) );
  MUX21X1 U104 ( .IN1(\fifo[6][16] ), .IN2(data_in[16]), .S(n51), .Q(n942) );
  MUX21X1 U105 ( .IN1(\fifo[6][15] ), .IN2(data_in[15]), .S(n51), .Q(n941) );
  MUX21X1 U106 ( .IN1(\fifo[6][14] ), .IN2(data_in[14]), .S(n51), .Q(n940) );
  MUX21X1 U107 ( .IN1(\fifo[6][13] ), .IN2(data_in[13]), .S(n51), .Q(n939) );
  MUX21X1 U108 ( .IN1(\fifo[6][12] ), .IN2(data_in[12]), .S(n51), .Q(n938) );
  MUX21X1 U109 ( .IN1(\fifo[6][11] ), .IN2(data_in[11]), .S(n51), .Q(n937) );
  MUX21X1 U110 ( .IN1(\fifo[6][10] ), .IN2(data_in[10]), .S(n51), .Q(n936) );
  MUX21X1 U111 ( .IN1(\fifo[6][9] ), .IN2(data_in[9]), .S(n51), .Q(n935) );
  MUX21X1 U112 ( .IN1(\fifo[6][8] ), .IN2(data_in[8]), .S(n51), .Q(n934) );
  MUX21X1 U113 ( .IN1(\fifo[6][7] ), .IN2(data_in[7]), .S(n51), .Q(n933) );
  MUX21X1 U114 ( .IN1(\fifo[6][6] ), .IN2(data_in[6]), .S(n51), .Q(n932) );
  MUX21X1 U115 ( .IN1(\fifo[6][5] ), .IN2(data_in[5]), .S(n51), .Q(n931) );
  MUX21X1 U116 ( .IN1(\fifo[6][4] ), .IN2(data_in[4]), .S(n51), .Q(n930) );
  MUX21X1 U117 ( .IN1(\fifo[6][3] ), .IN2(data_in[3]), .S(n51), .Q(n929) );
  MUX21X1 U118 ( .IN1(\fifo[6][2] ), .IN2(data_in[2]), .S(n51), .Q(n928) );
  MUX21X1 U119 ( .IN1(\fifo[6][1] ), .IN2(data_in[1]), .S(n51), .Q(n927) );
  MUX21X1 U120 ( .IN1(\fifo[6][0] ), .IN2(data_in[0]), .S(n51), .Q(n926) );
  AND2X1 U121 ( .IN1(n52), .IN2(n50), .Q(n51) );
  MUX21X1 U122 ( .IN1(\fifo[7][31] ), .IN2(data_in[31]), .S(n53), .Q(n925) );
  MUX21X1 U123 ( .IN1(\fifo[7][30] ), .IN2(data_in[30]), .S(n53), .Q(n924) );
  MUX21X1 U124 ( .IN1(\fifo[7][29] ), .IN2(data_in[29]), .S(n53), .Q(n923) );
  MUX21X1 U125 ( .IN1(\fifo[7][28] ), .IN2(data_in[28]), .S(n53), .Q(n922) );
  MUX21X1 U126 ( .IN1(\fifo[7][27] ), .IN2(data_in[27]), .S(n53), .Q(n921) );
  MUX21X1 U127 ( .IN1(\fifo[7][26] ), .IN2(data_in[26]), .S(n53), .Q(n920) );
  MUX21X1 U128 ( .IN1(\fifo[7][25] ), .IN2(data_in[25]), .S(n53), .Q(n919) );
  MUX21X1 U129 ( .IN1(\fifo[7][24] ), .IN2(data_in[24]), .S(n53), .Q(n918) );
  MUX21X1 U130 ( .IN1(\fifo[7][23] ), .IN2(data_in[23]), .S(n53), .Q(n917) );
  MUX21X1 U131 ( .IN1(\fifo[7][22] ), .IN2(data_in[22]), .S(n53), .Q(n916) );
  MUX21X1 U132 ( .IN1(\fifo[7][21] ), .IN2(data_in[21]), .S(n53), .Q(n915) );
  MUX21X1 U133 ( .IN1(\fifo[7][20] ), .IN2(data_in[20]), .S(n53), .Q(n914) );
  MUX21X1 U134 ( .IN1(\fifo[7][19] ), .IN2(data_in[19]), .S(n53), .Q(n913) );
  MUX21X1 U135 ( .IN1(\fifo[7][18] ), .IN2(data_in[18]), .S(n53), .Q(n912) );
  MUX21X1 U136 ( .IN1(\fifo[7][17] ), .IN2(data_in[17]), .S(n53), .Q(n911) );
  MUX21X1 U137 ( .IN1(\fifo[7][16] ), .IN2(data_in[16]), .S(n53), .Q(n910) );
  MUX21X1 U138 ( .IN1(\fifo[7][15] ), .IN2(data_in[15]), .S(n53), .Q(n909) );
  MUX21X1 U139 ( .IN1(\fifo[7][14] ), .IN2(data_in[14]), .S(n53), .Q(n908) );
  MUX21X1 U140 ( .IN1(\fifo[7][13] ), .IN2(data_in[13]), .S(n53), .Q(n907) );
  MUX21X1 U141 ( .IN1(\fifo[7][12] ), .IN2(data_in[12]), .S(n53), .Q(n906) );
  MUX21X1 U142 ( .IN1(\fifo[7][11] ), .IN2(data_in[11]), .S(n53), .Q(n905) );
  MUX21X1 U143 ( .IN1(\fifo[7][10] ), .IN2(data_in[10]), .S(n53), .Q(n904) );
  MUX21X1 U144 ( .IN1(\fifo[7][9] ), .IN2(data_in[9]), .S(n53), .Q(n903) );
  MUX21X1 U145 ( .IN1(\fifo[7][8] ), .IN2(data_in[8]), .S(n53), .Q(n902) );
  MUX21X1 U146 ( .IN1(\fifo[7][7] ), .IN2(data_in[7]), .S(n53), .Q(n901) );
  MUX21X1 U147 ( .IN1(\fifo[7][6] ), .IN2(data_in[6]), .S(n53), .Q(n900) );
  MUX21X1 U148 ( .IN1(\fifo[7][5] ), .IN2(data_in[5]), .S(n53), .Q(n899) );
  MUX21X1 U149 ( .IN1(\fifo[7][4] ), .IN2(data_in[4]), .S(n53), .Q(n898) );
  MUX21X1 U150 ( .IN1(\fifo[7][3] ), .IN2(data_in[3]), .S(n53), .Q(n897) );
  MUX21X1 U151 ( .IN1(\fifo[7][2] ), .IN2(data_in[2]), .S(n53), .Q(n896) );
  MUX21X1 U152 ( .IN1(\fifo[7][1] ), .IN2(data_in[1]), .S(n53), .Q(n895) );
  MUX21X1 U153 ( .IN1(\fifo[7][0] ), .IN2(data_in[0]), .S(n53), .Q(n894) );
  MUX21X1 U154 ( .IN1(\fifo[8][31] ), .IN2(data_in[31]), .S(n54), .Q(n893) );
  MUX21X1 U155 ( .IN1(\fifo[8][30] ), .IN2(data_in[30]), .S(n54), .Q(n892) );
  MUX21X1 U156 ( .IN1(\fifo[8][29] ), .IN2(data_in[29]), .S(n54), .Q(n891) );
  MUX21X1 U157 ( .IN1(\fifo[8][28] ), .IN2(data_in[28]), .S(n54), .Q(n890) );
  MUX21X1 U158 ( .IN1(\fifo[8][27] ), .IN2(data_in[27]), .S(n54), .Q(n889) );
  MUX21X1 U159 ( .IN1(\fifo[8][26] ), .IN2(data_in[26]), .S(n54), .Q(n888) );
  MUX21X1 U160 ( .IN1(\fifo[8][25] ), .IN2(data_in[25]), .S(n54), .Q(n887) );
  MUX21X1 U161 ( .IN1(\fifo[8][24] ), .IN2(data_in[24]), .S(n54), .Q(n886) );
  MUX21X1 U162 ( .IN1(\fifo[8][23] ), .IN2(data_in[23]), .S(n54), .Q(n885) );
  MUX21X1 U163 ( .IN1(\fifo[8][22] ), .IN2(data_in[22]), .S(n54), .Q(n884) );
  MUX21X1 U164 ( .IN1(\fifo[8][21] ), .IN2(data_in[21]), .S(n54), .Q(n883) );
  MUX21X1 U165 ( .IN1(\fifo[8][20] ), .IN2(data_in[20]), .S(n54), .Q(n882) );
  MUX21X1 U166 ( .IN1(\fifo[8][19] ), .IN2(data_in[19]), .S(n54), .Q(n881) );
  MUX21X1 U167 ( .IN1(\fifo[8][18] ), .IN2(data_in[18]), .S(n54), .Q(n880) );
  MUX21X1 U168 ( .IN1(\fifo[8][17] ), .IN2(data_in[17]), .S(n54), .Q(n879) );
  MUX21X1 U169 ( .IN1(\fifo[8][16] ), .IN2(data_in[16]), .S(n54), .Q(n878) );
  MUX21X1 U170 ( .IN1(\fifo[8][15] ), .IN2(data_in[15]), .S(n54), .Q(n877) );
  MUX21X1 U171 ( .IN1(\fifo[8][14] ), .IN2(data_in[14]), .S(n54), .Q(n876) );
  MUX21X1 U172 ( .IN1(\fifo[8][13] ), .IN2(data_in[13]), .S(n54), .Q(n875) );
  MUX21X1 U173 ( .IN1(\fifo[8][12] ), .IN2(data_in[12]), .S(n54), .Q(n874) );
  MUX21X1 U174 ( .IN1(\fifo[8][11] ), .IN2(data_in[11]), .S(n54), .Q(n873) );
  MUX21X1 U175 ( .IN1(\fifo[8][10] ), .IN2(data_in[10]), .S(n54), .Q(n872) );
  MUX21X1 U176 ( .IN1(\fifo[8][9] ), .IN2(data_in[9]), .S(n54), .Q(n871) );
  MUX21X1 U177 ( .IN1(\fifo[8][8] ), .IN2(data_in[8]), .S(n54), .Q(n870) );
  MUX21X1 U178 ( .IN1(\fifo[8][7] ), .IN2(data_in[7]), .S(n54), .Q(n869) );
  MUX21X1 U179 ( .IN1(\fifo[8][6] ), .IN2(data_in[6]), .S(n54), .Q(n868) );
  MUX21X1 U180 ( .IN1(\fifo[8][5] ), .IN2(data_in[5]), .S(n54), .Q(n867) );
  MUX21X1 U181 ( .IN1(\fifo[8][4] ), .IN2(data_in[4]), .S(n54), .Q(n866) );
  MUX21X1 U182 ( .IN1(\fifo[8][3] ), .IN2(data_in[3]), .S(n54), .Q(n865) );
  MUX21X1 U183 ( .IN1(\fifo[8][2] ), .IN2(data_in[2]), .S(n54), .Q(n864) );
  MUX21X1 U184 ( .IN1(\fifo[8][1] ), .IN2(data_in[1]), .S(n54), .Q(n863) );
  MUX21X1 U185 ( .IN1(\fifo[8][0] ), .IN2(data_in[0]), .S(n54), .Q(n862) );
  AND2X1 U186 ( .IN1(n55), .IN2(n56), .Q(n54) );
  MUX21X1 U187 ( .IN1(\fifo[9][31] ), .IN2(data_in[31]), .S(n57), .Q(n861) );
  MUX21X1 U188 ( .IN1(\fifo[9][30] ), .IN2(data_in[30]), .S(n57), .Q(n860) );
  MUX21X1 U189 ( .IN1(\fifo[9][29] ), .IN2(data_in[29]), .S(n57), .Q(n859) );
  MUX21X1 U190 ( .IN1(\fifo[9][28] ), .IN2(data_in[28]), .S(n57), .Q(n858) );
  MUX21X1 U191 ( .IN1(\fifo[9][27] ), .IN2(data_in[27]), .S(n57), .Q(n857) );
  MUX21X1 U192 ( .IN1(\fifo[9][26] ), .IN2(data_in[26]), .S(n57), .Q(n856) );
  MUX21X1 U193 ( .IN1(\fifo[9][25] ), .IN2(data_in[25]), .S(n57), .Q(n855) );
  MUX21X1 U194 ( .IN1(\fifo[9][24] ), .IN2(data_in[24]), .S(n57), .Q(n854) );
  MUX21X1 U195 ( .IN1(\fifo[9][23] ), .IN2(data_in[23]), .S(n57), .Q(n853) );
  MUX21X1 U196 ( .IN1(\fifo[9][22] ), .IN2(data_in[22]), .S(n57), .Q(n852) );
  MUX21X1 U197 ( .IN1(\fifo[9][21] ), .IN2(data_in[21]), .S(n57), .Q(n851) );
  MUX21X1 U198 ( .IN1(\fifo[9][20] ), .IN2(data_in[20]), .S(n57), .Q(n850) );
  MUX21X1 U199 ( .IN1(\fifo[9][19] ), .IN2(data_in[19]), .S(n57), .Q(n849) );
  MUX21X1 U200 ( .IN1(\fifo[9][18] ), .IN2(data_in[18]), .S(n57), .Q(n848) );
  MUX21X1 U201 ( .IN1(\fifo[9][17] ), .IN2(data_in[17]), .S(n57), .Q(n847) );
  MUX21X1 U202 ( .IN1(\fifo[9][16] ), .IN2(data_in[16]), .S(n57), .Q(n846) );
  MUX21X1 U203 ( .IN1(\fifo[9][15] ), .IN2(data_in[15]), .S(n57), .Q(n845) );
  MUX21X1 U204 ( .IN1(\fifo[9][14] ), .IN2(data_in[14]), .S(n57), .Q(n844) );
  MUX21X1 U205 ( .IN1(\fifo[9][13] ), .IN2(data_in[13]), .S(n57), .Q(n843) );
  MUX21X1 U206 ( .IN1(\fifo[9][12] ), .IN2(data_in[12]), .S(n57), .Q(n842) );
  MUX21X1 U207 ( .IN1(\fifo[9][11] ), .IN2(data_in[11]), .S(n57), .Q(n841) );
  MUX21X1 U208 ( .IN1(\fifo[9][10] ), .IN2(data_in[10]), .S(n57), .Q(n840) );
  MUX21X1 U209 ( .IN1(\fifo[9][9] ), .IN2(data_in[9]), .S(n57), .Q(n839) );
  MUX21X1 U210 ( .IN1(\fifo[9][8] ), .IN2(data_in[8]), .S(n57), .Q(n838) );
  MUX21X1 U211 ( .IN1(\fifo[9][7] ), .IN2(data_in[7]), .S(n57), .Q(n837) );
  MUX21X1 U212 ( .IN1(\fifo[9][6] ), .IN2(data_in[6]), .S(n57), .Q(n836) );
  MUX21X1 U213 ( .IN1(\fifo[9][5] ), .IN2(data_in[5]), .S(n57), .Q(n835) );
  MUX21X1 U214 ( .IN1(\fifo[9][4] ), .IN2(data_in[4]), .S(n57), .Q(n834) );
  MUX21X1 U215 ( .IN1(\fifo[9][3] ), .IN2(data_in[3]), .S(n57), .Q(n833) );
  MUX21X1 U216 ( .IN1(\fifo[9][2] ), .IN2(data_in[2]), .S(n57), .Q(n832) );
  MUX21X1 U217 ( .IN1(\fifo[9][1] ), .IN2(data_in[1]), .S(n57), .Q(n831) );
  MUX21X1 U218 ( .IN1(\fifo[9][0] ), .IN2(data_in[0]), .S(n57), .Q(n830) );
  AND2X1 U219 ( .IN1(n55), .IN2(n49), .Q(n57) );
  MUX21X1 U220 ( .IN1(\fifo[10][31] ), .IN2(data_in[31]), .S(n58), .Q(n829) );
  MUX21X1 U221 ( .IN1(\fifo[10][30] ), .IN2(data_in[30]), .S(n58), .Q(n828) );
  MUX21X1 U222 ( .IN1(\fifo[10][29] ), .IN2(data_in[29]), .S(n58), .Q(n827) );
  MUX21X1 U223 ( .IN1(\fifo[10][28] ), .IN2(data_in[28]), .S(n58), .Q(n826) );
  MUX21X1 U224 ( .IN1(\fifo[10][27] ), .IN2(data_in[27]), .S(n58), .Q(n825) );
  MUX21X1 U225 ( .IN1(\fifo[10][26] ), .IN2(data_in[26]), .S(n58), .Q(n824) );
  MUX21X1 U226 ( .IN1(\fifo[10][25] ), .IN2(data_in[25]), .S(n58), .Q(n823) );
  MUX21X1 U227 ( .IN1(\fifo[10][24] ), .IN2(data_in[24]), .S(n58), .Q(n822) );
  MUX21X1 U228 ( .IN1(\fifo[10][23] ), .IN2(data_in[23]), .S(n58), .Q(n821) );
  MUX21X1 U229 ( .IN1(\fifo[10][22] ), .IN2(data_in[22]), .S(n58), .Q(n820) );
  MUX21X1 U230 ( .IN1(\fifo[10][21] ), .IN2(data_in[21]), .S(n58), .Q(n819) );
  MUX21X1 U231 ( .IN1(\fifo[10][20] ), .IN2(data_in[20]), .S(n58), .Q(n818) );
  MUX21X1 U232 ( .IN1(\fifo[10][19] ), .IN2(data_in[19]), .S(n58), .Q(n817) );
  MUX21X1 U233 ( .IN1(\fifo[10][18] ), .IN2(data_in[18]), .S(n58), .Q(n816) );
  MUX21X1 U234 ( .IN1(\fifo[10][17] ), .IN2(data_in[17]), .S(n58), .Q(n815) );
  MUX21X1 U235 ( .IN1(\fifo[10][16] ), .IN2(data_in[16]), .S(n58), .Q(n814) );
  MUX21X1 U236 ( .IN1(\fifo[10][15] ), .IN2(data_in[15]), .S(n58), .Q(n813) );
  MUX21X1 U237 ( .IN1(\fifo[10][14] ), .IN2(data_in[14]), .S(n58), .Q(n812) );
  MUX21X1 U238 ( .IN1(\fifo[10][13] ), .IN2(data_in[13]), .S(n58), .Q(n811) );
  MUX21X1 U239 ( .IN1(\fifo[10][12] ), .IN2(data_in[12]), .S(n58), .Q(n810) );
  MUX21X1 U240 ( .IN1(\fifo[10][11] ), .IN2(data_in[11]), .S(n58), .Q(n809) );
  MUX21X1 U241 ( .IN1(\fifo[10][10] ), .IN2(data_in[10]), .S(n58), .Q(n808) );
  MUX21X1 U242 ( .IN1(\fifo[10][9] ), .IN2(data_in[9]), .S(n58), .Q(n807) );
  MUX21X1 U243 ( .IN1(\fifo[10][8] ), .IN2(data_in[8]), .S(n58), .Q(n806) );
  MUX21X1 U244 ( .IN1(\fifo[10][7] ), .IN2(data_in[7]), .S(n58), .Q(n805) );
  MUX21X1 U245 ( .IN1(\fifo[10][6] ), .IN2(data_in[6]), .S(n58), .Q(n804) );
  MUX21X1 U246 ( .IN1(\fifo[10][5] ), .IN2(data_in[5]), .S(n58), .Q(n803) );
  MUX21X1 U247 ( .IN1(\fifo[10][4] ), .IN2(data_in[4]), .S(n58), .Q(n802) );
  MUX21X1 U248 ( .IN1(\fifo[10][3] ), .IN2(data_in[3]), .S(n58), .Q(n801) );
  MUX21X1 U249 ( .IN1(\fifo[10][2] ), .IN2(data_in[2]), .S(n58), .Q(n800) );
  MUX21X1 U250 ( .IN1(\fifo[10][1] ), .IN2(data_in[1]), .S(n58), .Q(n799) );
  MUX21X1 U251 ( .IN1(\fifo[10][0] ), .IN2(data_in[0]), .S(n58), .Q(n798) );
  AND2X1 U252 ( .IN1(n55), .IN2(n52), .Q(n58) );
  MUX21X1 U253 ( .IN1(\fifo[11][31] ), .IN2(data_in[31]), .S(n59), .Q(n797) );
  MUX21X1 U254 ( .IN1(\fifo[11][30] ), .IN2(data_in[30]), .S(n59), .Q(n796) );
  MUX21X1 U255 ( .IN1(\fifo[11][29] ), .IN2(data_in[29]), .S(n59), .Q(n795) );
  MUX21X1 U256 ( .IN1(\fifo[11][28] ), .IN2(data_in[28]), .S(n59), .Q(n794) );
  MUX21X1 U257 ( .IN1(\fifo[11][27] ), .IN2(data_in[27]), .S(n59), .Q(n793) );
  MUX21X1 U258 ( .IN1(\fifo[11][26] ), .IN2(data_in[26]), .S(n59), .Q(n792) );
  MUX21X1 U259 ( .IN1(\fifo[11][25] ), .IN2(data_in[25]), .S(n59), .Q(n791) );
  MUX21X1 U260 ( .IN1(\fifo[11][24] ), .IN2(data_in[24]), .S(n59), .Q(n790) );
  MUX21X1 U261 ( .IN1(\fifo[11][23] ), .IN2(data_in[23]), .S(n59), .Q(n789) );
  MUX21X1 U262 ( .IN1(\fifo[11][22] ), .IN2(data_in[22]), .S(n59), .Q(n788) );
  MUX21X1 U263 ( .IN1(\fifo[11][21] ), .IN2(data_in[21]), .S(n59), .Q(n787) );
  MUX21X1 U264 ( .IN1(\fifo[11][20] ), .IN2(data_in[20]), .S(n59), .Q(n786) );
  MUX21X1 U265 ( .IN1(\fifo[11][19] ), .IN2(data_in[19]), .S(n59), .Q(n785) );
  MUX21X1 U266 ( .IN1(\fifo[11][18] ), .IN2(data_in[18]), .S(n59), .Q(n784) );
  MUX21X1 U267 ( .IN1(\fifo[11][17] ), .IN2(data_in[17]), .S(n59), .Q(n783) );
  MUX21X1 U268 ( .IN1(\fifo[11][16] ), .IN2(data_in[16]), .S(n59), .Q(n782) );
  MUX21X1 U269 ( .IN1(\fifo[11][15] ), .IN2(data_in[15]), .S(n59), .Q(n781) );
  MUX21X1 U270 ( .IN1(\fifo[11][14] ), .IN2(data_in[14]), .S(n59), .Q(n780) );
  MUX21X1 U271 ( .IN1(\fifo[11][13] ), .IN2(data_in[13]), .S(n59), .Q(n779) );
  MUX21X1 U272 ( .IN1(\fifo[11][12] ), .IN2(data_in[12]), .S(n59), .Q(n778) );
  MUX21X1 U273 ( .IN1(\fifo[11][11] ), .IN2(data_in[11]), .S(n59), .Q(n777) );
  MUX21X1 U274 ( .IN1(\fifo[11][10] ), .IN2(data_in[10]), .S(n59), .Q(n776) );
  MUX21X1 U275 ( .IN1(\fifo[11][9] ), .IN2(data_in[9]), .S(n59), .Q(n775) );
  MUX21X1 U276 ( .IN1(\fifo[11][8] ), .IN2(data_in[8]), .S(n59), .Q(n774) );
  MUX21X1 U277 ( .IN1(\fifo[11][7] ), .IN2(data_in[7]), .S(n59), .Q(n773) );
  MUX21X1 U278 ( .IN1(\fifo[11][6] ), .IN2(data_in[6]), .S(n59), .Q(n772) );
  MUX21X1 U279 ( .IN1(\fifo[11][5] ), .IN2(data_in[5]), .S(n59), .Q(n771) );
  MUX21X1 U280 ( .IN1(\fifo[11][4] ), .IN2(data_in[4]), .S(n59), .Q(n770) );
  MUX21X1 U281 ( .IN1(\fifo[11][3] ), .IN2(data_in[3]), .S(n59), .Q(n769) );
  MUX21X1 U282 ( .IN1(\fifo[11][2] ), .IN2(data_in[2]), .S(n59), .Q(n768) );
  MUX21X1 U283 ( .IN1(\fifo[11][1] ), .IN2(data_in[1]), .S(n59), .Q(n767) );
  MUX21X1 U284 ( .IN1(\fifo[11][0] ), .IN2(data_in[0]), .S(n59), .Q(n766) );
  AND2X1 U285 ( .IN1(n55), .IN2(n60), .Q(n59) );
  MUX21X1 U286 ( .IN1(\fifo[12][31] ), .IN2(data_in[31]), .S(n61), .Q(n765) );
  MUX21X1 U287 ( .IN1(\fifo[12][30] ), .IN2(data_in[30]), .S(n61), .Q(n764) );
  MUX21X1 U288 ( .IN1(\fifo[12][29] ), .IN2(data_in[29]), .S(n61), .Q(n763) );
  MUX21X1 U289 ( .IN1(\fifo[12][28] ), .IN2(data_in[28]), .S(n61), .Q(n762) );
  MUX21X1 U290 ( .IN1(\fifo[12][27] ), .IN2(data_in[27]), .S(n61), .Q(n761) );
  MUX21X1 U291 ( .IN1(\fifo[12][26] ), .IN2(data_in[26]), .S(n61), .Q(n760) );
  MUX21X1 U292 ( .IN1(\fifo[12][25] ), .IN2(data_in[25]), .S(n61), .Q(n759) );
  MUX21X1 U293 ( .IN1(\fifo[12][24] ), .IN2(data_in[24]), .S(n61), .Q(n758) );
  MUX21X1 U294 ( .IN1(\fifo[12][23] ), .IN2(data_in[23]), .S(n61), .Q(n757) );
  MUX21X1 U295 ( .IN1(\fifo[12][22] ), .IN2(data_in[22]), .S(n61), .Q(n756) );
  MUX21X1 U296 ( .IN1(\fifo[12][21] ), .IN2(data_in[21]), .S(n61), .Q(n755) );
  MUX21X1 U297 ( .IN1(\fifo[12][20] ), .IN2(data_in[20]), .S(n61), .Q(n754) );
  MUX21X1 U298 ( .IN1(\fifo[12][19] ), .IN2(data_in[19]), .S(n61), .Q(n753) );
  MUX21X1 U299 ( .IN1(\fifo[12][18] ), .IN2(data_in[18]), .S(n61), .Q(n752) );
  MUX21X1 U300 ( .IN1(\fifo[12][17] ), .IN2(data_in[17]), .S(n61), .Q(n751) );
  MUX21X1 U301 ( .IN1(\fifo[12][16] ), .IN2(data_in[16]), .S(n61), .Q(n750) );
  MUX21X1 U302 ( .IN1(\fifo[12][15] ), .IN2(data_in[15]), .S(n61), .Q(n749) );
  MUX21X1 U303 ( .IN1(\fifo[12][14] ), .IN2(data_in[14]), .S(n61), .Q(n748) );
  MUX21X1 U304 ( .IN1(\fifo[12][13] ), .IN2(data_in[13]), .S(n61), .Q(n747) );
  MUX21X1 U305 ( .IN1(\fifo[12][12] ), .IN2(data_in[12]), .S(n61), .Q(n746) );
  MUX21X1 U306 ( .IN1(\fifo[12][11] ), .IN2(data_in[11]), .S(n61), .Q(n745) );
  MUX21X1 U307 ( .IN1(\fifo[12][10] ), .IN2(data_in[10]), .S(n61), .Q(n744) );
  MUX21X1 U308 ( .IN1(\fifo[12][9] ), .IN2(data_in[9]), .S(n61), .Q(n743) );
  MUX21X1 U309 ( .IN1(\fifo[12][8] ), .IN2(data_in[8]), .S(n61), .Q(n742) );
  MUX21X1 U310 ( .IN1(\fifo[12][7] ), .IN2(data_in[7]), .S(n61), .Q(n741) );
  MUX21X1 U311 ( .IN1(\fifo[12][6] ), .IN2(data_in[6]), .S(n61), .Q(n740) );
  MUX21X1 U312 ( .IN1(\fifo[12][5] ), .IN2(data_in[5]), .S(n61), .Q(n739) );
  MUX21X1 U313 ( .IN1(\fifo[12][4] ), .IN2(data_in[4]), .S(n61), .Q(n738) );
  MUX21X1 U314 ( .IN1(\fifo[12][3] ), .IN2(data_in[3]), .S(n61), .Q(n737) );
  MUX21X1 U315 ( .IN1(\fifo[12][2] ), .IN2(data_in[2]), .S(n61), .Q(n736) );
  MUX21X1 U316 ( .IN1(\fifo[12][1] ), .IN2(data_in[1]), .S(n61), .Q(n735) );
  MUX21X1 U317 ( .IN1(\fifo[12][0] ), .IN2(data_in[0]), .S(n61), .Q(n734) );
  AND2X1 U318 ( .IN1(n62), .IN2(n56), .Q(n61) );
  MUX21X1 U319 ( .IN1(\fifo[13][31] ), .IN2(data_in[31]), .S(n63), .Q(n733) );
  MUX21X1 U320 ( .IN1(\fifo[13][30] ), .IN2(data_in[30]), .S(n63), .Q(n732) );
  MUX21X1 U321 ( .IN1(\fifo[13][29] ), .IN2(data_in[29]), .S(n63), .Q(n731) );
  MUX21X1 U322 ( .IN1(\fifo[13][28] ), .IN2(data_in[28]), .S(n63), .Q(n730) );
  MUX21X1 U323 ( .IN1(\fifo[13][27] ), .IN2(data_in[27]), .S(n63), .Q(n729) );
  MUX21X1 U324 ( .IN1(\fifo[13][26] ), .IN2(data_in[26]), .S(n63), .Q(n728) );
  MUX21X1 U325 ( .IN1(\fifo[13][25] ), .IN2(data_in[25]), .S(n63), .Q(n727) );
  MUX21X1 U326 ( .IN1(\fifo[13][24] ), .IN2(data_in[24]), .S(n63), .Q(n726) );
  MUX21X1 U327 ( .IN1(\fifo[13][23] ), .IN2(data_in[23]), .S(n63), .Q(n725) );
  MUX21X1 U328 ( .IN1(\fifo[13][22] ), .IN2(data_in[22]), .S(n63), .Q(n724) );
  MUX21X1 U329 ( .IN1(\fifo[13][21] ), .IN2(data_in[21]), .S(n63), .Q(n723) );
  MUX21X1 U330 ( .IN1(\fifo[13][20] ), .IN2(data_in[20]), .S(n63), .Q(n722) );
  MUX21X1 U331 ( .IN1(\fifo[13][19] ), .IN2(data_in[19]), .S(n63), .Q(n721) );
  MUX21X1 U332 ( .IN1(\fifo[13][18] ), .IN2(data_in[18]), .S(n63), .Q(n720) );
  MUX21X1 U333 ( .IN1(\fifo[13][17] ), .IN2(data_in[17]), .S(n63), .Q(n719) );
  MUX21X1 U334 ( .IN1(\fifo[13][16] ), .IN2(data_in[16]), .S(n63), .Q(n718) );
  MUX21X1 U335 ( .IN1(\fifo[13][15] ), .IN2(data_in[15]), .S(n63), .Q(n717) );
  MUX21X1 U336 ( .IN1(\fifo[13][14] ), .IN2(data_in[14]), .S(n63), .Q(n716) );
  MUX21X1 U337 ( .IN1(\fifo[13][13] ), .IN2(data_in[13]), .S(n63), .Q(n715) );
  MUX21X1 U338 ( .IN1(\fifo[13][12] ), .IN2(data_in[12]), .S(n63), .Q(n714) );
  MUX21X1 U339 ( .IN1(\fifo[13][11] ), .IN2(data_in[11]), .S(n63), .Q(n713) );
  MUX21X1 U340 ( .IN1(\fifo[13][10] ), .IN2(data_in[10]), .S(n63), .Q(n712) );
  MUX21X1 U341 ( .IN1(\fifo[13][9] ), .IN2(data_in[9]), .S(n63), .Q(n711) );
  MUX21X1 U342 ( .IN1(\fifo[13][8] ), .IN2(data_in[8]), .S(n63), .Q(n710) );
  MUX21X1 U343 ( .IN1(\fifo[13][7] ), .IN2(data_in[7]), .S(n63), .Q(n709) );
  MUX21X1 U344 ( .IN1(\fifo[13][6] ), .IN2(data_in[6]), .S(n63), .Q(n708) );
  MUX21X1 U345 ( .IN1(\fifo[13][5] ), .IN2(data_in[5]), .S(n63), .Q(n707) );
  MUX21X1 U346 ( .IN1(\fifo[13][4] ), .IN2(data_in[4]), .S(n63), .Q(n706) );
  MUX21X1 U347 ( .IN1(\fifo[13][3] ), .IN2(data_in[3]), .S(n63), .Q(n705) );
  MUX21X1 U348 ( .IN1(\fifo[13][2] ), .IN2(data_in[2]), .S(n63), .Q(n704) );
  MUX21X1 U349 ( .IN1(\fifo[13][1] ), .IN2(data_in[1]), .S(n63), .Q(n703) );
  MUX21X1 U350 ( .IN1(\fifo[13][0] ), .IN2(data_in[0]), .S(n63), .Q(n702) );
  AND2X1 U351 ( .IN1(n62), .IN2(n49), .Q(n63) );
  MUX21X1 U352 ( .IN1(\fifo[14][31] ), .IN2(data_in[31]), .S(n64), .Q(n701) );
  MUX21X1 U353 ( .IN1(\fifo[14][30] ), .IN2(data_in[30]), .S(n64), .Q(n700) );
  MUX21X1 U354 ( .IN1(\fifo[14][29] ), .IN2(data_in[29]), .S(n64), .Q(n699) );
  MUX21X1 U355 ( .IN1(\fifo[14][28] ), .IN2(data_in[28]), .S(n64), .Q(n698) );
  MUX21X1 U356 ( .IN1(\fifo[14][27] ), .IN2(data_in[27]), .S(n64), .Q(n697) );
  MUX21X1 U357 ( .IN1(\fifo[14][26] ), .IN2(data_in[26]), .S(n64), .Q(n696) );
  MUX21X1 U358 ( .IN1(\fifo[14][25] ), .IN2(data_in[25]), .S(n64), .Q(n695) );
  MUX21X1 U359 ( .IN1(\fifo[14][24] ), .IN2(data_in[24]), .S(n64), .Q(n694) );
  MUX21X1 U360 ( .IN1(\fifo[14][23] ), .IN2(data_in[23]), .S(n64), .Q(n693) );
  MUX21X1 U361 ( .IN1(\fifo[14][22] ), .IN2(data_in[22]), .S(n64), .Q(n692) );
  MUX21X1 U362 ( .IN1(\fifo[14][21] ), .IN2(data_in[21]), .S(n64), .Q(n691) );
  MUX21X1 U363 ( .IN1(\fifo[14][20] ), .IN2(data_in[20]), .S(n64), .Q(n690) );
  MUX21X1 U364 ( .IN1(\fifo[14][19] ), .IN2(data_in[19]), .S(n64), .Q(n689) );
  MUX21X1 U365 ( .IN1(\fifo[14][18] ), .IN2(data_in[18]), .S(n64), .Q(n688) );
  MUX21X1 U366 ( .IN1(\fifo[14][17] ), .IN2(data_in[17]), .S(n64), .Q(n687) );
  MUX21X1 U367 ( .IN1(\fifo[14][16] ), .IN2(data_in[16]), .S(n64), .Q(n686) );
  MUX21X1 U368 ( .IN1(\fifo[14][15] ), .IN2(data_in[15]), .S(n64), .Q(n685) );
  MUX21X1 U369 ( .IN1(\fifo[14][14] ), .IN2(data_in[14]), .S(n64), .Q(n684) );
  MUX21X1 U370 ( .IN1(\fifo[14][13] ), .IN2(data_in[13]), .S(n64), .Q(n683) );
  MUX21X1 U371 ( .IN1(\fifo[14][12] ), .IN2(data_in[12]), .S(n64), .Q(n682) );
  MUX21X1 U372 ( .IN1(\fifo[14][11] ), .IN2(data_in[11]), .S(n64), .Q(n681) );
  MUX21X1 U373 ( .IN1(\fifo[14][10] ), .IN2(data_in[10]), .S(n64), .Q(n680) );
  MUX21X1 U374 ( .IN1(\fifo[14][9] ), .IN2(data_in[9]), .S(n64), .Q(n679) );
  MUX21X1 U375 ( .IN1(\fifo[14][8] ), .IN2(data_in[8]), .S(n64), .Q(n678) );
  MUX21X1 U376 ( .IN1(\fifo[14][7] ), .IN2(data_in[7]), .S(n64), .Q(n677) );
  MUX21X1 U377 ( .IN1(\fifo[14][6] ), .IN2(data_in[6]), .S(n64), .Q(n676) );
  MUX21X1 U378 ( .IN1(\fifo[14][5] ), .IN2(data_in[5]), .S(n64), .Q(n675) );
  MUX21X1 U379 ( .IN1(\fifo[14][4] ), .IN2(data_in[4]), .S(n64), .Q(n674) );
  MUX21X1 U380 ( .IN1(\fifo[14][3] ), .IN2(data_in[3]), .S(n64), .Q(n673) );
  MUX21X1 U381 ( .IN1(\fifo[14][2] ), .IN2(data_in[2]), .S(n64), .Q(n672) );
  MUX21X1 U382 ( .IN1(\fifo[14][1] ), .IN2(data_in[1]), .S(n64), .Q(n671) );
  MUX21X1 U383 ( .IN1(\fifo[14][0] ), .IN2(data_in[0]), .S(n64), .Q(n670) );
  AND2X1 U384 ( .IN1(n62), .IN2(n52), .Q(n64) );
  MUX21X1 U385 ( .IN1(\fifo[15][31] ), .IN2(data_in[31]), .S(n65), .Q(n669) );
  MUX21X1 U386 ( .IN1(\fifo[15][30] ), .IN2(data_in[30]), .S(n65), .Q(n668) );
  MUX21X1 U387 ( .IN1(\fifo[15][29] ), .IN2(data_in[29]), .S(n65), .Q(n667) );
  MUX21X1 U388 ( .IN1(\fifo[15][28] ), .IN2(data_in[28]), .S(n65), .Q(n666) );
  MUX21X1 U389 ( .IN1(\fifo[15][27] ), .IN2(data_in[27]), .S(n65), .Q(n665) );
  MUX21X1 U390 ( .IN1(\fifo[15][26] ), .IN2(data_in[26]), .S(n65), .Q(n664) );
  MUX21X1 U391 ( .IN1(\fifo[15][25] ), .IN2(data_in[25]), .S(n65), .Q(n663) );
  MUX21X1 U392 ( .IN1(\fifo[15][24] ), .IN2(data_in[24]), .S(n65), .Q(n662) );
  MUX21X1 U393 ( .IN1(\fifo[15][23] ), .IN2(data_in[23]), .S(n65), .Q(n661) );
  MUX21X1 U394 ( .IN1(\fifo[15][22] ), .IN2(data_in[22]), .S(n65), .Q(n660) );
  MUX21X1 U395 ( .IN1(\fifo[15][21] ), .IN2(data_in[21]), .S(n65), .Q(n659) );
  MUX21X1 U396 ( .IN1(\fifo[15][20] ), .IN2(data_in[20]), .S(n65), .Q(n658) );
  MUX21X1 U397 ( .IN1(\fifo[15][19] ), .IN2(data_in[19]), .S(n65), .Q(n657) );
  MUX21X1 U398 ( .IN1(\fifo[15][18] ), .IN2(data_in[18]), .S(n65), .Q(n656) );
  MUX21X1 U399 ( .IN1(\fifo[15][17] ), .IN2(data_in[17]), .S(n65), .Q(n655) );
  MUX21X1 U400 ( .IN1(\fifo[15][16] ), .IN2(data_in[16]), .S(n65), .Q(n654) );
  MUX21X1 U401 ( .IN1(\fifo[15][15] ), .IN2(data_in[15]), .S(n65), .Q(n653) );
  MUX21X1 U402 ( .IN1(\fifo[15][14] ), .IN2(data_in[14]), .S(n65), .Q(n652) );
  MUX21X1 U403 ( .IN1(\fifo[15][13] ), .IN2(data_in[13]), .S(n65), .Q(n651) );
  MUX21X1 U404 ( .IN1(\fifo[15][12] ), .IN2(data_in[12]), .S(n65), .Q(n650) );
  MUX21X1 U405 ( .IN1(\fifo[15][11] ), .IN2(data_in[11]), .S(n65), .Q(n649) );
  MUX21X1 U406 ( .IN1(\fifo[15][10] ), .IN2(data_in[10]), .S(n65), .Q(n648) );
  MUX21X1 U407 ( .IN1(\fifo[15][9] ), .IN2(data_in[9]), .S(n65), .Q(n647) );
  MUX21X1 U408 ( .IN1(\fifo[15][8] ), .IN2(data_in[8]), .S(n65), .Q(n646) );
  MUX21X1 U409 ( .IN1(\fifo[15][7] ), .IN2(data_in[7]), .S(n65), .Q(n645) );
  MUX21X1 U410 ( .IN1(\fifo[15][6] ), .IN2(data_in[6]), .S(n65), .Q(n644) );
  MUX21X1 U411 ( .IN1(\fifo[15][5] ), .IN2(data_in[5]), .S(n65), .Q(n643) );
  MUX21X1 U412 ( .IN1(\fifo[15][4] ), .IN2(data_in[4]), .S(n65), .Q(n642) );
  MUX21X1 U413 ( .IN1(\fifo[15][3] ), .IN2(data_in[3]), .S(n65), .Q(n641) );
  MUX21X1 U414 ( .IN1(\fifo[15][2] ), .IN2(data_in[2]), .S(n65), .Q(n640) );
  MUX21X1 U415 ( .IN1(\fifo[15][1] ), .IN2(data_in[1]), .S(n65), .Q(n639) );
  MUX21X1 U416 ( .IN1(\fifo[15][0] ), .IN2(data_in[0]), .S(n65), .Q(n638) );
  AND2X1 U417 ( .IN1(n62), .IN2(n60), .Q(n65) );
  NOR2X0 U418 ( .IN1(n3), .IN2(n1), .QN(n62) );
  AO21X1 U419 ( .IN1(clear), .IN2(n66), .IN3(n67), .Q(n1162) );
  MUX21X1 U420 ( .IN1(n68), .IN2(n69), .S(n1311), .Q(n67) );
  AO22X1 U421 ( .IN1(n68), .IN2(cnt[1]), .IN3(n69), .IN4(n70), .Q(n1161) );
  AO21X1 U422 ( .IN1(n71), .IN2(\U3/U1/Z_0 ), .IN3(n72), .Q(n70) );
  MUX21X1 U423 ( .IN1(n73), .IN2(n74), .S(n584), .Q(n72) );
  XOR2X1 U424 ( .IN1(cnt[0]), .IN2(\U3/U1/Z_0 ), .Q(n74) );
  NOR2X0 U425 ( .IN1(\U3/U1/Z_0 ), .IN2(cnt[0]), .QN(n73) );
  AO22X1 U426 ( .IN1(n68), .IN2(cnt[2]), .IN3(n69), .IN4(n75), .Q(n1160) );
  XOR3X1 U427 ( .IN1(\U3/U1/Z_0 ), .IN2(cnt[2]), .IN3(n76), .Q(n75) );
  AO22X1 U428 ( .IN1(n68), .IN2(cnt[3]), .IN3(n69), .IN4(n77), .Q(n1159) );
  XOR3X1 U429 ( .IN1(n1313), .IN2(\U3/U1/Z_0 ), .IN3(n78), .Q(n77) );
  AO22X1 U430 ( .IN1(n68), .IN2(cnt[4]), .IN3(n69), .IN4(n79), .Q(n1158) );
  XOR3X1 U431 ( .IN1(n564), .IN2(\U3/U1/Z_0 ), .IN3(n80), .Q(n79) );
  OA22X1 U432 ( .IN1(n1313), .IN2(n81), .IN3(n78), .IN4(n82), .Q(n80) );
  INVX0 U433 ( .INP(n83), .ZN(n78) );
  NOR2X0 U434 ( .IN1(\U3/U1/Z_0 ), .IN2(n83), .QN(n81) );
  AO22X1 U435 ( .IN1(\U3/U1/Z_0 ), .IN2(n76), .IN3(n84), .IN4(cnt[2]), .Q(n83)
         );
  OR2X1 U436 ( .IN1(n76), .IN2(\U3/U1/Z_0 ), .Q(n84) );
  AO21X1 U437 ( .IN1(\U3/U1/Z_0 ), .IN2(n85), .IN3(n71), .Q(n76) );
  NAND2X0 U438 ( .IN1(n1311), .IN2(n584), .QN(n85) );
  NOR2X0 U439 ( .IN1(n69), .IN2(clear), .QN(n68) );
  AND2X1 U440 ( .IN1(n66), .IN2(n86), .Q(n69) );
  XNOR2X1 U441 ( .IN1(write), .IN2(n82), .Q(n66) );
  INVX0 U442 ( .INP(\U3/U1/Z_0 ), .ZN(n82) );
  AO21X1 U443 ( .IN1(clear), .IN2(\U3/U1/Z_0 ), .IN3(n87), .Q(n1157) );
  MUX21X1 U444 ( .IN1(n88), .IN2(n89), .S(n588), .Q(n87) );
  AO22X1 U445 ( .IN1(n88), .IN2(N15), .IN3(n89), .IN4(n90), .Q(n1156) );
  OR2X1 U446 ( .IN1(n91), .IN2(n92), .Q(n90) );
  MUX21X1 U447 ( .IN1(n93), .IN2(n94), .S(n586), .Q(n1155) );
  NOR2X0 U448 ( .IN1(n95), .IN2(n96), .QN(n94) );
  AO22X1 U449 ( .IN1(n93), .IN2(N17), .IN3(n89), .IN4(n97), .Q(n1154) );
  NAND2X0 U450 ( .IN1(n98), .IN2(n99), .QN(n97) );
  AO21X1 U451 ( .IN1(n89), .IN2(n96), .IN3(n88), .Q(n93) );
  NOR2X0 U452 ( .IN1(n89), .IN2(clear), .QN(n88) );
  INVX0 U453 ( .INP(n95), .ZN(n89) );
  NAND3X0 U454 ( .IN1(n45), .IN2(n86), .IN3(\U3/U1/Z_0 ), .QN(n95) );
  NAND3X0 U455 ( .IN1(n1311), .IN2(n100), .IN3(n564), .QN(n45) );
  AO221X1 U456 ( .IN1(n101), .IN2(write_pointer[0]), .IN3(clear), .IN4(write), 
        .IN5(n102), .Q(n1153) );
  NAND3X0 U457 ( .IN1(n103), .IN2(n104), .IN3(n105), .QN(n1152) );
  NAND2X0 U458 ( .IN1(n101), .IN2(write_pointer[1]), .QN(n105) );
  INVX0 U459 ( .INP(n106), .ZN(n101) );
  MUX21X1 U460 ( .IN1(n60), .IN2(n107), .S(write_pointer[2]), .Q(n1151) );
  AO221X1 U461 ( .IN1(write_pointer[3]), .IN2(n107), .IN3(n55), .IN4(n108), 
        .IN5(n53), .Q(n1150) );
  AND2X1 U462 ( .IN1(n60), .IN2(n50), .Q(n53) );
  NOR2X0 U463 ( .IN1(n3), .IN2(write_pointer[2]), .QN(n55) );
  NAND3X0 U464 ( .IN1(n106), .IN2(n109), .IN3(n110), .QN(n107) );
  NAND2X0 U465 ( .IN1(n108), .IN2(n4), .QN(n110) );
  NAND2X0 U466 ( .IN1(n111), .IN2(n86), .QN(n106) );
  MUX21X1 U467 ( .IN1(data_in[31]), .IN2(\fifo[0][31] ), .S(n112), .Q(n1149)
         );
  MUX21X1 U468 ( .IN1(data_in[30]), .IN2(\fifo[0][30] ), .S(n112), .Q(n1148)
         );
  MUX21X1 U469 ( .IN1(data_in[29]), .IN2(\fifo[0][29] ), .S(n112), .Q(n1147)
         );
  MUX21X1 U470 ( .IN1(data_in[28]), .IN2(\fifo[0][28] ), .S(n112), .Q(n1146)
         );
  MUX21X1 U471 ( .IN1(data_in[27]), .IN2(\fifo[0][27] ), .S(n112), .Q(n1145)
         );
  MUX21X1 U472 ( .IN1(data_in[26]), .IN2(\fifo[0][26] ), .S(n112), .Q(n1144)
         );
  MUX21X1 U473 ( .IN1(data_in[25]), .IN2(\fifo[0][25] ), .S(n112), .Q(n1143)
         );
  MUX21X1 U474 ( .IN1(data_in[24]), .IN2(\fifo[0][24] ), .S(n112), .Q(n1142)
         );
  MUX21X1 U475 ( .IN1(data_in[23]), .IN2(\fifo[0][23] ), .S(n112), .Q(n1141)
         );
  MUX21X1 U476 ( .IN1(data_in[22]), .IN2(\fifo[0][22] ), .S(n112), .Q(n1140)
         );
  MUX21X1 U477 ( .IN1(data_in[21]), .IN2(\fifo[0][21] ), .S(n112), .Q(n1139)
         );
  MUX21X1 U478 ( .IN1(data_in[20]), .IN2(\fifo[0][20] ), .S(n112), .Q(n1138)
         );
  MUX21X1 U479 ( .IN1(data_in[19]), .IN2(\fifo[0][19] ), .S(n112), .Q(n1137)
         );
  MUX21X1 U480 ( .IN1(data_in[18]), .IN2(\fifo[0][18] ), .S(n112), .Q(n1136)
         );
  MUX21X1 U481 ( .IN1(data_in[17]), .IN2(\fifo[0][17] ), .S(n112), .Q(n1135)
         );
  MUX21X1 U482 ( .IN1(data_in[16]), .IN2(\fifo[0][16] ), .S(n112), .Q(n1134)
         );
  MUX21X1 U483 ( .IN1(data_in[15]), .IN2(\fifo[0][15] ), .S(n112), .Q(n1133)
         );
  MUX21X1 U484 ( .IN1(data_in[14]), .IN2(\fifo[0][14] ), .S(n112), .Q(n1132)
         );
  MUX21X1 U485 ( .IN1(data_in[13]), .IN2(\fifo[0][13] ), .S(n112), .Q(n1131)
         );
  MUX21X1 U486 ( .IN1(data_in[12]), .IN2(\fifo[0][12] ), .S(n112), .Q(n1130)
         );
  MUX21X1 U487 ( .IN1(data_in[11]), .IN2(\fifo[0][11] ), .S(n112), .Q(n1129)
         );
  MUX21X1 U488 ( .IN1(data_in[10]), .IN2(\fifo[0][10] ), .S(n112), .Q(n1128)
         );
  MUX21X1 U489 ( .IN1(data_in[9]), .IN2(\fifo[0][9] ), .S(n112), .Q(n1127) );
  MUX21X1 U490 ( .IN1(data_in[8]), .IN2(\fifo[0][8] ), .S(n112), .Q(n1126) );
  MUX21X1 U491 ( .IN1(data_in[7]), .IN2(\fifo[0][7] ), .S(n112), .Q(n1125) );
  MUX21X1 U492 ( .IN1(data_in[6]), .IN2(\fifo[0][6] ), .S(n112), .Q(n1124) );
  MUX21X1 U493 ( .IN1(data_in[5]), .IN2(\fifo[0][5] ), .S(n112), .Q(n1123) );
  MUX21X1 U494 ( .IN1(data_in[4]), .IN2(\fifo[0][4] ), .S(n112), .Q(n1122) );
  MUX21X1 U495 ( .IN1(data_in[3]), .IN2(\fifo[0][3] ), .S(n112), .Q(n1121) );
  MUX21X1 U496 ( .IN1(data_in[2]), .IN2(\fifo[0][2] ), .S(n112), .Q(n1120) );
  MUX21X1 U497 ( .IN1(data_in[1]), .IN2(\fifo[0][1] ), .S(n112), .Q(n1119) );
  MUX21X1 U498 ( .IN1(data_in[0]), .IN2(\fifo[0][0] ), .S(n112), .Q(n1118) );
  AOI22X1 U499 ( .IN1(clear), .IN2(write), .IN3(n113), .IN4(n56), .QN(n112) );
  MUX21X1 U500 ( .IN1(\fifo[1][31] ), .IN2(data_in[31]), .S(n114), .Q(n1117)
         );
  MUX21X1 U501 ( .IN1(\fifo[1][30] ), .IN2(data_in[30]), .S(n114), .Q(n1116)
         );
  MUX21X1 U502 ( .IN1(\fifo[1][29] ), .IN2(data_in[29]), .S(n114), .Q(n1115)
         );
  MUX21X1 U503 ( .IN1(\fifo[1][28] ), .IN2(data_in[28]), .S(n114), .Q(n1114)
         );
  MUX21X1 U504 ( .IN1(\fifo[1][27] ), .IN2(data_in[27]), .S(n114), .Q(n1113)
         );
  MUX21X1 U505 ( .IN1(\fifo[1][26] ), .IN2(data_in[26]), .S(n114), .Q(n1112)
         );
  MUX21X1 U506 ( .IN1(\fifo[1][25] ), .IN2(data_in[25]), .S(n114), .Q(n1111)
         );
  MUX21X1 U507 ( .IN1(\fifo[1][24] ), .IN2(data_in[24]), .S(n114), .Q(n1110)
         );
  MUX21X1 U508 ( .IN1(\fifo[1][23] ), .IN2(data_in[23]), .S(n114), .Q(n1109)
         );
  MUX21X1 U509 ( .IN1(\fifo[1][22] ), .IN2(data_in[22]), .S(n114), .Q(n1108)
         );
  MUX21X1 U510 ( .IN1(\fifo[1][21] ), .IN2(data_in[21]), .S(n114), .Q(n1107)
         );
  MUX21X1 U511 ( .IN1(\fifo[1][20] ), .IN2(data_in[20]), .S(n114), .Q(n1106)
         );
  MUX21X1 U512 ( .IN1(\fifo[1][19] ), .IN2(data_in[19]), .S(n114), .Q(n1105)
         );
  MUX21X1 U513 ( .IN1(\fifo[1][18] ), .IN2(data_in[18]), .S(n114), .Q(n1104)
         );
  MUX21X1 U514 ( .IN1(\fifo[1][17] ), .IN2(data_in[17]), .S(n114), .Q(n1103)
         );
  MUX21X1 U515 ( .IN1(\fifo[1][16] ), .IN2(data_in[16]), .S(n114), .Q(n1102)
         );
  MUX21X1 U516 ( .IN1(\fifo[1][15] ), .IN2(data_in[15]), .S(n114), .Q(n1101)
         );
  MUX21X1 U517 ( .IN1(\fifo[1][14] ), .IN2(data_in[14]), .S(n114), .Q(n1100)
         );
  MUX21X1 U518 ( .IN1(\fifo[1][13] ), .IN2(data_in[13]), .S(n114), .Q(n1099)
         );
  MUX21X1 U519 ( .IN1(\fifo[1][12] ), .IN2(data_in[12]), .S(n114), .Q(n1098)
         );
  MUX21X1 U520 ( .IN1(\fifo[1][11] ), .IN2(data_in[11]), .S(n114), .Q(n1097)
         );
  MUX21X1 U521 ( .IN1(\fifo[1][10] ), .IN2(data_in[10]), .S(n114), .Q(n1096)
         );
  MUX21X1 U522 ( .IN1(\fifo[1][9] ), .IN2(data_in[9]), .S(n114), .Q(n1095) );
  MUX21X1 U523 ( .IN1(\fifo[1][8] ), .IN2(data_in[8]), .S(n114), .Q(n1094) );
  MUX21X1 U524 ( .IN1(\fifo[1][7] ), .IN2(data_in[7]), .S(n114), .Q(n1093) );
  MUX21X1 U525 ( .IN1(\fifo[1][6] ), .IN2(data_in[6]), .S(n114), .Q(n1092) );
  MUX21X1 U526 ( .IN1(\fifo[1][5] ), .IN2(data_in[5]), .S(n114), .Q(n1091) );
  MUX21X1 U527 ( .IN1(\fifo[1][4] ), .IN2(data_in[4]), .S(n114), .Q(n1090) );
  MUX21X1 U528 ( .IN1(\fifo[1][3] ), .IN2(data_in[3]), .S(n114), .Q(n1089) );
  MUX21X1 U529 ( .IN1(\fifo[1][2] ), .IN2(data_in[2]), .S(n114), .Q(n1088) );
  MUX21X1 U530 ( .IN1(\fifo[1][1] ), .IN2(data_in[1]), .S(n114), .Q(n1087) );
  MUX21X1 U531 ( .IN1(\fifo[1][0] ), .IN2(data_in[0]), .S(n114), .Q(n1086) );
  AND2X1 U532 ( .IN1(n113), .IN2(n49), .Q(n114) );
  INVX0 U533 ( .INP(n103), .ZN(n49) );
  NAND3X0 U534 ( .IN1(n108), .IN2(n4), .IN3(write_pointer[0]), .QN(n103) );
  MUX21X1 U535 ( .IN1(\fifo[2][31] ), .IN2(data_in[31]), .S(n115), .Q(n1085)
         );
  MUX21X1 U536 ( .IN1(\fifo[2][30] ), .IN2(data_in[30]), .S(n115), .Q(n1084)
         );
  MUX21X1 U537 ( .IN1(\fifo[2][29] ), .IN2(data_in[29]), .S(n115), .Q(n1083)
         );
  MUX21X1 U538 ( .IN1(\fifo[2][28] ), .IN2(data_in[28]), .S(n115), .Q(n1082)
         );
  MUX21X1 U539 ( .IN1(\fifo[2][27] ), .IN2(data_in[27]), .S(n115), .Q(n1081)
         );
  MUX21X1 U540 ( .IN1(\fifo[2][26] ), .IN2(data_in[26]), .S(n115), .Q(n1080)
         );
  MUX21X1 U541 ( .IN1(\fifo[2][25] ), .IN2(data_in[25]), .S(n115), .Q(n1079)
         );
  MUX21X1 U542 ( .IN1(\fifo[2][24] ), .IN2(data_in[24]), .S(n115), .Q(n1078)
         );
  MUX21X1 U543 ( .IN1(\fifo[2][23] ), .IN2(data_in[23]), .S(n115), .Q(n1077)
         );
  MUX21X1 U544 ( .IN1(\fifo[2][22] ), .IN2(data_in[22]), .S(n115), .Q(n1076)
         );
  MUX21X1 U545 ( .IN1(\fifo[2][21] ), .IN2(data_in[21]), .S(n115), .Q(n1075)
         );
  MUX21X1 U546 ( .IN1(\fifo[2][20] ), .IN2(data_in[20]), .S(n115), .Q(n1074)
         );
  MUX21X1 U547 ( .IN1(\fifo[2][19] ), .IN2(data_in[19]), .S(n115), .Q(n1073)
         );
  MUX21X1 U548 ( .IN1(\fifo[2][18] ), .IN2(data_in[18]), .S(n115), .Q(n1072)
         );
  MUX21X1 U549 ( .IN1(\fifo[2][17] ), .IN2(data_in[17]), .S(n115), .Q(n1071)
         );
  MUX21X1 U550 ( .IN1(\fifo[2][16] ), .IN2(data_in[16]), .S(n115), .Q(n1070)
         );
  MUX21X1 U551 ( .IN1(\fifo[2][15] ), .IN2(data_in[15]), .S(n115), .Q(n1069)
         );
  MUX21X1 U552 ( .IN1(\fifo[2][14] ), .IN2(data_in[14]), .S(n115), .Q(n1068)
         );
  MUX21X1 U553 ( .IN1(\fifo[2][13] ), .IN2(data_in[13]), .S(n115), .Q(n1067)
         );
  MUX21X1 U554 ( .IN1(\fifo[2][12] ), .IN2(data_in[12]), .S(n115), .Q(n1066)
         );
  MUX21X1 U555 ( .IN1(\fifo[2][11] ), .IN2(data_in[11]), .S(n115), .Q(n1065)
         );
  MUX21X1 U556 ( .IN1(\fifo[2][10] ), .IN2(data_in[10]), .S(n115), .Q(n1064)
         );
  MUX21X1 U557 ( .IN1(\fifo[2][9] ), .IN2(data_in[9]), .S(n115), .Q(n1063) );
  MUX21X1 U558 ( .IN1(\fifo[2][8] ), .IN2(data_in[8]), .S(n115), .Q(n1062) );
  MUX21X1 U559 ( .IN1(\fifo[2][7] ), .IN2(data_in[7]), .S(n115), .Q(n1061) );
  MUX21X1 U560 ( .IN1(\fifo[2][6] ), .IN2(data_in[6]), .S(n115), .Q(n1060) );
  MUX21X1 U561 ( .IN1(\fifo[2][5] ), .IN2(data_in[5]), .S(n115), .Q(n1059) );
  MUX21X1 U562 ( .IN1(\fifo[2][4] ), .IN2(data_in[4]), .S(n115), .Q(n1058) );
  MUX21X1 U563 ( .IN1(\fifo[2][3] ), .IN2(data_in[3]), .S(n115), .Q(n1057) );
  MUX21X1 U564 ( .IN1(\fifo[2][2] ), .IN2(data_in[2]), .S(n115), .Q(n1056) );
  MUX21X1 U565 ( .IN1(\fifo[2][1] ), .IN2(data_in[1]), .S(n115), .Q(n1055) );
  MUX21X1 U566 ( .IN1(\fifo[2][0] ), .IN2(data_in[0]), .S(n115), .Q(n1054) );
  AND2X1 U567 ( .IN1(n113), .IN2(n52), .Q(n115) );
  INVX0 U568 ( .INP(n104), .ZN(n52) );
  NAND2X0 U569 ( .IN1(write_pointer[1]), .IN2(n102), .QN(n104) );
  MUX21X1 U570 ( .IN1(\fifo[3][31] ), .IN2(data_in[31]), .S(n116), .Q(n1053)
         );
  MUX21X1 U571 ( .IN1(\fifo[3][30] ), .IN2(data_in[30]), .S(n116), .Q(n1052)
         );
  MUX21X1 U572 ( .IN1(\fifo[3][29] ), .IN2(data_in[29]), .S(n116), .Q(n1051)
         );
  MUX21X1 U573 ( .IN1(\fifo[3][28] ), .IN2(data_in[28]), .S(n116), .Q(n1050)
         );
  MUX21X1 U574 ( .IN1(\fifo[3][27] ), .IN2(data_in[27]), .S(n116), .Q(n1049)
         );
  MUX21X1 U575 ( .IN1(\fifo[3][26] ), .IN2(data_in[26]), .S(n116), .Q(n1048)
         );
  MUX21X1 U576 ( .IN1(\fifo[3][25] ), .IN2(data_in[25]), .S(n116), .Q(n1047)
         );
  MUX21X1 U577 ( .IN1(\fifo[3][24] ), .IN2(data_in[24]), .S(n116), .Q(n1046)
         );
  MUX21X1 U578 ( .IN1(\fifo[3][23] ), .IN2(data_in[23]), .S(n116), .Q(n1045)
         );
  MUX21X1 U579 ( .IN1(\fifo[3][22] ), .IN2(data_in[22]), .S(n116), .Q(n1044)
         );
  MUX21X1 U580 ( .IN1(\fifo[3][21] ), .IN2(data_in[21]), .S(n116), .Q(n1043)
         );
  MUX21X1 U581 ( .IN1(\fifo[3][20] ), .IN2(data_in[20]), .S(n116), .Q(n1042)
         );
  MUX21X1 U582 ( .IN1(\fifo[3][19] ), .IN2(data_in[19]), .S(n116), .Q(n1041)
         );
  MUX21X1 U583 ( .IN1(\fifo[3][18] ), .IN2(data_in[18]), .S(n116), .Q(n1040)
         );
  MUX21X1 U584 ( .IN1(\fifo[3][17] ), .IN2(data_in[17]), .S(n116), .Q(n1039)
         );
  MUX21X1 U585 ( .IN1(\fifo[3][16] ), .IN2(data_in[16]), .S(n116), .Q(n1038)
         );
  MUX21X1 U586 ( .IN1(\fifo[3][15] ), .IN2(data_in[15]), .S(n116), .Q(n1037)
         );
  MUX21X1 U587 ( .IN1(\fifo[3][14] ), .IN2(data_in[14]), .S(n116), .Q(n1036)
         );
  MUX21X1 U588 ( .IN1(\fifo[3][13] ), .IN2(data_in[13]), .S(n116), .Q(n1035)
         );
  MUX21X1 U589 ( .IN1(\fifo[3][12] ), .IN2(data_in[12]), .S(n116), .Q(n1034)
         );
  MUX21X1 U590 ( .IN1(\fifo[3][11] ), .IN2(data_in[11]), .S(n116), .Q(n1033)
         );
  MUX21X1 U591 ( .IN1(\fifo[3][10] ), .IN2(data_in[10]), .S(n116), .Q(n1032)
         );
  MUX21X1 U592 ( .IN1(\fifo[3][9] ), .IN2(data_in[9]), .S(n116), .Q(n1031) );
  MUX21X1 U593 ( .IN1(\fifo[3][8] ), .IN2(data_in[8]), .S(n116), .Q(n1030) );
  MUX21X1 U594 ( .IN1(\fifo[3][7] ), .IN2(data_in[7]), .S(n116), .Q(n1029) );
  MUX21X1 U595 ( .IN1(\fifo[3][6] ), .IN2(data_in[6]), .S(n116), .Q(n1028) );
  MUX21X1 U596 ( .IN1(\fifo[3][5] ), .IN2(data_in[5]), .S(n116), .Q(n1027) );
  MUX21X1 U597 ( .IN1(\fifo[3][4] ), .IN2(data_in[4]), .S(n116), .Q(n1026) );
  MUX21X1 U598 ( .IN1(\fifo[3][3] ), .IN2(data_in[3]), .S(n116), .Q(n1025) );
  MUX21X1 U599 ( .IN1(\fifo[3][2] ), .IN2(data_in[2]), .S(n116), .Q(n1024) );
  MUX21X1 U600 ( .IN1(\fifo[3][1] ), .IN2(data_in[1]), .S(n116), .Q(n1023) );
  MUX21X1 U601 ( .IN1(\fifo[3][0] ), .IN2(data_in[0]), .S(n116), .Q(n1022) );
  AND2X1 U602 ( .IN1(n113), .IN2(n60), .Q(n116) );
  AND3X1 U603 ( .IN1(write_pointer[0]), .IN2(n108), .IN3(write_pointer[1]), 
        .Q(n60) );
  INVX0 U604 ( .INP(n111), .ZN(n108) );
  NOR2X0 U605 ( .IN1(write_pointer[3]), .IN2(write_pointer[2]), .QN(n113) );
  MUX21X1 U606 ( .IN1(\fifo[4][31] ), .IN2(data_in[31]), .S(n47), .Q(n1021) );
  MUX21X1 U607 ( .IN1(\fifo[4][30] ), .IN2(data_in[30]), .S(n47), .Q(n1020) );
  MUX21X1 U608 ( .IN1(\fifo[4][29] ), .IN2(data_in[29]), .S(n47), .Q(n1019) );
  MUX21X1 U609 ( .IN1(\fifo[4][28] ), .IN2(data_in[28]), .S(n47), .Q(n1018) );
  MUX21X1 U610 ( .IN1(\fifo[4][27] ), .IN2(data_in[27]), .S(n47), .Q(n1017) );
  MUX21X1 U611 ( .IN1(\fifo[4][26] ), .IN2(data_in[26]), .S(n47), .Q(n1016) );
  MUX21X1 U612 ( .IN1(\fifo[4][25] ), .IN2(data_in[25]), .S(n47), .Q(n1015) );
  MUX21X1 U613 ( .IN1(\fifo[4][24] ), .IN2(data_in[24]), .S(n47), .Q(n1014) );
  MUX21X1 U614 ( .IN1(\fifo[4][23] ), .IN2(data_in[23]), .S(n47), .Q(n1013) );
  MUX21X1 U615 ( .IN1(\fifo[4][22] ), .IN2(data_in[22]), .S(n47), .Q(n1012) );
  MUX21X1 U616 ( .IN1(\fifo[4][21] ), .IN2(data_in[21]), .S(n47), .Q(n1011) );
  MUX21X1 U617 ( .IN1(\fifo[4][20] ), .IN2(data_in[20]), .S(n47), .Q(n1010) );
  MUX21X1 U618 ( .IN1(\fifo[4][19] ), .IN2(data_in[19]), .S(n47), .Q(n1009) );
  MUX21X1 U619 ( .IN1(\fifo[4][18] ), .IN2(data_in[18]), .S(n47), .Q(n1008) );
  MUX21X1 U620 ( .IN1(\fifo[4][17] ), .IN2(data_in[17]), .S(n47), .Q(n1007) );
  MUX21X1 U621 ( .IN1(\fifo[4][16] ), .IN2(data_in[16]), .S(n47), .Q(n1006) );
  MUX21X1 U622 ( .IN1(\fifo[4][15] ), .IN2(data_in[15]), .S(n47), .Q(n1005) );
  MUX21X1 U623 ( .IN1(\fifo[4][14] ), .IN2(data_in[14]), .S(n47), .Q(n1004) );
  MUX21X1 U624 ( .IN1(\fifo[4][13] ), .IN2(data_in[13]), .S(n47), .Q(n1003) );
  MUX21X1 U625 ( .IN1(\fifo[4][12] ), .IN2(data_in[12]), .S(n47), .Q(n1002) );
  MUX21X1 U626 ( .IN1(\fifo[4][11] ), .IN2(data_in[11]), .S(n47), .Q(n1001) );
  MUX21X1 U627 ( .IN1(\fifo[4][10] ), .IN2(data_in[10]), .S(n47), .Q(n1000) );
  AND2X1 U628 ( .IN1(n56), .IN2(n50), .Q(n47) );
  NOR2X0 U629 ( .IN1(n1), .IN2(write_pointer[3]), .QN(n50) );
  NOR2X0 U630 ( .IN1(n109), .IN2(write_pointer[1]), .QN(n56) );
  INVX0 U631 ( .INP(n102), .ZN(n109) );
  NOR2X0 U632 ( .IN1(n111), .IN2(write_pointer[0]), .QN(n102) );
  NAND3X0 U633 ( .IN1(n46), .IN2(n86), .IN3(write), .QN(n111) );
  INVX0 U634 ( .INP(clear), .ZN(n86) );
  NAND3X0 U635 ( .IN1(n100), .IN2(cnt[4]), .IN3(n1311), .QN(n46) );
  AND3X1 U636 ( .IN1(cnt[2]), .IN2(cnt[3]), .IN3(n71), .Q(almost_full) );
  NOR2X0 U637 ( .IN1(n1311), .IN2(n584), .QN(n71) );
  AND3X1 U638 ( .IN1(n564), .IN2(cnt[0]), .IN3(n100), .Q(almost_empty) );
  AND3X1 U639 ( .IN1(n1313), .IN2(n1312), .IN3(n584), .Q(n100) );
  MUX21X1 U640 ( .IN1(n117), .IN2(\fifo[0][31] ), .S(clear), .Q(N155) );
  NAND4X0 U641 ( .IN1(n118), .IN2(n119), .IN3(n120), .IN4(n121), .QN(n117) );
  OA221X1 U642 ( .IN1(n1917), .IN2(n122), .IN3(n1565), .IN4(n123), .IN5(n124), 
        .Q(n121) );
  OA22X1 U643 ( .IN1(n1693), .IN2(n125), .IN3(n1939), .IN4(n126), .Q(n124) );
  OA221X1 U644 ( .IN1(n1597), .IN2(n127), .IN3(n1469), .IN4(n128), .IN5(n129), 
        .Q(n120) );
  OA22X1 U645 ( .IN1(n1821), .IN2(n130), .IN3(n1725), .IN4(n131), .Q(n129) );
  OA221X1 U646 ( .IN1(n1629), .IN2(n132), .IN3(n1501), .IN4(n133), .IN5(n134), 
        .Q(n119) );
  OA22X1 U647 ( .IN1(n1853), .IN2(n135), .IN3(n1757), .IN4(n136), .Q(n134) );
  OA221X1 U648 ( .IN1(n1789), .IN2(n137), .IN3(n1885), .IN4(n138), .IN5(n139), 
        .Q(n118) );
  OA22X1 U649 ( .IN1(n1661), .IN2(n140), .IN3(n1533), .IN4(n98), .Q(n139) );
  MUX21X1 U650 ( .IN1(n141), .IN2(\fifo[0][30] ), .S(clear), .Q(N154) );
  NAND4X0 U651 ( .IN1(n142), .IN2(n143), .IN3(n144), .IN4(n145), .QN(n141) );
  OA221X1 U652 ( .IN1(n1918), .IN2(n122), .IN3(n1566), .IN4(n123), .IN5(n146), 
        .Q(n145) );
  OA22X1 U653 ( .IN1(n1694), .IN2(n125), .IN3(n1940), .IN4(n126), .Q(n146) );
  OA221X1 U654 ( .IN1(n1598), .IN2(n127), .IN3(n1470), .IN4(n128), .IN5(n147), 
        .Q(n144) );
  OA22X1 U655 ( .IN1(n1822), .IN2(n130), .IN3(n1726), .IN4(n131), .Q(n147) );
  OA221X1 U656 ( .IN1(n1630), .IN2(n132), .IN3(n1502), .IN4(n133), .IN5(n148), 
        .Q(n143) );
  OA22X1 U657 ( .IN1(n1854), .IN2(n135), .IN3(n1758), .IN4(n136), .Q(n148) );
  OA221X1 U658 ( .IN1(n1790), .IN2(n137), .IN3(n1886), .IN4(n138), .IN5(n149), 
        .Q(n142) );
  OA22X1 U659 ( .IN1(n1662), .IN2(n140), .IN3(n1534), .IN4(n98), .Q(n149) );
  MUX21X1 U660 ( .IN1(n150), .IN2(\fifo[0][29] ), .S(clear), .Q(N153) );
  NAND4X0 U661 ( .IN1(n151), .IN2(n152), .IN3(n153), .IN4(n154), .QN(n150) );
  OA221X1 U662 ( .IN1(n1919), .IN2(n122), .IN3(n1567), .IN4(n123), .IN5(n155), 
        .Q(n154) );
  OA22X1 U663 ( .IN1(n1695), .IN2(n125), .IN3(n1941), .IN4(n126), .Q(n155) );
  OA221X1 U664 ( .IN1(n1599), .IN2(n127), .IN3(n1471), .IN4(n128), .IN5(n156), 
        .Q(n153) );
  OA22X1 U665 ( .IN1(n1823), .IN2(n130), .IN3(n1727), .IN4(n131), .Q(n156) );
  OA221X1 U666 ( .IN1(n1631), .IN2(n132), .IN3(n1503), .IN4(n133), .IN5(n157), 
        .Q(n152) );
  OA22X1 U667 ( .IN1(n1855), .IN2(n135), .IN3(n1759), .IN4(n136), .Q(n157) );
  OA221X1 U668 ( .IN1(n1791), .IN2(n137), .IN3(n1887), .IN4(n138), .IN5(n158), 
        .Q(n151) );
  OA22X1 U669 ( .IN1(n1663), .IN2(n140), .IN3(n1535), .IN4(n98), .Q(n158) );
  MUX21X1 U670 ( .IN1(n159), .IN2(\fifo[0][28] ), .S(clear), .Q(N152) );
  NAND4X0 U671 ( .IN1(n160), .IN2(n161), .IN3(n162), .IN4(n163), .QN(n159) );
  OA221X1 U672 ( .IN1(n1920), .IN2(n122), .IN3(n1568), .IN4(n123), .IN5(n164), 
        .Q(n163) );
  OA22X1 U673 ( .IN1(n1696), .IN2(n125), .IN3(n1942), .IN4(n126), .Q(n164) );
  OA221X1 U674 ( .IN1(n1600), .IN2(n127), .IN3(n1472), .IN4(n128), .IN5(n165), 
        .Q(n162) );
  OA22X1 U675 ( .IN1(n1824), .IN2(n130), .IN3(n1728), .IN4(n131), .Q(n165) );
  OA221X1 U676 ( .IN1(n1632), .IN2(n132), .IN3(n1504), .IN4(n133), .IN5(n166), 
        .Q(n161) );
  OA22X1 U677 ( .IN1(n1856), .IN2(n135), .IN3(n1760), .IN4(n136), .Q(n166) );
  OA221X1 U678 ( .IN1(n1792), .IN2(n137), .IN3(n1888), .IN4(n138), .IN5(n167), 
        .Q(n160) );
  OA22X1 U679 ( .IN1(n1664), .IN2(n140), .IN3(n1536), .IN4(n98), .Q(n167) );
  MUX21X1 U680 ( .IN1(n168), .IN2(\fifo[0][27] ), .S(clear), .Q(N151) );
  NAND4X0 U681 ( .IN1(n169), .IN2(n170), .IN3(n171), .IN4(n172), .QN(n168) );
  OA221X1 U682 ( .IN1(n1921), .IN2(n122), .IN3(n1569), .IN4(n123), .IN5(n173), 
        .Q(n172) );
  OA22X1 U683 ( .IN1(n1697), .IN2(n125), .IN3(n1943), .IN4(n126), .Q(n173) );
  OA221X1 U684 ( .IN1(n1601), .IN2(n127), .IN3(n1473), .IN4(n128), .IN5(n174), 
        .Q(n171) );
  OA22X1 U685 ( .IN1(n1825), .IN2(n130), .IN3(n1729), .IN4(n131), .Q(n174) );
  OA221X1 U686 ( .IN1(n1633), .IN2(n132), .IN3(n1505), .IN4(n133), .IN5(n175), 
        .Q(n170) );
  OA22X1 U687 ( .IN1(n1857), .IN2(n135), .IN3(n1761), .IN4(n136), .Q(n175) );
  OA221X1 U688 ( .IN1(n1793), .IN2(n137), .IN3(n1889), .IN4(n138), .IN5(n176), 
        .Q(n169) );
  OA22X1 U689 ( .IN1(n1665), .IN2(n140), .IN3(n1537), .IN4(n98), .Q(n176) );
  MUX21X1 U690 ( .IN1(n177), .IN2(\fifo[0][26] ), .S(clear), .Q(N150) );
  NAND4X0 U691 ( .IN1(n178), .IN2(n179), .IN3(n180), .IN4(n181), .QN(n177) );
  OA221X1 U692 ( .IN1(n1922), .IN2(n122), .IN3(n1570), .IN4(n123), .IN5(n182), 
        .Q(n181) );
  OA22X1 U693 ( .IN1(n1698), .IN2(n125), .IN3(n1944), .IN4(n126), .Q(n182) );
  OA221X1 U694 ( .IN1(n1602), .IN2(n127), .IN3(n1474), .IN4(n128), .IN5(n183), 
        .Q(n180) );
  OA22X1 U695 ( .IN1(n1826), .IN2(n130), .IN3(n1730), .IN4(n131), .Q(n183) );
  OA221X1 U696 ( .IN1(n1634), .IN2(n132), .IN3(n1506), .IN4(n133), .IN5(n184), 
        .Q(n179) );
  OA22X1 U697 ( .IN1(n1858), .IN2(n135), .IN3(n1762), .IN4(n136), .Q(n184) );
  OA221X1 U698 ( .IN1(n1794), .IN2(n137), .IN3(n1890), .IN4(n138), .IN5(n185), 
        .Q(n178) );
  OA22X1 U699 ( .IN1(n1666), .IN2(n140), .IN3(n1538), .IN4(n98), .Q(n185) );
  MUX21X1 U700 ( .IN1(n186), .IN2(\fifo[0][25] ), .S(clear), .Q(N149) );
  NAND4X0 U701 ( .IN1(n187), .IN2(n188), .IN3(n189), .IN4(n190), .QN(n186) );
  OA221X1 U702 ( .IN1(n1923), .IN2(n122), .IN3(n1571), .IN4(n123), .IN5(n191), 
        .Q(n190) );
  OA22X1 U703 ( .IN1(n1699), .IN2(n125), .IN3(n1945), .IN4(n126), .Q(n191) );
  OA221X1 U704 ( .IN1(n1603), .IN2(n127), .IN3(n1475), .IN4(n128), .IN5(n192), 
        .Q(n189) );
  OA22X1 U705 ( .IN1(n1827), .IN2(n130), .IN3(n1731), .IN4(n131), .Q(n192) );
  OA221X1 U706 ( .IN1(n1635), .IN2(n132), .IN3(n1507), .IN4(n133), .IN5(n193), 
        .Q(n188) );
  OA22X1 U707 ( .IN1(n1859), .IN2(n135), .IN3(n1763), .IN4(n136), .Q(n193) );
  OA221X1 U708 ( .IN1(n1795), .IN2(n137), .IN3(n1891), .IN4(n138), .IN5(n194), 
        .Q(n187) );
  OA22X1 U709 ( .IN1(n1667), .IN2(n140), .IN3(n1539), .IN4(n98), .Q(n194) );
  MUX21X1 U710 ( .IN1(n195), .IN2(\fifo[0][24] ), .S(clear), .Q(N148) );
  NAND4X0 U711 ( .IN1(n196), .IN2(n197), .IN3(n198), .IN4(n199), .QN(n195) );
  OA221X1 U712 ( .IN1(n1924), .IN2(n122), .IN3(n1572), .IN4(n123), .IN5(n200), 
        .Q(n199) );
  OA22X1 U713 ( .IN1(n1700), .IN2(n125), .IN3(n1946), .IN4(n126), .Q(n200) );
  OA221X1 U714 ( .IN1(n1604), .IN2(n127), .IN3(n1476), .IN4(n128), .IN5(n201), 
        .Q(n198) );
  OA22X1 U715 ( .IN1(n1828), .IN2(n130), .IN3(n1732), .IN4(n131), .Q(n201) );
  OA221X1 U716 ( .IN1(n1636), .IN2(n132), .IN3(n1508), .IN4(n133), .IN5(n202), 
        .Q(n197) );
  OA22X1 U717 ( .IN1(n1860), .IN2(n135), .IN3(n1764), .IN4(n136), .Q(n202) );
  OA221X1 U718 ( .IN1(n1796), .IN2(n137), .IN3(n1892), .IN4(n138), .IN5(n203), 
        .Q(n196) );
  OA22X1 U719 ( .IN1(n1668), .IN2(n140), .IN3(n1540), .IN4(n98), .Q(n203) );
  MUX21X1 U720 ( .IN1(n204), .IN2(\fifo[0][23] ), .S(clear), .Q(N147) );
  NAND4X0 U721 ( .IN1(n205), .IN2(n206), .IN3(n207), .IN4(n208), .QN(n204) );
  OA221X1 U722 ( .IN1(n1925), .IN2(n122), .IN3(n1573), .IN4(n123), .IN5(n209), 
        .Q(n208) );
  OA22X1 U723 ( .IN1(n1701), .IN2(n125), .IN3(n1947), .IN4(n126), .Q(n209) );
  OA221X1 U724 ( .IN1(n1605), .IN2(n127), .IN3(n1477), .IN4(n128), .IN5(n210), 
        .Q(n207) );
  OA22X1 U725 ( .IN1(n1829), .IN2(n130), .IN3(n1733), .IN4(n131), .Q(n210) );
  OA221X1 U726 ( .IN1(n1637), .IN2(n132), .IN3(n1509), .IN4(n133), .IN5(n211), 
        .Q(n206) );
  OA22X1 U727 ( .IN1(n1861), .IN2(n135), .IN3(n1765), .IN4(n136), .Q(n211) );
  OA221X1 U728 ( .IN1(n1797), .IN2(n137), .IN3(n1893), .IN4(n138), .IN5(n212), 
        .Q(n205) );
  OA22X1 U729 ( .IN1(n1669), .IN2(n140), .IN3(n1541), .IN4(n98), .Q(n212) );
  MUX21X1 U730 ( .IN1(n213), .IN2(\fifo[0][22] ), .S(clear), .Q(N146) );
  NAND4X0 U731 ( .IN1(n214), .IN2(n215), .IN3(n216), .IN4(n217), .QN(n213) );
  OA221X1 U732 ( .IN1(n1926), .IN2(n122), .IN3(n1574), .IN4(n123), .IN5(n218), 
        .Q(n217) );
  OA22X1 U733 ( .IN1(n1702), .IN2(n125), .IN3(n1948), .IN4(n126), .Q(n218) );
  OA221X1 U734 ( .IN1(n1606), .IN2(n127), .IN3(n1478), .IN4(n128), .IN5(n219), 
        .Q(n216) );
  OA22X1 U735 ( .IN1(n1830), .IN2(n130), .IN3(n1734), .IN4(n131), .Q(n219) );
  OA221X1 U736 ( .IN1(n1638), .IN2(n132), .IN3(n1510), .IN4(n133), .IN5(n220), 
        .Q(n215) );
  OA22X1 U737 ( .IN1(n1862), .IN2(n135), .IN3(n1766), .IN4(n136), .Q(n220) );
  OA221X1 U738 ( .IN1(n1798), .IN2(n137), .IN3(n1894), .IN4(n138), .IN5(n221), 
        .Q(n214) );
  OA22X1 U739 ( .IN1(n1670), .IN2(n140), .IN3(n1542), .IN4(n98), .Q(n221) );
  MUX21X1 U740 ( .IN1(n222), .IN2(\fifo[0][21] ), .S(clear), .Q(N145) );
  NAND4X0 U741 ( .IN1(n223), .IN2(n224), .IN3(n225), .IN4(n226), .QN(n222) );
  OA221X1 U742 ( .IN1(n1927), .IN2(n122), .IN3(n1575), .IN4(n123), .IN5(n227), 
        .Q(n226) );
  OA22X1 U743 ( .IN1(n1703), .IN2(n125), .IN3(n1949), .IN4(n126), .Q(n227) );
  OA221X1 U744 ( .IN1(n1607), .IN2(n127), .IN3(n1479), .IN4(n128), .IN5(n228), 
        .Q(n225) );
  OA22X1 U745 ( .IN1(n1831), .IN2(n130), .IN3(n1735), .IN4(n131), .Q(n228) );
  OA221X1 U746 ( .IN1(n1639), .IN2(n132), .IN3(n1511), .IN4(n133), .IN5(n229), 
        .Q(n224) );
  OA22X1 U747 ( .IN1(n1863), .IN2(n135), .IN3(n1767), .IN4(n136), .Q(n229) );
  OA221X1 U748 ( .IN1(n1799), .IN2(n137), .IN3(n1895), .IN4(n138), .IN5(n230), 
        .Q(n223) );
  OA22X1 U749 ( .IN1(n1671), .IN2(n140), .IN3(n1543), .IN4(n98), .Q(n230) );
  MUX21X1 U750 ( .IN1(n231), .IN2(\fifo[0][20] ), .S(clear), .Q(N144) );
  NAND4X0 U751 ( .IN1(n232), .IN2(n233), .IN3(n234), .IN4(n235), .QN(n231) );
  OA221X1 U752 ( .IN1(n1928), .IN2(n122), .IN3(n1576), .IN4(n123), .IN5(n236), 
        .Q(n235) );
  OA22X1 U753 ( .IN1(n1704), .IN2(n125), .IN3(n1950), .IN4(n126), .Q(n236) );
  OA221X1 U754 ( .IN1(n1608), .IN2(n127), .IN3(n1480), .IN4(n128), .IN5(n237), 
        .Q(n234) );
  OA22X1 U755 ( .IN1(n1832), .IN2(n130), .IN3(n1736), .IN4(n131), .Q(n237) );
  OA221X1 U756 ( .IN1(n1640), .IN2(n132), .IN3(n1512), .IN4(n133), .IN5(n238), 
        .Q(n233) );
  OA22X1 U757 ( .IN1(n1864), .IN2(n135), .IN3(n1768), .IN4(n136), .Q(n238) );
  OA221X1 U758 ( .IN1(n1800), .IN2(n137), .IN3(n1896), .IN4(n138), .IN5(n239), 
        .Q(n232) );
  OA22X1 U759 ( .IN1(n1672), .IN2(n140), .IN3(n1544), .IN4(n98), .Q(n239) );
  MUX21X1 U760 ( .IN1(n240), .IN2(\fifo[0][19] ), .S(clear), .Q(N143) );
  NAND4X0 U761 ( .IN1(n241), .IN2(n242), .IN3(n243), .IN4(n244), .QN(n240) );
  OA221X1 U762 ( .IN1(n1929), .IN2(n122), .IN3(n1577), .IN4(n123), .IN5(n245), 
        .Q(n244) );
  OA22X1 U763 ( .IN1(n1705), .IN2(n125), .IN3(n1951), .IN4(n126), .Q(n245) );
  OA221X1 U764 ( .IN1(n1609), .IN2(n127), .IN3(n1481), .IN4(n128), .IN5(n246), 
        .Q(n243) );
  OA22X1 U765 ( .IN1(n1833), .IN2(n130), .IN3(n1737), .IN4(n131), .Q(n246) );
  OA221X1 U766 ( .IN1(n1641), .IN2(n132), .IN3(n1513), .IN4(n133), .IN5(n247), 
        .Q(n242) );
  OA22X1 U767 ( .IN1(n1865), .IN2(n135), .IN3(n1769), .IN4(n136), .Q(n247) );
  OA221X1 U768 ( .IN1(n1801), .IN2(n137), .IN3(n1897), .IN4(n138), .IN5(n248), 
        .Q(n241) );
  OA22X1 U769 ( .IN1(n1673), .IN2(n140), .IN3(n1545), .IN4(n98), .Q(n248) );
  MUX21X1 U770 ( .IN1(n249), .IN2(\fifo[0][18] ), .S(clear), .Q(N142) );
  NAND4X0 U771 ( .IN1(n250), .IN2(n251), .IN3(n252), .IN4(n253), .QN(n249) );
  OA221X1 U772 ( .IN1(n1930), .IN2(n122), .IN3(n1578), .IN4(n123), .IN5(n254), 
        .Q(n253) );
  OA22X1 U773 ( .IN1(n1706), .IN2(n125), .IN3(n1952), .IN4(n126), .Q(n254) );
  OA221X1 U774 ( .IN1(n1610), .IN2(n127), .IN3(n1482), .IN4(n128), .IN5(n255), 
        .Q(n252) );
  OA22X1 U775 ( .IN1(n1834), .IN2(n130), .IN3(n1738), .IN4(n131), .Q(n255) );
  OA221X1 U776 ( .IN1(n1642), .IN2(n132), .IN3(n1514), .IN4(n133), .IN5(n256), 
        .Q(n251) );
  OA22X1 U777 ( .IN1(n1866), .IN2(n135), .IN3(n1770), .IN4(n136), .Q(n256) );
  OA221X1 U778 ( .IN1(n1802), .IN2(n137), .IN3(n1898), .IN4(n138), .IN5(n257), 
        .Q(n250) );
  OA22X1 U779 ( .IN1(n1674), .IN2(n140), .IN3(n1546), .IN4(n98), .Q(n257) );
  MUX21X1 U780 ( .IN1(n258), .IN2(\fifo[0][17] ), .S(clear), .Q(N141) );
  NAND4X0 U781 ( .IN1(n259), .IN2(n260), .IN3(n261), .IN4(n262), .QN(n258) );
  OA221X1 U782 ( .IN1(n1931), .IN2(n122), .IN3(n1579), .IN4(n123), .IN5(n263), 
        .Q(n262) );
  OA22X1 U783 ( .IN1(n1707), .IN2(n125), .IN3(n1953), .IN4(n126), .Q(n263) );
  OA221X1 U784 ( .IN1(n1611), .IN2(n127), .IN3(n1483), .IN4(n128), .IN5(n264), 
        .Q(n261) );
  OA22X1 U785 ( .IN1(n1835), .IN2(n130), .IN3(n1739), .IN4(n131), .Q(n264) );
  OA221X1 U786 ( .IN1(n1643), .IN2(n132), .IN3(n1515), .IN4(n133), .IN5(n265), 
        .Q(n260) );
  OA22X1 U787 ( .IN1(n1867), .IN2(n135), .IN3(n1771), .IN4(n136), .Q(n265) );
  OA221X1 U788 ( .IN1(n1803), .IN2(n137), .IN3(n1899), .IN4(n138), .IN5(n266), 
        .Q(n259) );
  OA22X1 U789 ( .IN1(n1675), .IN2(n140), .IN3(n1547), .IN4(n98), .Q(n266) );
  MUX21X1 U790 ( .IN1(n267), .IN2(\fifo[0][16] ), .S(clear), .Q(N140) );
  NAND4X0 U791 ( .IN1(n268), .IN2(n269), .IN3(n270), .IN4(n271), .QN(n267) );
  OA221X1 U792 ( .IN1(n1932), .IN2(n122), .IN3(n1580), .IN4(n123), .IN5(n272), 
        .Q(n271) );
  OA22X1 U793 ( .IN1(n1708), .IN2(n125), .IN3(n1954), .IN4(n126), .Q(n272) );
  OA221X1 U794 ( .IN1(n1612), .IN2(n127), .IN3(n1484), .IN4(n128), .IN5(n273), 
        .Q(n270) );
  OA22X1 U795 ( .IN1(n1836), .IN2(n130), .IN3(n1740), .IN4(n131), .Q(n273) );
  OA221X1 U796 ( .IN1(n1644), .IN2(n132), .IN3(n1516), .IN4(n133), .IN5(n274), 
        .Q(n269) );
  OA22X1 U797 ( .IN1(n1868), .IN2(n135), .IN3(n1772), .IN4(n136), .Q(n274) );
  OA221X1 U798 ( .IN1(n1804), .IN2(n137), .IN3(n1900), .IN4(n138), .IN5(n275), 
        .Q(n268) );
  OA22X1 U799 ( .IN1(n1676), .IN2(n140), .IN3(n1548), .IN4(n98), .Q(n275) );
  MUX21X1 U800 ( .IN1(n276), .IN2(\fifo[0][15] ), .S(clear), .Q(N139) );
  NAND4X0 U801 ( .IN1(n277), .IN2(n278), .IN3(n279), .IN4(n280), .QN(n276) );
  OA221X1 U802 ( .IN1(n1933), .IN2(n122), .IN3(n1581), .IN4(n123), .IN5(n281), 
        .Q(n280) );
  OA22X1 U803 ( .IN1(n1709), .IN2(n125), .IN3(n1955), .IN4(n126), .Q(n281) );
  OA221X1 U804 ( .IN1(n1613), .IN2(n127), .IN3(n1485), .IN4(n128), .IN5(n282), 
        .Q(n279) );
  OA22X1 U805 ( .IN1(n1837), .IN2(n130), .IN3(n1741), .IN4(n131), .Q(n282) );
  OA221X1 U806 ( .IN1(n1645), .IN2(n132), .IN3(n1517), .IN4(n133), .IN5(n283), 
        .Q(n278) );
  OA22X1 U807 ( .IN1(n1869), .IN2(n135), .IN3(n1773), .IN4(n136), .Q(n283) );
  OA221X1 U808 ( .IN1(n1805), .IN2(n137), .IN3(n1901), .IN4(n138), .IN5(n284), 
        .Q(n277) );
  OA22X1 U809 ( .IN1(n1677), .IN2(n140), .IN3(n1549), .IN4(n98), .Q(n284) );
  MUX21X1 U810 ( .IN1(n285), .IN2(\fifo[0][14] ), .S(clear), .Q(N138) );
  NAND4X0 U811 ( .IN1(n286), .IN2(n287), .IN3(n288), .IN4(n289), .QN(n285) );
  OA221X1 U812 ( .IN1(n1934), .IN2(n122), .IN3(n1582), .IN4(n123), .IN5(n290), 
        .Q(n289) );
  OA22X1 U813 ( .IN1(n1710), .IN2(n125), .IN3(n1956), .IN4(n126), .Q(n290) );
  OA221X1 U814 ( .IN1(n1614), .IN2(n127), .IN3(n1486), .IN4(n128), .IN5(n291), 
        .Q(n288) );
  OA22X1 U815 ( .IN1(n1838), .IN2(n130), .IN3(n1742), .IN4(n131), .Q(n291) );
  OA221X1 U816 ( .IN1(n1646), .IN2(n132), .IN3(n1518), .IN4(n133), .IN5(n292), 
        .Q(n287) );
  OA22X1 U817 ( .IN1(n1870), .IN2(n135), .IN3(n1774), .IN4(n136), .Q(n292) );
  OA221X1 U818 ( .IN1(n1806), .IN2(n137), .IN3(n1902), .IN4(n138), .IN5(n293), 
        .Q(n286) );
  OA22X1 U819 ( .IN1(n1678), .IN2(n140), .IN3(n1550), .IN4(n98), .Q(n293) );
  MUX21X1 U820 ( .IN1(n294), .IN2(\fifo[0][13] ), .S(clear), .Q(N137) );
  NAND4X0 U821 ( .IN1(n295), .IN2(n296), .IN3(n297), .IN4(n298), .QN(n294) );
  OA221X1 U822 ( .IN1(n1935), .IN2(n122), .IN3(n1583), .IN4(n123), .IN5(n299), 
        .Q(n298) );
  OA22X1 U823 ( .IN1(n1711), .IN2(n125), .IN3(n1957), .IN4(n126), .Q(n299) );
  OA221X1 U824 ( .IN1(n1615), .IN2(n127), .IN3(n1487), .IN4(n128), .IN5(n300), 
        .Q(n297) );
  OA22X1 U825 ( .IN1(n1839), .IN2(n130), .IN3(n1743), .IN4(n131), .Q(n300) );
  OA221X1 U826 ( .IN1(n1647), .IN2(n132), .IN3(n1519), .IN4(n133), .IN5(n301), 
        .Q(n296) );
  OA22X1 U827 ( .IN1(n1871), .IN2(n135), .IN3(n1775), .IN4(n136), .Q(n301) );
  OA221X1 U828 ( .IN1(n1807), .IN2(n137), .IN3(n1903), .IN4(n138), .IN5(n302), 
        .Q(n295) );
  OA22X1 U829 ( .IN1(n1679), .IN2(n140), .IN3(n1551), .IN4(n98), .Q(n302) );
  MUX21X1 U830 ( .IN1(n303), .IN2(\fifo[0][12] ), .S(clear), .Q(N136) );
  NAND4X0 U831 ( .IN1(n304), .IN2(n305), .IN3(n306), .IN4(n307), .QN(n303) );
  OA221X1 U832 ( .IN1(n1936), .IN2(n122), .IN3(n1584), .IN4(n123), .IN5(n308), 
        .Q(n307) );
  OA22X1 U833 ( .IN1(n1712), .IN2(n125), .IN3(n1958), .IN4(n126), .Q(n308) );
  OA221X1 U834 ( .IN1(n1616), .IN2(n127), .IN3(n1488), .IN4(n128), .IN5(n309), 
        .Q(n306) );
  OA22X1 U835 ( .IN1(n1840), .IN2(n130), .IN3(n1744), .IN4(n131), .Q(n309) );
  OA221X1 U836 ( .IN1(n1648), .IN2(n132), .IN3(n1520), .IN4(n133), .IN5(n310), 
        .Q(n305) );
  OA22X1 U837 ( .IN1(n1872), .IN2(n135), .IN3(n1776), .IN4(n136), .Q(n310) );
  OA221X1 U838 ( .IN1(n1808), .IN2(n137), .IN3(n1904), .IN4(n138), .IN5(n311), 
        .Q(n304) );
  OA22X1 U839 ( .IN1(n1680), .IN2(n140), .IN3(n1552), .IN4(n98), .Q(n311) );
  MUX21X1 U840 ( .IN1(n312), .IN2(\fifo[0][11] ), .S(clear), .Q(N135) );
  NAND4X0 U841 ( .IN1(n313), .IN2(n314), .IN3(n315), .IN4(n316), .QN(n312) );
  OA221X1 U842 ( .IN1(n1937), .IN2(n122), .IN3(n1585), .IN4(n123), .IN5(n317), 
        .Q(n316) );
  OA22X1 U843 ( .IN1(n1713), .IN2(n125), .IN3(n1959), .IN4(n126), .Q(n317) );
  OA221X1 U844 ( .IN1(n1617), .IN2(n127), .IN3(n1489), .IN4(n128), .IN5(n318), 
        .Q(n315) );
  OA22X1 U845 ( .IN1(n1841), .IN2(n130), .IN3(n1745), .IN4(n131), .Q(n318) );
  OA221X1 U846 ( .IN1(n1649), .IN2(n132), .IN3(n1521), .IN4(n133), .IN5(n319), 
        .Q(n314) );
  OA22X1 U847 ( .IN1(n1873), .IN2(n135), .IN3(n1777), .IN4(n136), .Q(n319) );
  OA221X1 U848 ( .IN1(n1809), .IN2(n137), .IN3(n1905), .IN4(n138), .IN5(n320), 
        .Q(n313) );
  OA22X1 U849 ( .IN1(n1681), .IN2(n140), .IN3(n1553), .IN4(n98), .Q(n320) );
  MUX21X1 U850 ( .IN1(n321), .IN2(\fifo[0][10] ), .S(clear), .Q(N134) );
  NAND4X0 U851 ( .IN1(n322), .IN2(n323), .IN3(n324), .IN4(n325), .QN(n321) );
  OA221X1 U852 ( .IN1(n1938), .IN2(n122), .IN3(n1586), .IN4(n123), .IN5(n326), 
        .Q(n325) );
  OA22X1 U853 ( .IN1(n1714), .IN2(n125), .IN3(n1960), .IN4(n126), .Q(n326) );
  OA221X1 U854 ( .IN1(n1618), .IN2(n127), .IN3(n1490), .IN4(n128), .IN5(n327), 
        .Q(n324) );
  OA22X1 U855 ( .IN1(n1842), .IN2(n130), .IN3(n1746), .IN4(n131), .Q(n327) );
  OA221X1 U856 ( .IN1(n1650), .IN2(n132), .IN3(n1522), .IN4(n133), .IN5(n328), 
        .Q(n323) );
  OA22X1 U857 ( .IN1(n1874), .IN2(n135), .IN3(n1778), .IN4(n136), .Q(n328) );
  OA221X1 U858 ( .IN1(n1810), .IN2(n137), .IN3(n1906), .IN4(n138), .IN5(n329), 
        .Q(n322) );
  OA22X1 U859 ( .IN1(n1682), .IN2(n140), .IN3(n1554), .IN4(n98), .Q(n329) );
  MUX21X1 U860 ( .IN1(n330), .IN2(\fifo[0][9] ), .S(clear), .Q(N133) );
  NAND4X0 U861 ( .IN1(n331), .IN2(n332), .IN3(n333), .IN4(n334), .QN(n330) );
  OA221X1 U862 ( .IN1(n1459), .IN2(n122), .IN3(n1587), .IN4(n123), .IN5(n335), 
        .Q(n334) );
  OA22X1 U863 ( .IN1(n1715), .IN2(n125), .IN3(n1961), .IN4(n126), .Q(n335) );
  OA221X1 U864 ( .IN1(n1619), .IN2(n127), .IN3(n1491), .IN4(n128), .IN5(n336), 
        .Q(n333) );
  OA22X1 U865 ( .IN1(n1843), .IN2(n130), .IN3(n1747), .IN4(n131), .Q(n336) );
  OA221X1 U866 ( .IN1(n1651), .IN2(n132), .IN3(n1523), .IN4(n133), .IN5(n337), 
        .Q(n332) );
  OA22X1 U867 ( .IN1(n1875), .IN2(n135), .IN3(n1779), .IN4(n136), .Q(n337) );
  OA221X1 U868 ( .IN1(n1811), .IN2(n137), .IN3(n1907), .IN4(n138), .IN5(n338), 
        .Q(n331) );
  OA22X1 U869 ( .IN1(n1683), .IN2(n140), .IN3(n1555), .IN4(n98), .Q(n338) );
  MUX21X1 U870 ( .IN1(n339), .IN2(\fifo[0][8] ), .S(clear), .Q(N132) );
  NAND4X0 U871 ( .IN1(n340), .IN2(n341), .IN3(n342), .IN4(n343), .QN(n339) );
  OA221X1 U872 ( .IN1(n1460), .IN2(n122), .IN3(n1588), .IN4(n123), .IN5(n344), 
        .Q(n343) );
  OA22X1 U873 ( .IN1(n1716), .IN2(n125), .IN3(n1962), .IN4(n126), .Q(n344) );
  OA221X1 U874 ( .IN1(n1620), .IN2(n127), .IN3(n1492), .IN4(n128), .IN5(n345), 
        .Q(n342) );
  OA22X1 U875 ( .IN1(n1844), .IN2(n130), .IN3(n1748), .IN4(n131), .Q(n345) );
  OA221X1 U876 ( .IN1(n1652), .IN2(n132), .IN3(n1524), .IN4(n133), .IN5(n346), 
        .Q(n341) );
  OA22X1 U877 ( .IN1(n1876), .IN2(n135), .IN3(n1780), .IN4(n136), .Q(n346) );
  OA221X1 U878 ( .IN1(n1812), .IN2(n137), .IN3(n1908), .IN4(n138), .IN5(n347), 
        .Q(n340) );
  OA22X1 U879 ( .IN1(n1684), .IN2(n140), .IN3(n1556), .IN4(n98), .Q(n347) );
  MUX21X1 U880 ( .IN1(n348), .IN2(\fifo[0][7] ), .S(clear), .Q(N131) );
  NAND4X0 U881 ( .IN1(n349), .IN2(n350), .IN3(n351), .IN4(n352), .QN(n348) );
  OA221X1 U882 ( .IN1(n1461), .IN2(n122), .IN3(n1589), .IN4(n123), .IN5(n353), 
        .Q(n352) );
  OA22X1 U883 ( .IN1(n1717), .IN2(n125), .IN3(n1963), .IN4(n126), .Q(n353) );
  OA221X1 U884 ( .IN1(n1621), .IN2(n127), .IN3(n1493), .IN4(n128), .IN5(n354), 
        .Q(n351) );
  OA22X1 U885 ( .IN1(n1845), .IN2(n130), .IN3(n1749), .IN4(n131), .Q(n354) );
  OA221X1 U886 ( .IN1(n1653), .IN2(n132), .IN3(n1525), .IN4(n133), .IN5(n355), 
        .Q(n350) );
  OA22X1 U887 ( .IN1(n1877), .IN2(n135), .IN3(n1781), .IN4(n136), .Q(n355) );
  OA221X1 U888 ( .IN1(n1813), .IN2(n137), .IN3(n1909), .IN4(n138), .IN5(n356), 
        .Q(n349) );
  OA22X1 U889 ( .IN1(n1685), .IN2(n140), .IN3(n1557), .IN4(n98), .Q(n356) );
  MUX21X1 U890 ( .IN1(n357), .IN2(\fifo[0][6] ), .S(clear), .Q(N130) );
  NAND4X0 U891 ( .IN1(n358), .IN2(n359), .IN3(n360), .IN4(n361), .QN(n357) );
  OA221X1 U892 ( .IN1(n1462), .IN2(n122), .IN3(n1590), .IN4(n123), .IN5(n362), 
        .Q(n361) );
  OA22X1 U893 ( .IN1(n1718), .IN2(n125), .IN3(n1964), .IN4(n126), .Q(n362) );
  OA221X1 U894 ( .IN1(n1622), .IN2(n127), .IN3(n1494), .IN4(n128), .IN5(n363), 
        .Q(n360) );
  OA22X1 U895 ( .IN1(n1846), .IN2(n130), .IN3(n1750), .IN4(n131), .Q(n363) );
  OA221X1 U896 ( .IN1(n1654), .IN2(n132), .IN3(n1526), .IN4(n133), .IN5(n364), 
        .Q(n359) );
  OA22X1 U897 ( .IN1(n1878), .IN2(n135), .IN3(n1782), .IN4(n136), .Q(n364) );
  OA221X1 U898 ( .IN1(n1814), .IN2(n137), .IN3(n1910), .IN4(n138), .IN5(n365), 
        .Q(n358) );
  OA22X1 U899 ( .IN1(n1686), .IN2(n140), .IN3(n1558), .IN4(n98), .Q(n365) );
  MUX21X1 U900 ( .IN1(n366), .IN2(\fifo[0][5] ), .S(clear), .Q(N129) );
  NAND4X0 U901 ( .IN1(n367), .IN2(n368), .IN3(n369), .IN4(n370), .QN(n366) );
  OA221X1 U902 ( .IN1(n1463), .IN2(n122), .IN3(n1591), .IN4(n123), .IN5(n371), 
        .Q(n370) );
  OA22X1 U903 ( .IN1(n1719), .IN2(n125), .IN3(n1965), .IN4(n126), .Q(n371) );
  OA221X1 U904 ( .IN1(n1623), .IN2(n127), .IN3(n1495), .IN4(n128), .IN5(n372), 
        .Q(n369) );
  OA22X1 U905 ( .IN1(n1847), .IN2(n130), .IN3(n1751), .IN4(n131), .Q(n372) );
  OA221X1 U906 ( .IN1(n1655), .IN2(n132), .IN3(n1527), .IN4(n133), .IN5(n373), 
        .Q(n368) );
  OA22X1 U907 ( .IN1(n1879), .IN2(n135), .IN3(n1783), .IN4(n136), .Q(n373) );
  OA221X1 U908 ( .IN1(n1815), .IN2(n137), .IN3(n1911), .IN4(n138), .IN5(n374), 
        .Q(n367) );
  OA22X1 U909 ( .IN1(n1687), .IN2(n140), .IN3(n1559), .IN4(n98), .Q(n374) );
  MUX21X1 U910 ( .IN1(n375), .IN2(\fifo[0][4] ), .S(clear), .Q(N128) );
  NAND4X0 U911 ( .IN1(n376), .IN2(n377), .IN3(n378), .IN4(n379), .QN(n375) );
  OA221X1 U912 ( .IN1(n1464), .IN2(n122), .IN3(n1592), .IN4(n123), .IN5(n380), 
        .Q(n379) );
  OA22X1 U913 ( .IN1(n1720), .IN2(n125), .IN3(n1966), .IN4(n126), .Q(n380) );
  OA221X1 U914 ( .IN1(n1624), .IN2(n127), .IN3(n1496), .IN4(n128), .IN5(n381), 
        .Q(n378) );
  OA22X1 U915 ( .IN1(n1848), .IN2(n130), .IN3(n1752), .IN4(n131), .Q(n381) );
  OA221X1 U916 ( .IN1(n1656), .IN2(n132), .IN3(n1528), .IN4(n133), .IN5(n382), 
        .Q(n377) );
  OA22X1 U917 ( .IN1(n1880), .IN2(n135), .IN3(n1784), .IN4(n136), .Q(n382) );
  OA221X1 U918 ( .IN1(n1816), .IN2(n137), .IN3(n1912), .IN4(n138), .IN5(n383), 
        .Q(n376) );
  OA22X1 U919 ( .IN1(n1688), .IN2(n140), .IN3(n1560), .IN4(n98), .Q(n383) );
  MUX21X1 U920 ( .IN1(n384), .IN2(\fifo[0][3] ), .S(clear), .Q(N127) );
  NAND4X0 U921 ( .IN1(n385), .IN2(n386), .IN3(n387), .IN4(n388), .QN(n384) );
  OA221X1 U922 ( .IN1(n1465), .IN2(n122), .IN3(n1593), .IN4(n123), .IN5(n389), 
        .Q(n388) );
  OA22X1 U923 ( .IN1(n1721), .IN2(n125), .IN3(n1967), .IN4(n126), .Q(n389) );
  OA221X1 U924 ( .IN1(n1625), .IN2(n127), .IN3(n1497), .IN4(n128), .IN5(n390), 
        .Q(n387) );
  OA22X1 U925 ( .IN1(n1849), .IN2(n130), .IN3(n1753), .IN4(n131), .Q(n390) );
  OA221X1 U926 ( .IN1(n1657), .IN2(n132), .IN3(n1529), .IN4(n133), .IN5(n391), 
        .Q(n386) );
  OA22X1 U927 ( .IN1(n1881), .IN2(n135), .IN3(n1785), .IN4(n136), .Q(n391) );
  OA221X1 U928 ( .IN1(n1817), .IN2(n137), .IN3(n1913), .IN4(n138), .IN5(n392), 
        .Q(n385) );
  OA22X1 U929 ( .IN1(n1689), .IN2(n140), .IN3(n1561), .IN4(n98), .Q(n392) );
  MUX21X1 U930 ( .IN1(n393), .IN2(\fifo[0][2] ), .S(clear), .Q(N126) );
  NAND4X0 U931 ( .IN1(n394), .IN2(n395), .IN3(n396), .IN4(n397), .QN(n393) );
  OA221X1 U932 ( .IN1(n1466), .IN2(n122), .IN3(n1594), .IN4(n123), .IN5(n398), 
        .Q(n397) );
  OA22X1 U933 ( .IN1(n1722), .IN2(n125), .IN3(n1968), .IN4(n126), .Q(n398) );
  OA221X1 U934 ( .IN1(n1626), .IN2(n127), .IN3(n1498), .IN4(n128), .IN5(n399), 
        .Q(n396) );
  OA22X1 U935 ( .IN1(n1850), .IN2(n130), .IN3(n1754), .IN4(n131), .Q(n399) );
  OA221X1 U936 ( .IN1(n1658), .IN2(n132), .IN3(n1530), .IN4(n133), .IN5(n400), 
        .Q(n395) );
  OA22X1 U937 ( .IN1(n1882), .IN2(n135), .IN3(n1786), .IN4(n136), .Q(n400) );
  OA221X1 U938 ( .IN1(n1818), .IN2(n137), .IN3(n1914), .IN4(n138), .IN5(n401), 
        .Q(n394) );
  OA22X1 U939 ( .IN1(n1690), .IN2(n140), .IN3(n1562), .IN4(n98), .Q(n401) );
  MUX21X1 U940 ( .IN1(n402), .IN2(\fifo[0][1] ), .S(clear), .Q(N125) );
  NAND4X0 U941 ( .IN1(n403), .IN2(n404), .IN3(n405), .IN4(n406), .QN(n402) );
  OA221X1 U942 ( .IN1(n1467), .IN2(n122), .IN3(n1595), .IN4(n123), .IN5(n407), 
        .Q(n406) );
  OA22X1 U943 ( .IN1(n1723), .IN2(n125), .IN3(n1969), .IN4(n126), .Q(n407) );
  OA221X1 U944 ( .IN1(n1627), .IN2(n127), .IN3(n1499), .IN4(n128), .IN5(n408), 
        .Q(n405) );
  OA22X1 U945 ( .IN1(n1851), .IN2(n130), .IN3(n1755), .IN4(n131), .Q(n408) );
  OA221X1 U946 ( .IN1(n1659), .IN2(n132), .IN3(n1531), .IN4(n133), .IN5(n409), 
        .Q(n404) );
  OA22X1 U947 ( .IN1(n1883), .IN2(n135), .IN3(n1787), .IN4(n136), .Q(n409) );
  OA221X1 U948 ( .IN1(n1819), .IN2(n137), .IN3(n1915), .IN4(n138), .IN5(n410), 
        .Q(n403) );
  OA22X1 U949 ( .IN1(n1691), .IN2(n140), .IN3(n1563), .IN4(n98), .Q(n410) );
  MUX21X1 U950 ( .IN1(n411), .IN2(\fifo[0][0] ), .S(clear), .Q(N124) );
  NAND4X0 U951 ( .IN1(n412), .IN2(n413), .IN3(n414), .IN4(n415), .QN(n411) );
  OA221X1 U952 ( .IN1(n1468), .IN2(n122), .IN3(n1596), .IN4(n123), .IN5(n416), 
        .Q(n415) );
  OA22X1 U953 ( .IN1(n1724), .IN2(n125), .IN3(n1970), .IN4(n126), .Q(n416) );
  NAND2X0 U954 ( .IN1(n417), .IN2(n418), .QN(n126) );
  NAND2X0 U955 ( .IN1(n419), .IN2(n418), .QN(n125) );
  NAND2X0 U956 ( .IN1(n420), .IN2(n418), .QN(n123) );
  NAND2X0 U957 ( .IN1(n418), .IN2(n421), .QN(n122) );
  NOR2X0 U958 ( .IN1(N15), .IN2(n2), .QN(n418) );
  OA221X1 U959 ( .IN1(n1628), .IN2(n127), .IN3(n1500), .IN4(n128), .IN5(n422), 
        .Q(n414) );
  OA22X1 U960 ( .IN1(n1852), .IN2(n130), .IN3(n1756), .IN4(n131), .Q(n422) );
  NAND2X0 U961 ( .IN1(n92), .IN2(n419), .QN(n131) );
  NAND2X0 U962 ( .IN1(n92), .IN2(n417), .QN(n130) );
  NAND2X0 U963 ( .IN1(n92), .IN2(n421), .QN(n128) );
  NAND2X0 U964 ( .IN1(n92), .IN2(n420), .QN(n127) );
  NOR2X0 U965 ( .IN1(N15), .IN2(n588), .QN(n92) );
  OA221X1 U966 ( .IN1(n1660), .IN2(n132), .IN3(n1532), .IN4(n133), .IN5(n423), 
        .Q(n413) );
  OA22X1 U967 ( .IN1(n1884), .IN2(n135), .IN3(n1788), .IN4(n136), .Q(n423) );
  NAND2X0 U968 ( .IN1(n91), .IN2(n419), .QN(n136) );
  NAND2X0 U969 ( .IN1(n91), .IN2(n417), .QN(n135) );
  NAND2X0 U970 ( .IN1(n91), .IN2(n421), .QN(n133) );
  NAND2X0 U971 ( .IN1(n91), .IN2(n420), .QN(n132) );
  NOR2X0 U972 ( .IN1(n2), .IN2(n587), .QN(n91) );
  OA221X1 U973 ( .IN1(n1820), .IN2(n137), .IN3(n1916), .IN4(n138), .IN5(n424), 
        .Q(n412) );
  OA22X1 U974 ( .IN1(n1692), .IN2(n140), .IN3(n1564), .IN4(n98), .Q(n424) );
  NAND2X0 U975 ( .IN1(n421), .IN2(n425), .QN(n98) );
  NOR2X0 U976 ( .IN1(N17), .IN2(n586), .QN(n421) );
  NAND2X0 U977 ( .IN1(n420), .IN2(n425), .QN(n140) );
  INVX0 U978 ( .INP(n99), .ZN(n420) );
  NAND2X0 U979 ( .IN1(n586), .IN2(N17), .QN(n99) );
  NAND2X0 U980 ( .IN1(n417), .IN2(n425), .QN(n138) );
  AND2X1 U981 ( .IN1(n585), .IN2(n586), .Q(n417) );
  NAND2X0 U982 ( .IN1(n419), .IN2(n425), .QN(n137) );
  INVX0 U983 ( .INP(n96), .ZN(n425) );
  NAND2X0 U984 ( .IN1(n2), .IN2(N15), .QN(n96) );
  NOR2X0 U985 ( .IN1(n586), .IN2(n585), .QN(n419) );
endmodule


module eth_fifo_DATA_WIDTH32_DEPTH16_CNT_WIDTH5_test_1 ( data_in, data_out, 
        clk, reset, write, read, clear, almost_full, full, almost_empty, empty, 
        cnt, eth_top_test_point_11887_in, test_si2, test_si1, test_so1, 
        test_se );
  input [31:0] data_in;
  output [31:0] data_out;
  output [4:0] cnt;
  input clk, reset, write, read, clear, eth_top_test_point_11887_in, test_si2,
         test_si1, test_se;
  output almost_full, full, almost_empty, empty, test_so1;
  wire   N15, N16, N17, \fifo[0][31] , \fifo[0][30] , \fifo[0][29] ,
         \fifo[0][28] , \fifo[0][27] , \fifo[0][26] , \fifo[0][25] ,
         \fifo[0][24] , \fifo[0][23] , \fifo[0][22] , \fifo[0][21] ,
         \fifo[0][20] , \fifo[0][19] , \fifo[0][18] , \fifo[0][17] ,
         \fifo[0][16] , \fifo[0][15] , \fifo[0][14] , \fifo[0][13] ,
         \fifo[0][12] , \fifo[0][11] , \fifo[0][10] , \fifo[0][9] ,
         \fifo[0][8] , \fifo[0][7] , \fifo[0][6] , \fifo[0][5] , \fifo[0][4] ,
         \fifo[0][3] , \fifo[0][2] , \fifo[0][1] , \fifo[0][0] , \fifo[1][31] ,
         \fifo[1][30] , \fifo[1][29] , \fifo[1][28] , \fifo[1][27] ,
         \fifo[1][26] , \fifo[1][25] , \fifo[1][24] , \fifo[1][23] ,
         \fifo[1][22] , \fifo[1][21] , \fifo[1][20] , \fifo[1][19] ,
         \fifo[1][18] , \fifo[1][17] , \fifo[1][16] , \fifo[1][15] ,
         \fifo[1][14] , \fifo[1][13] , \fifo[1][12] , \fifo[1][11] ,
         \fifo[1][10] , \fifo[1][9] , \fifo[1][8] , \fifo[1][7] , \fifo[1][6] ,
         \fifo[1][5] , \fifo[1][4] , \fifo[1][3] , \fifo[1][2] , \fifo[1][1] ,
         \fifo[1][0] , \fifo[2][31] , \fifo[2][30] , \fifo[2][29] ,
         \fifo[2][28] , \fifo[2][27] , \fifo[2][26] , \fifo[2][25] ,
         \fifo[2][24] , \fifo[2][23] , \fifo[2][22] , \fifo[2][21] ,
         \fifo[2][20] , \fifo[2][19] , \fifo[2][18] , \fifo[2][17] ,
         \fifo[2][16] , \fifo[2][15] , \fifo[2][14] , \fifo[2][13] ,
         \fifo[2][12] , \fifo[2][11] , \fifo[2][10] , \fifo[2][9] ,
         \fifo[2][8] , \fifo[2][7] , \fifo[2][6] , \fifo[2][5] , \fifo[2][4] ,
         \fifo[2][3] , \fifo[2][2] , \fifo[2][1] , \fifo[2][0] , \fifo[3][31] ,
         \fifo[3][30] , \fifo[3][29] , \fifo[3][28] , \fifo[3][27] ,
         \fifo[3][26] , \fifo[3][25] , \fifo[3][24] , \fifo[3][23] ,
         \fifo[3][22] , \fifo[3][21] , \fifo[3][20] , \fifo[3][19] ,
         \fifo[3][18] , \fifo[3][17] , \fifo[3][16] , \fifo[3][15] ,
         \fifo[3][14] , \fifo[3][13] , \fifo[3][12] , \fifo[3][11] ,
         \fifo[3][10] , \fifo[3][9] , \fifo[3][8] , \fifo[3][7] , \fifo[3][6] ,
         \fifo[3][5] , \fifo[3][4] , \fifo[3][3] , \fifo[3][2] , \fifo[3][1] ,
         \fifo[3][0] , \fifo[4][31] , \fifo[4][30] , \fifo[4][29] ,
         \fifo[4][28] , \fifo[4][27] , \fifo[4][26] , \fifo[4][25] ,
         \fifo[4][24] , \fifo[4][23] , \fifo[4][22] , \fifo[4][21] ,
         \fifo[4][20] , \fifo[4][19] , \fifo[4][18] , \fifo[4][17] ,
         \fifo[4][16] , \fifo[4][15] , \fifo[4][14] , \fifo[4][13] ,
         \fifo[4][12] , \fifo[4][11] , \fifo[4][10] , \fifo[4][9] ,
         \fifo[4][8] , \fifo[4][7] , \fifo[4][6] , \fifo[4][5] , \fifo[4][4] ,
         \fifo[4][3] , \fifo[4][2] , \fifo[4][1] , \fifo[4][0] , \fifo[5][31] ,
         \fifo[5][30] , \fifo[5][29] , \fifo[5][28] , \fifo[5][27] ,
         \fifo[5][26] , \fifo[5][25] , \fifo[5][24] , \fifo[5][23] ,
         \fifo[5][22] , \fifo[5][21] , \fifo[5][20] , \fifo[5][19] ,
         \fifo[5][18] , \fifo[5][17] , \fifo[5][16] , \fifo[5][15] ,
         \fifo[5][14] , \fifo[5][13] , \fifo[5][12] , \fifo[5][11] ,
         \fifo[5][10] , \fifo[5][9] , \fifo[5][8] , \fifo[5][7] , \fifo[5][6] ,
         \fifo[5][5] , \fifo[5][4] , \fifo[5][3] , \fifo[5][2] , \fifo[5][1] ,
         \fifo[5][0] , \fifo[6][31] , \fifo[6][30] , \fifo[6][29] ,
         \fifo[6][28] , \fifo[6][27] , \fifo[6][26] , \fifo[6][25] ,
         \fifo[6][24] , \fifo[6][23] , \fifo[6][22] , \fifo[6][21] ,
         \fifo[6][20] , \fifo[6][19] , \fifo[6][18] , \fifo[6][17] ,
         \fifo[6][16] , \fifo[6][15] , \fifo[6][14] , \fifo[6][13] ,
         \fifo[6][12] , \fifo[6][11] , \fifo[6][10] , \fifo[6][9] ,
         \fifo[6][8] , \fifo[6][7] , \fifo[6][6] , \fifo[6][5] , \fifo[6][4] ,
         \fifo[6][3] , \fifo[6][2] , \fifo[6][1] , \fifo[6][0] , \fifo[7][31] ,
         \fifo[7][30] , \fifo[7][29] , \fifo[7][28] , \fifo[7][27] ,
         \fifo[7][26] , \fifo[7][25] , \fifo[7][24] , \fifo[7][23] ,
         \fifo[7][22] , \fifo[7][21] , \fifo[7][20] , \fifo[7][19] ,
         \fifo[7][18] , \fifo[7][17] , \fifo[7][16] , \fifo[7][15] ,
         \fifo[7][14] , \fifo[7][13] , \fifo[7][12] , \fifo[7][11] ,
         \fifo[7][10] , \fifo[7][9] , \fifo[7][8] , \fifo[7][7] , \fifo[7][6] ,
         \fifo[7][5] , \fifo[7][4] , \fifo[7][3] , \fifo[7][2] , \fifo[7][1] ,
         \fifo[7][0] , \fifo[8][31] , \fifo[8][30] , \fifo[8][29] ,
         \fifo[8][28] , \fifo[8][27] , \fifo[8][26] , \fifo[8][25] ,
         \fifo[8][24] , \fifo[8][23] , \fifo[8][22] , \fifo[8][21] ,
         \fifo[8][20] , \fifo[8][19] , \fifo[8][18] , \fifo[8][17] ,
         \fifo[8][16] , \fifo[8][15] , \fifo[8][14] , \fifo[8][13] ,
         \fifo[8][12] , \fifo[8][11] , \fifo[8][10] , \fifo[8][9] ,
         \fifo[8][8] , \fifo[8][7] , \fifo[8][6] , \fifo[8][5] , \fifo[8][4] ,
         \fifo[8][3] , \fifo[8][2] , \fifo[8][1] , \fifo[8][0] , \fifo[9][31] ,
         \fifo[9][30] , \fifo[9][29] , \fifo[9][28] , \fifo[9][27] ,
         \fifo[9][26] , \fifo[9][25] , \fifo[9][24] , \fifo[9][23] ,
         \fifo[9][22] , \fifo[9][21] , \fifo[9][20] , \fifo[9][19] ,
         \fifo[9][18] , \fifo[9][17] , \fifo[9][16] , \fifo[9][15] ,
         \fifo[9][14] , \fifo[9][13] , \fifo[9][12] , \fifo[9][11] ,
         \fifo[9][10] , \fifo[9][9] , \fifo[9][8] , \fifo[9][7] , \fifo[9][6] ,
         \fifo[9][5] , \fifo[9][4] , \fifo[9][3] , \fifo[9][2] , \fifo[9][1] ,
         \fifo[9][0] , \fifo[10][31] , \fifo[10][30] , \fifo[10][29] ,
         \fifo[10][28] , \fifo[10][27] , \fifo[10][26] , \fifo[10][25] ,
         \fifo[10][24] , \fifo[10][23] , \fifo[10][22] , \fifo[10][21] ,
         \fifo[10][20] , \fifo[10][19] , \fifo[10][18] , \fifo[10][17] ,
         \fifo[10][16] , \fifo[10][15] , \fifo[10][14] , \fifo[10][13] ,
         \fifo[10][12] , \fifo[10][11] , \fifo[10][10] , \fifo[10][9] ,
         \fifo[10][8] , \fifo[10][7] , \fifo[10][6] , \fifo[10][5] ,
         \fifo[10][4] , \fifo[10][3] , \fifo[10][2] , \fifo[10][1] ,
         \fifo[10][0] , \fifo[11][31] , \fifo[11][30] , \fifo[11][29] ,
         \fifo[11][28] , \fifo[11][27] , \fifo[11][26] , \fifo[11][25] ,
         \fifo[11][24] , \fifo[11][23] , \fifo[11][22] , \fifo[11][21] ,
         \fifo[11][20] , \fifo[11][19] , \fifo[11][18] , \fifo[11][17] ,
         \fifo[11][16] , \fifo[11][15] , \fifo[11][14] , \fifo[11][13] ,
         \fifo[11][12] , \fifo[11][11] , \fifo[11][10] , \fifo[11][9] ,
         \fifo[11][8] , \fifo[11][7] , \fifo[11][6] , \fifo[11][5] ,
         \fifo[11][4] , \fifo[11][3] , \fifo[11][2] , \fifo[11][1] ,
         \fifo[11][0] , \fifo[12][31] , \fifo[12][30] , \fifo[12][29] ,
         \fifo[12][28] , \fifo[12][27] , \fifo[12][26] , \fifo[12][25] ,
         \fifo[12][24] , \fifo[12][23] , \fifo[12][22] , \fifo[12][21] ,
         \fifo[12][20] , \fifo[12][19] , \fifo[12][18] , \fifo[12][17] ,
         \fifo[12][16] , \fifo[12][15] , \fifo[12][14] , \fifo[12][13] ,
         \fifo[12][12] , \fifo[12][11] , \fifo[12][10] , \fifo[12][9] ,
         \fifo[12][8] , \fifo[12][7] , \fifo[12][6] , \fifo[12][5] ,
         \fifo[12][4] , \fifo[12][3] , \fifo[12][2] , \fifo[12][1] ,
         \fifo[12][0] , \fifo[13][31] , \fifo[13][30] , \fifo[13][29] ,
         \fifo[13][28] , \fifo[13][27] , \fifo[13][26] , \fifo[13][25] ,
         \fifo[13][24] , \fifo[13][23] , \fifo[13][22] , \fifo[13][21] ,
         \fifo[13][20] , \fifo[13][19] , \fifo[13][18] , \fifo[13][17] ,
         \fifo[13][16] , \fifo[13][15] , \fifo[13][14] , \fifo[13][13] ,
         \fifo[13][12] , \fifo[13][11] , \fifo[13][10] , \fifo[13][9] ,
         \fifo[13][8] , \fifo[13][7] , \fifo[13][6] , \fifo[13][5] ,
         \fifo[13][4] , \fifo[13][3] , \fifo[13][2] , \fifo[13][1] ,
         \fifo[13][0] , \fifo[14][31] , \fifo[14][30] , \fifo[14][29] ,
         \fifo[14][28] , \fifo[14][27] , \fifo[14][26] , \fifo[14][25] ,
         \fifo[14][24] , \fifo[14][23] , \fifo[14][22] , \fifo[14][21] ,
         \fifo[14][20] , \fifo[14][19] , \fifo[14][18] , \fifo[14][17] ,
         \fifo[14][16] , \fifo[14][15] , \fifo[14][14] , \fifo[14][13] ,
         \fifo[14][12] , \fifo[14][11] , \fifo[14][10] , \fifo[14][9] ,
         \fifo[14][8] , \fifo[14][7] , \fifo[14][6] , \fifo[14][5] ,
         \fifo[14][4] , \fifo[14][3] , \fifo[14][2] , \fifo[14][1] ,
         \fifo[14][0] , \fifo[15][31] , \fifo[15][30] , \fifo[15][29] ,
         \fifo[15][28] , \fifo[15][27] , \fifo[15][26] , \fifo[15][25] ,
         \fifo[15][24] , \fifo[15][23] , \fifo[15][22] , \fifo[15][21] ,
         \fifo[15][20] , \fifo[15][19] , \fifo[15][18] , \fifo[15][17] ,
         \fifo[15][16] , \fifo[15][15] , \fifo[15][14] , \fifo[15][13] ,
         \fifo[15][12] , \fifo[15][11] , \fifo[15][10] , \fifo[15][9] ,
         \fifo[15][8] , \fifo[15][7] , \fifo[15][6] , \fifo[15][5] ,
         \fifo[15][4] , \fifo[15][3] , \fifo[15][2] , \fifo[15][1] ,
         \fifo[15][0] , N124, N125, N126, N127, N128, N129, N130, N131, N132,
         N133, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, \U3/U1/Z_0 , n2, n1311, n1312, n1313, n1318, n1319, n1320,
         n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
         n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
         n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
         n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
         n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
         n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
         n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
         n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
         n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
         n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
         n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
         n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
         n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
         n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
         n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
         n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
         n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
         n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
         n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
         n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
         n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
         n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
         n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
         n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
         n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
         n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
         n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
         n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
         n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
         n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
         n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
         n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
         n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
         n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
         n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
         n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
         n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
         n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
         n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
         n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
         n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
         n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740,
         n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750,
         n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
         n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
         n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
         n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
         n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
         n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
         n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
         n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
         n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
         n1841, n1842, n1844, n1845, n1846, n1847, n1848, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
         n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1314,
         n1315, n1316, n1317, n1843, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n428;
  wire   [3:0] write_pointer;
  assign test_so1 = write_pointer[3];
  assign \U3/U1/Z_0  = read;

  SDFFARX1 \cnt_reg[0]  ( .D(n1318), .SI(test_si1), .SE(test_se), .CLK(n5), 
        .RSTB(n428), .Q(cnt[0]), .QN(n1311) );
  SDFFARX1 \cnt_reg[1]  ( .D(n1319), .SI(cnt[0]), .SE(test_se), .CLK(n5), 
        .RSTB(n428), .Q(cnt[1]), .QN(n1847) );
  SDFFARX1 \cnt_reg[2]  ( .D(n1320), .SI(cnt[1]), .SE(test_se), .CLK(n5), 
        .RSTB(n428), .Q(cnt[2]), .QN(n1312) );
  SDFFARX1 \cnt_reg[3]  ( .D(n1321), .SI(cnt[2]), .SE(test_se), .CLK(n5), 
        .RSTB(n428), .Q(cnt[3]), .QN(n1313) );
  SDFFARX1 \cnt_reg[4]  ( .D(n1322), .SI(cnt[3]), .SE(test_se), .CLK(n5), 
        .RSTB(n428), .Q(cnt[4]), .QN(n1848) );
  SDFFARX1 \read_pointer_reg[0]  ( .D(n1323), .SI(\fifo[15][31] ), .SE(test_se), .CLK(n5), .RSTB(n428), .Q(n2), .QN(n426) );
  SDFFARX1 \read_pointer_reg[1]  ( .D(n1324), .SI(n2), .SE(test_se), .CLK(n6), 
        .RSTB(n428), .Q(N15), .QN(n1844) );
  SDFFARX1 \read_pointer_reg[2]  ( .D(n1325), .SI(N15), .SE(test_se), .CLK(n5), 
        .RSTB(n428), .Q(N16), .QN(n1845) );
  SDFFARX1 \read_pointer_reg[3]  ( .D(n1326), .SI(N16), .SE(test_se), .CLK(n5), 
        .RSTB(n428), .Q(N17), .QN(n1846) );
  SDFFARX1 \write_pointer_reg[0]  ( .D(n1327), .SI(N17), .SE(test_se), .CLK(n5), .RSTB(n428), .Q(write_pointer[0]) );
  SDFFARX1 \write_pointer_reg[1]  ( .D(n1328), .SI(write_pointer[0]), .SE(
        test_se), .CLK(n5), .RSTB(n428), .Q(write_pointer[1]), .QN(n4) );
  SDFFARX1 \write_pointer_reg[2]  ( .D(n1329), .SI(write_pointer[1]), .SE(
        test_se), .CLK(n5), .RSTB(n428), .Q(write_pointer[2]), .QN(n1) );
  SDFFARX1 \write_pointer_reg[3]  ( .D(n1330), .SI(write_pointer[2]), .SE(
        test_se), .CLK(n5), .RSTB(n428), .Q(write_pointer[3]), .QN(n3) );
  SDFFX1 \fifo_reg[0][31]  ( .D(n1331), .SI(\fifo[0][30] ), .SE(test_se), 
        .CLK(n20), .Q(\fifo[0][31] ), .QN(n1935) );
  SDFFX1 \fifo_reg[0][30]  ( .D(n1332), .SI(\fifo[0][29] ), .SE(test_se), 
        .CLK(n35), .Q(\fifo[0][30] ), .QN(n1936) );
  SDFFX1 \fifo_reg[0][29]  ( .D(n1333), .SI(\fifo[0][28] ), .SE(test_se), 
        .CLK(n35), .Q(\fifo[0][29] ), .QN(n1937) );
  SDFFX1 \fifo_reg[0][28]  ( .D(n1334), .SI(\fifo[0][27] ), .SE(test_se), 
        .CLK(n34), .Q(\fifo[0][28] ), .QN(n1938) );
  SDFFX1 \fifo_reg[0][27]  ( .D(n1335), .SI(\fifo[0][26] ), .SE(test_se), 
        .CLK(n34), .Q(\fifo[0][27] ), .QN(n1939) );
  SDFFX1 \fifo_reg[0][26]  ( .D(n1336), .SI(\fifo[0][25] ), .SE(test_se), 
        .CLK(n34), .Q(\fifo[0][26] ), .QN(n1940) );
  SDFFX1 \fifo_reg[0][25]  ( .D(n1337), .SI(\fifo[0][24] ), .SE(test_se), 
        .CLK(n34), .Q(\fifo[0][25] ), .QN(n1941) );
  SDFFX1 \fifo_reg[0][24]  ( .D(n1338), .SI(\fifo[0][23] ), .SE(test_se), 
        .CLK(n34), .Q(\fifo[0][24] ), .QN(n1942) );
  SDFFX1 \fifo_reg[0][23]  ( .D(n1339), .SI(\fifo[0][22] ), .SE(test_se), 
        .CLK(n34), .Q(\fifo[0][23] ), .QN(n1943) );
  SDFFX1 \fifo_reg[0][22]  ( .D(n1340), .SI(\fifo[0][21] ), .SE(test_se), 
        .CLK(n34), .Q(\fifo[0][22] ), .QN(n1944) );
  SDFFX1 \fifo_reg[0][21]  ( .D(n1341), .SI(\fifo[0][20] ), .SE(test_se), 
        .CLK(n34), .Q(\fifo[0][21] ), .QN(n1945) );
  SDFFX1 \fifo_reg[0][20]  ( .D(n1342), .SI(\fifo[0][19] ), .SE(test_se), 
        .CLK(n34), .Q(\fifo[0][20] ), .QN(n1946) );
  SDFFX1 \fifo_reg[0][19]  ( .D(n1343), .SI(\fifo[0][18] ), .SE(test_se), 
        .CLK(n34), .Q(\fifo[0][19] ), .QN(n1947) );
  SDFFX1 \fifo_reg[0][18]  ( .D(n1344), .SI(\fifo[0][17] ), .SE(test_se), 
        .CLK(n34), .Q(\fifo[0][18] ), .QN(n1948) );
  SDFFX1 \fifo_reg[0][17]  ( .D(n1345), .SI(\fifo[0][16] ), .SE(test_se), 
        .CLK(n34), .Q(\fifo[0][17] ), .QN(n1949) );
  SDFFX1 \fifo_reg[0][16]  ( .D(n1346), .SI(\fifo[0][15] ), .SE(test_se), 
        .CLK(n34), .Q(\fifo[0][16] ), .QN(n1950) );
  SDFFX1 \fifo_reg[0][15]  ( .D(n1347), .SI(\fifo[0][14] ), .SE(test_se), 
        .CLK(n34), .Q(\fifo[0][15] ), .QN(n1951) );
  SDFFX1 \fifo_reg[0][14]  ( .D(n1348), .SI(\fifo[0][13] ), .SE(test_se), 
        .CLK(n33), .Q(\fifo[0][14] ), .QN(n1952) );
  SDFFX1 \fifo_reg[0][13]  ( .D(n1349), .SI(\fifo[0][12] ), .SE(test_se), 
        .CLK(n33), .Q(\fifo[0][13] ), .QN(n1953) );
  SDFFX1 \fifo_reg[0][12]  ( .D(n1350), .SI(\fifo[0][11] ), .SE(test_se), 
        .CLK(n33), .Q(\fifo[0][12] ), .QN(n1954) );
  SDFFX1 \fifo_reg[0][11]  ( .D(n1351), .SI(\fifo[0][10] ), .SE(test_se), 
        .CLK(n33), .Q(\fifo[0][11] ), .QN(n1955) );
  SDFFX1 \fifo_reg[0][10]  ( .D(n1352), .SI(\fifo[0][9] ), .SE(test_se), .CLK(
        n33), .Q(\fifo[0][10] ), .QN(n1956) );
  SDFFX1 \fifo_reg[0][9]  ( .D(n1353), .SI(\fifo[0][8] ), .SE(test_se), .CLK(
        n33), .Q(\fifo[0][9] ), .QN(n1957) );
  SDFFX1 \fifo_reg[0][8]  ( .D(n1354), .SI(\fifo[0][7] ), .SE(test_se), .CLK(
        n33), .Q(\fifo[0][8] ), .QN(n1958) );
  SDFFX1 \fifo_reg[0][7]  ( .D(n1355), .SI(\fifo[0][6] ), .SE(test_se), .CLK(
        n33), .Q(\fifo[0][7] ), .QN(n1959) );
  SDFFX1 \fifo_reg[0][6]  ( .D(n1356), .SI(\fifo[0][5] ), .SE(test_se), .CLK(
        n33), .Q(\fifo[0][6] ), .QN(n1960) );
  SDFFX1 \fifo_reg[0][5]  ( .D(n1357), .SI(\fifo[0][4] ), .SE(test_se), .CLK(
        n33), .Q(\fifo[0][5] ), .QN(n1961) );
  SDFFX1 \fifo_reg[0][4]  ( .D(n1358), .SI(\fifo[0][3] ), .SE(test_se), .CLK(
        n33), .Q(\fifo[0][4] ), .QN(n1962) );
  SDFFX1 \fifo_reg[0][3]  ( .D(n1359), .SI(\fifo[0][2] ), .SE(test_se), .CLK(
        n33), .Q(\fifo[0][3] ), .QN(n1963) );
  SDFFX1 \fifo_reg[0][2]  ( .D(n1360), .SI(\fifo[0][1] ), .SE(test_se), .CLK(
        n33), .Q(\fifo[0][2] ), .QN(n1964) );
  SDFFX1 \fifo_reg[0][1]  ( .D(n1361), .SI(\fifo[0][0] ), .SE(test_se), .CLK(
        n33), .Q(\fifo[0][1] ), .QN(n1965) );
  SDFFX1 \fifo_reg[0][0]  ( .D(n1362), .SI(data_out[30]), .SE(test_se), .CLK(
        n32), .Q(\fifo[0][0] ), .QN(n1966) );
  SDFFX1 \fifo_reg[1][31]  ( .D(n1363), .SI(\fifo[1][30] ), .SE(test_se), 
        .CLK(n17), .Q(\fifo[1][31] ), .QN(n1284) );
  SDFFX1 \fifo_reg[1][30]  ( .D(n1364), .SI(\fifo[1][29] ), .SE(test_se), 
        .CLK(n17), .Q(\fifo[1][30] ), .QN(n1285) );
  SDFFX1 \fifo_reg[1][29]  ( .D(n1365), .SI(\fifo[1][28] ), .SE(test_se), 
        .CLK(n17), .Q(\fifo[1][29] ), .QN(n1286) );
  SDFFX1 \fifo_reg[1][28]  ( .D(n1366), .SI(\fifo[1][27] ), .SE(test_se), 
        .CLK(n17), .Q(\fifo[1][28] ), .QN(n1287) );
  SDFFX1 \fifo_reg[1][27]  ( .D(n1367), .SI(\fifo[1][26] ), .SE(test_se), 
        .CLK(n17), .Q(\fifo[1][27] ), .QN(n1288) );
  SDFFX1 \fifo_reg[1][26]  ( .D(n1368), .SI(\fifo[1][25] ), .SE(test_se), 
        .CLK(n17), .Q(\fifo[1][26] ), .QN(n1289) );
  SDFFX1 \fifo_reg[1][25]  ( .D(n1369), .SI(\fifo[1][24] ), .SE(test_se), 
        .CLK(n17), .Q(\fifo[1][25] ), .QN(n1290) );
  SDFFX1 \fifo_reg[1][24]  ( .D(n1370), .SI(\fifo[1][23] ), .SE(test_se), 
        .CLK(n17), .Q(\fifo[1][24] ), .QN(n1291) );
  SDFFX1 \fifo_reg[1][23]  ( .D(n1371), .SI(\fifo[1][22] ), .SE(test_se), 
        .CLK(n17), .Q(\fifo[1][23] ), .QN(n1292) );
  SDFFX1 \fifo_reg[1][22]  ( .D(n1372), .SI(\fifo[1][21] ), .SE(test_se), 
        .CLK(n17), .Q(\fifo[1][22] ), .QN(n1293) );
  SDFFX1 \fifo_reg[1][21]  ( .D(n1373), .SI(\fifo[1][20] ), .SE(test_se), 
        .CLK(n17), .Q(\fifo[1][21] ), .QN(n1294) );
  SDFFX1 \fifo_reg[1][20]  ( .D(n1374), .SI(\fifo[1][19] ), .SE(test_se), 
        .CLK(n17), .Q(\fifo[1][20] ), .QN(n1295) );
  SDFFX1 \fifo_reg[1][19]  ( .D(n1375), .SI(\fifo[1][18] ), .SE(test_se), 
        .CLK(n17), .Q(\fifo[1][19] ), .QN(n1296) );
  SDFFX1 \fifo_reg[1][18]  ( .D(n1376), .SI(\fifo[1][17] ), .SE(test_se), 
        .CLK(n17), .Q(\fifo[1][18] ), .QN(n1297) );
  SDFFX1 \fifo_reg[1][17]  ( .D(n1377), .SI(\fifo[1][16] ), .SE(test_se), 
        .CLK(n16), .Q(\fifo[1][17] ), .QN(n1298) );
  SDFFX1 \fifo_reg[1][16]  ( .D(n1378), .SI(\fifo[1][15] ), .SE(test_se), 
        .CLK(n16), .Q(\fifo[1][16] ), .QN(n1299) );
  SDFFX1 \fifo_reg[1][15]  ( .D(n1379), .SI(\fifo[1][14] ), .SE(test_se), 
        .CLK(n16), .Q(\fifo[1][15] ), .QN(n1300) );
  SDFFX1 \fifo_reg[1][14]  ( .D(n1380), .SI(\fifo[1][13] ), .SE(test_se), 
        .CLK(n16), .Q(\fifo[1][14] ), .QN(n1301) );
  SDFFX1 \fifo_reg[1][13]  ( .D(n1381), .SI(\fifo[1][12] ), .SE(test_se), 
        .CLK(n16), .Q(\fifo[1][13] ), .QN(n1302) );
  SDFFX1 \fifo_reg[1][12]  ( .D(n1382), .SI(\fifo[1][11] ), .SE(test_se), 
        .CLK(n16), .Q(\fifo[1][12] ), .QN(n1303) );
  SDFFX1 \fifo_reg[1][11]  ( .D(n1383), .SI(\fifo[1][10] ), .SE(test_se), 
        .CLK(n16), .Q(\fifo[1][11] ), .QN(n1304) );
  SDFFX1 \fifo_reg[1][10]  ( .D(n1384), .SI(\fifo[1][9] ), .SE(test_se), .CLK(
        n16), .Q(\fifo[1][10] ), .QN(n1305) );
  SDFFX1 \fifo_reg[1][9]  ( .D(n1385), .SI(\fifo[1][8] ), .SE(test_se), .CLK(
        n16), .Q(\fifo[1][9] ), .QN(n1306) );
  SDFFX1 \fifo_reg[1][8]  ( .D(n1386), .SI(\fifo[1][7] ), .SE(test_se), .CLK(
        n16), .Q(\fifo[1][8] ), .QN(n1307) );
  SDFFX1 \fifo_reg[1][7]  ( .D(n1387), .SI(\fifo[1][6] ), .SE(test_se), .CLK(
        n16), .Q(\fifo[1][7] ), .QN(n1308) );
  SDFFX1 \fifo_reg[1][6]  ( .D(n1388), .SI(\fifo[1][5] ), .SE(test_se), .CLK(
        n16), .Q(\fifo[1][6] ), .QN(n1309) );
  SDFFX1 \fifo_reg[1][5]  ( .D(n1389), .SI(\fifo[1][4] ), .SE(test_se), .CLK(
        n16), .Q(\fifo[1][5] ), .QN(n1310) );
  SDFFX1 \fifo_reg[1][4]  ( .D(n1390), .SI(\fifo[1][3] ), .SE(test_se), .CLK(
        n16), .Q(\fifo[1][4] ), .QN(n1314) );
  SDFFX1 \fifo_reg[1][3]  ( .D(n1391), .SI(\fifo[1][2] ), .SE(test_se), .CLK(
        n15), .Q(\fifo[1][3] ), .QN(n1315) );
  SDFFX1 \fifo_reg[1][2]  ( .D(n1392), .SI(\fifo[1][1] ), .SE(test_se), .CLK(
        n15), .Q(\fifo[1][2] ), .QN(n1316) );
  SDFFX1 \fifo_reg[1][1]  ( .D(n1393), .SI(\fifo[1][0] ), .SE(test_se), .CLK(
        n15), .Q(\fifo[1][1] ), .QN(n1317) );
  SDFFX1 \fifo_reg[1][0]  ( .D(n1394), .SI(\fifo[0][31] ), .SE(test_se), .CLK(
        n15), .Q(\fifo[1][0] ), .QN(n1843) );
  SDFFX1 \fifo_reg[2][31]  ( .D(n1395), .SI(\fifo[2][30] ), .SE(test_se), 
        .CLK(n20), .Q(\fifo[2][31] ), .QN(n1849) );
  SDFFX1 \fifo_reg[2][30]  ( .D(n1396), .SI(\fifo[2][29] ), .SE(test_se), 
        .CLK(n20), .Q(\fifo[2][30] ), .QN(n1850) );
  SDFFX1 \fifo_reg[2][29]  ( .D(n1397), .SI(\fifo[2][28] ), .SE(test_se), 
        .CLK(n20), .Q(\fifo[2][29] ), .QN(n1851) );
  SDFFX1 \fifo_reg[2][28]  ( .D(n1398), .SI(\fifo[2][27] ), .SE(test_se), 
        .CLK(n20), .Q(\fifo[2][28] ), .QN(n1852) );
  SDFFX1 \fifo_reg[2][27]  ( .D(n1399), .SI(\fifo[2][26] ), .SE(test_se), 
        .CLK(n19), .Q(\fifo[2][27] ), .QN(n1853) );
  SDFFX1 \fifo_reg[2][26]  ( .D(n1400), .SI(\fifo[2][25] ), .SE(test_se), 
        .CLK(n19), .Q(\fifo[2][26] ), .QN(n1854) );
  SDFFX1 \fifo_reg[2][25]  ( .D(n1401), .SI(\fifo[2][24] ), .SE(test_se), 
        .CLK(n19), .Q(\fifo[2][25] ), .QN(n1855) );
  SDFFX1 \fifo_reg[2][24]  ( .D(n1402), .SI(\fifo[2][23] ), .SE(test_se), 
        .CLK(n19), .Q(\fifo[2][24] ), .QN(n1856) );
  SDFFX1 \fifo_reg[2][23]  ( .D(n1403), .SI(\fifo[2][22] ), .SE(test_se), 
        .CLK(n19), .Q(\fifo[2][23] ), .QN(n1857) );
  SDFFX1 \fifo_reg[2][22]  ( .D(n1404), .SI(\fifo[2][21] ), .SE(test_se), 
        .CLK(n19), .Q(\fifo[2][22] ), .QN(n1858) );
  SDFFX1 \fifo_reg[2][21]  ( .D(n1405), .SI(\fifo[2][20] ), .SE(test_se), 
        .CLK(n19), .Q(\fifo[2][21] ), .QN(n1859) );
  SDFFX1 \fifo_reg[2][20]  ( .D(n1406), .SI(\fifo[2][19] ), .SE(test_se), 
        .CLK(n19), .Q(\fifo[2][20] ), .QN(n1860) );
  SDFFX1 \fifo_reg[2][19]  ( .D(n1407), .SI(\fifo[2][18] ), .SE(test_se), 
        .CLK(n19), .Q(\fifo[2][19] ), .QN(n1861) );
  SDFFX1 \fifo_reg[2][18]  ( .D(n1408), .SI(\fifo[2][17] ), .SE(test_se), 
        .CLK(n19), .Q(\fifo[2][18] ), .QN(n1862) );
  SDFFX1 \fifo_reg[2][17]  ( .D(n1409), .SI(\fifo[2][16] ), .SE(test_se), 
        .CLK(n19), .Q(\fifo[2][17] ), .QN(n1863) );
  SDFFX1 \fifo_reg[2][16]  ( .D(n1410), .SI(\fifo[2][15] ), .SE(test_se), 
        .CLK(n19), .Q(\fifo[2][16] ), .QN(n1864) );
  SDFFX1 \fifo_reg[2][15]  ( .D(n1411), .SI(\fifo[2][14] ), .SE(test_se), 
        .CLK(n19), .Q(\fifo[2][15] ), .QN(n1865) );
  SDFFX1 \fifo_reg[2][14]  ( .D(n1412), .SI(\fifo[2][13] ), .SE(test_se), 
        .CLK(n19), .Q(\fifo[2][14] ), .QN(n1866) );
  SDFFX1 \fifo_reg[2][13]  ( .D(n1413), .SI(\fifo[2][12] ), .SE(test_se), 
        .CLK(n18), .Q(\fifo[2][13] ), .QN(n1867) );
  SDFFX1 \fifo_reg[2][12]  ( .D(n1414), .SI(\fifo[2][11] ), .SE(test_se), 
        .CLK(n18), .Q(\fifo[2][12] ), .QN(n1868) );
  SDFFX1 \fifo_reg[2][11]  ( .D(n1415), .SI(\fifo[2][10] ), .SE(test_se), 
        .CLK(n18), .Q(\fifo[2][11] ), .QN(n1869) );
  SDFFX1 \fifo_reg[2][10]  ( .D(n1416), .SI(\fifo[2][9] ), .SE(test_se), .CLK(
        n18), .Q(\fifo[2][10] ), .QN(n1870) );
  SDFFX1 \fifo_reg[2][9]  ( .D(n1417), .SI(\fifo[2][8] ), .SE(test_se), .CLK(
        n18), .Q(\fifo[2][9] ), .QN(n1871) );
  SDFFX1 \fifo_reg[2][8]  ( .D(n1418), .SI(\fifo[2][7] ), .SE(test_se), .CLK(
        n18), .Q(\fifo[2][8] ), .QN(n1872) );
  SDFFX1 \fifo_reg[2][7]  ( .D(n1419), .SI(\fifo[2][6] ), .SE(test_se), .CLK(
        n18), .Q(\fifo[2][7] ), .QN(n1873) );
  SDFFX1 \fifo_reg[2][6]  ( .D(n1420), .SI(\fifo[2][5] ), .SE(test_se), .CLK(
        n18), .Q(\fifo[2][6] ), .QN(n1874) );
  SDFFX1 \fifo_reg[2][5]  ( .D(n1421), .SI(\fifo[2][4] ), .SE(test_se), .CLK(
        n18), .Q(\fifo[2][5] ), .QN(n1875) );
  SDFFX1 \fifo_reg[2][4]  ( .D(n1422), .SI(\fifo[2][3] ), .SE(test_se), .CLK(
        n18), .Q(\fifo[2][4] ), .QN(n1876) );
  SDFFX1 \fifo_reg[2][3]  ( .D(n1423), .SI(\fifo[2][2] ), .SE(test_se), .CLK(
        n18), .Q(\fifo[2][3] ), .QN(n1877) );
  SDFFX1 \fifo_reg[2][2]  ( .D(n1424), .SI(\fifo[2][1] ), .SE(test_se), .CLK(
        n18), .Q(\fifo[2][2] ), .QN(n1878) );
  SDFFX1 \fifo_reg[2][1]  ( .D(n1425), .SI(\fifo[2][0] ), .SE(test_se), .CLK(
        n18), .Q(\fifo[2][1] ), .QN(n1879) );
  SDFFX1 \fifo_reg[2][0]  ( .D(n1426), .SI(\fifo[1][31] ), .SE(test_se), .CLK(
        n18), .Q(\fifo[2][0] ), .QN(n1880) );
  SDFFX1 \fifo_reg[3][31]  ( .D(n1427), .SI(\fifo[3][30] ), .SE(test_se), 
        .CLK(n22), .Q(\fifo[3][31] ), .QN(n1881) );
  SDFFX1 \fifo_reg[3][30]  ( .D(n1428), .SI(\fifo[3][29] ), .SE(test_se), 
        .CLK(n22), .Q(\fifo[3][30] ), .QN(n1882) );
  SDFFX1 \fifo_reg[3][29]  ( .D(n1429), .SI(\fifo[3][28] ), .SE(test_se), 
        .CLK(n22), .Q(\fifo[3][29] ), .QN(n1883) );
  SDFFX1 \fifo_reg[3][28]  ( .D(n1430), .SI(\fifo[3][27] ), .SE(test_se), 
        .CLK(n22), .Q(\fifo[3][28] ), .QN(n1884) );
  SDFFX1 \fifo_reg[3][27]  ( .D(n1431), .SI(\fifo[3][26] ), .SE(test_se), 
        .CLK(n22), .Q(\fifo[3][27] ), .QN(n1885) );
  SDFFX1 \fifo_reg[3][26]  ( .D(n1432), .SI(\fifo[3][25] ), .SE(test_se), 
        .CLK(n22), .Q(\fifo[3][26] ), .QN(n1886) );
  SDFFX1 \fifo_reg[3][25]  ( .D(n1433), .SI(\fifo[3][24] ), .SE(test_se), 
        .CLK(n22), .Q(\fifo[3][25] ), .QN(n1887) );
  SDFFX1 \fifo_reg[3][24]  ( .D(n1434), .SI(\fifo[3][23] ), .SE(test_se), 
        .CLK(n22), .Q(\fifo[3][24] ), .QN(n1888) );
  SDFFX1 \fifo_reg[3][23]  ( .D(n1435), .SI(\fifo[3][22] ), .SE(test_se), 
        .CLK(n22), .Q(\fifo[3][23] ), .QN(n1889) );
  SDFFX1 \fifo_reg[3][22]  ( .D(n1436), .SI(\fifo[3][21] ), .SE(test_se), 
        .CLK(n21), .Q(\fifo[3][22] ), .QN(n1890) );
  SDFFX1 \fifo_reg[3][21]  ( .D(n1437), .SI(\fifo[3][20] ), .SE(test_se), 
        .CLK(n21), .Q(\fifo[3][21] ), .QN(n1891) );
  SDFFX1 \fifo_reg[3][20]  ( .D(n1438), .SI(\fifo[3][19] ), .SE(test_se), 
        .CLK(n21), .Q(\fifo[3][20] ), .QN(n1892) );
  SDFFX1 \fifo_reg[3][19]  ( .D(n1439), .SI(\fifo[3][18] ), .SE(test_se), 
        .CLK(n21), .Q(\fifo[3][19] ), .QN(n1893) );
  SDFFX1 \fifo_reg[3][18]  ( .D(n1440), .SI(\fifo[3][17] ), .SE(test_se), 
        .CLK(n21), .Q(\fifo[3][18] ), .QN(n1894) );
  SDFFX1 \fifo_reg[3][17]  ( .D(n1441), .SI(\fifo[3][16] ), .SE(test_se), 
        .CLK(n21), .Q(\fifo[3][17] ), .QN(n1895) );
  SDFFX1 \fifo_reg[3][16]  ( .D(n1442), .SI(\fifo[3][15] ), .SE(test_se), 
        .CLK(n21), .Q(\fifo[3][16] ), .QN(n1896) );
  SDFFX1 \fifo_reg[3][15]  ( .D(n1443), .SI(\fifo[3][14] ), .SE(test_se), 
        .CLK(n21), .Q(\fifo[3][15] ), .QN(n1897) );
  SDFFX1 \fifo_reg[3][14]  ( .D(n1444), .SI(\fifo[3][13] ), .SE(test_se), 
        .CLK(n21), .Q(\fifo[3][14] ), .QN(n1898) );
  SDFFX1 \fifo_reg[3][13]  ( .D(n1445), .SI(\fifo[3][12] ), .SE(test_se), 
        .CLK(n21), .Q(\fifo[3][13] ), .QN(n1899) );
  SDFFX1 \fifo_reg[3][12]  ( .D(n1446), .SI(\fifo[3][11] ), .SE(test_se), 
        .CLK(n21), .Q(\fifo[3][12] ), .QN(n1900) );
  SDFFX1 \fifo_reg[3][11]  ( .D(n1447), .SI(\fifo[3][10] ), .SE(test_se), 
        .CLK(n21), .Q(\fifo[3][11] ), .QN(n1901) );
  SDFFX1 \fifo_reg[3][10]  ( .D(n1448), .SI(\fifo[3][9] ), .SE(test_se), .CLK(
        n21), .Q(\fifo[3][10] ), .QN(n1902) );
  SDFFX1 \fifo_reg[3][9]  ( .D(n1449), .SI(\fifo[3][8] ), .SE(test_se), .CLK(
        n21), .Q(\fifo[3][9] ), .QN(n1903) );
  SDFFX1 \fifo_reg[3][8]  ( .D(n1450), .SI(\fifo[3][7] ), .SE(test_se), .CLK(
        n20), .Q(\fifo[3][8] ), .QN(n1904) );
  SDFFX1 \fifo_reg[3][7]  ( .D(n1451), .SI(\fifo[3][6] ), .SE(test_se), .CLK(
        n20), .Q(\fifo[3][7] ), .QN(n1905) );
  SDFFX1 \fifo_reg[3][6]  ( .D(n1452), .SI(\fifo[3][5] ), .SE(test_se), .CLK(
        n20), .Q(\fifo[3][6] ), .QN(n1906) );
  SDFFX1 \fifo_reg[3][5]  ( .D(n1453), .SI(\fifo[3][4] ), .SE(test_se), .CLK(
        n20), .Q(\fifo[3][5] ), .QN(n1907) );
  SDFFX1 \fifo_reg[3][4]  ( .D(n1454), .SI(\fifo[3][3] ), .SE(test_se), .CLK(
        n20), .Q(\fifo[3][4] ), .QN(n1908) );
  SDFFX1 \fifo_reg[3][3]  ( .D(n1455), .SI(\fifo[3][2] ), .SE(test_se), .CLK(
        n20), .Q(\fifo[3][3] ), .QN(n1909) );
  SDFFX1 \fifo_reg[3][2]  ( .D(n1456), .SI(\fifo[3][1] ), .SE(test_se), .CLK(
        n20), .Q(\fifo[3][2] ), .QN(n1910) );
  SDFFX1 \fifo_reg[3][1]  ( .D(n1457), .SI(\fifo[3][0] ), .SE(test_se), .CLK(
        n20), .Q(\fifo[3][1] ), .QN(n1911) );
  SDFFX1 \fifo_reg[3][0]  ( .D(n1458), .SI(\fifo[2][31] ), .SE(test_se), .CLK(
        n20), .Q(\fifo[3][0] ), .QN(n1912) );
  SDFFX1 \fifo_reg[4][31]  ( .D(n1459), .SI(\fifo[4][30] ), .SE(test_se), 
        .CLK(n24), .Q(\fifo[4][31] ), .QN(n1913) );
  SDFFX1 \fifo_reg[4][30]  ( .D(n1460), .SI(\fifo[4][29] ), .SE(test_se), 
        .CLK(n24), .Q(\fifo[4][30] ), .QN(n1914) );
  SDFFX1 \fifo_reg[4][29]  ( .D(n1461), .SI(\fifo[4][28] ), .SE(test_se), 
        .CLK(n24), .Q(\fifo[4][29] ), .QN(n1915) );
  SDFFX1 \fifo_reg[4][28]  ( .D(n1462), .SI(\fifo[4][27] ), .SE(test_se), 
        .CLK(n24), .Q(\fifo[4][28] ), .QN(n1916) );
  SDFFX1 \fifo_reg[4][27]  ( .D(n1463), .SI(\fifo[4][26] ), .SE(test_se), 
        .CLK(n24), .Q(\fifo[4][27] ), .QN(n1917) );
  SDFFX1 \fifo_reg[4][26]  ( .D(n1464), .SI(\fifo[4][25] ), .SE(test_se), 
        .CLK(n24), .Q(\fifo[4][26] ), .QN(n1918) );
  SDFFX1 \fifo_reg[4][25]  ( .D(n1465), .SI(\fifo[4][24] ), .SE(test_se), 
        .CLK(n24), .Q(\fifo[4][25] ), .QN(n1919) );
  SDFFX1 \fifo_reg[4][24]  ( .D(n1466), .SI(\fifo[4][23] ), .SE(test_se), 
        .CLK(n24), .Q(\fifo[4][24] ), .QN(n1920) );
  SDFFX1 \fifo_reg[4][23]  ( .D(n1467), .SI(\fifo[4][22] ), .SE(test_se), 
        .CLK(n24), .Q(\fifo[4][23] ), .QN(n1921) );
  SDFFX1 \fifo_reg[4][22]  ( .D(n1468), .SI(\fifo[4][21] ), .SE(test_se), 
        .CLK(n24), .Q(\fifo[4][22] ), .QN(n1922) );
  SDFFX1 \fifo_reg[4][21]  ( .D(n1469), .SI(\fifo[4][20] ), .SE(test_se), 
        .CLK(n24), .Q(\fifo[4][21] ), .QN(n1923) );
  SDFFX1 \fifo_reg[4][20]  ( .D(n1470), .SI(\fifo[4][19] ), .SE(test_se), 
        .CLK(n24), .Q(\fifo[4][20] ), .QN(n1924) );
  SDFFX1 \fifo_reg[4][19]  ( .D(n1471), .SI(\fifo[4][18] ), .SE(test_se), 
        .CLK(n24), .Q(\fifo[4][19] ), .QN(n1925) );
  SDFFX1 \fifo_reg[4][18]  ( .D(n1472), .SI(\fifo[4][17] ), .SE(test_se), 
        .CLK(n23), .Q(\fifo[4][18] ), .QN(n1926) );
  SDFFX1 \fifo_reg[4][17]  ( .D(n1473), .SI(\fifo[4][16] ), .SE(test_se), 
        .CLK(n23), .Q(\fifo[4][17] ), .QN(n1927) );
  SDFFX1 \fifo_reg[4][16]  ( .D(n1474), .SI(\fifo[4][15] ), .SE(test_se), 
        .CLK(n23), .Q(\fifo[4][16] ), .QN(n1928) );
  SDFFX1 \fifo_reg[4][15]  ( .D(n1475), .SI(\fifo[4][14] ), .SE(test_se), 
        .CLK(n23), .Q(\fifo[4][15] ), .QN(n1929) );
  SDFFX1 \fifo_reg[4][14]  ( .D(n1476), .SI(\fifo[4][13] ), .SE(test_se), 
        .CLK(n23), .Q(\fifo[4][14] ), .QN(n1930) );
  SDFFX1 \fifo_reg[4][13]  ( .D(n1477), .SI(\fifo[4][12] ), .SE(test_se), 
        .CLK(n23), .Q(\fifo[4][13] ), .QN(n1931) );
  SDFFX1 \fifo_reg[4][12]  ( .D(n1478), .SI(\fifo[4][11] ), .SE(test_se), 
        .CLK(n23), .Q(\fifo[4][12] ), .QN(n1932) );
  SDFFX1 \fifo_reg[4][11]  ( .D(n1479), .SI(\fifo[4][10] ), .SE(test_se), 
        .CLK(n23), .Q(\fifo[4][11] ), .QN(n1933) );
  SDFFX1 \fifo_reg[4][10]  ( .D(n1480), .SI(\fifo[4][9] ), .SE(test_se), .CLK(
        n23), .Q(\fifo[4][10] ), .QN(n1934) );
  SDFFX1 \fifo_reg[4][9]  ( .D(n1481), .SI(\fifo[4][8] ), .SE(test_se), .CLK(
        n23), .Q(\fifo[4][9] ), .QN(n922) );
  SDFFX1 \fifo_reg[4][8]  ( .D(n1482), .SI(\fifo[4][7] ), .SE(test_se), .CLK(
        n23), .Q(\fifo[4][8] ), .QN(n923) );
  SDFFX1 \fifo_reg[4][7]  ( .D(n1483), .SI(\fifo[4][6] ), .SE(test_se), .CLK(
        n23), .Q(\fifo[4][7] ), .QN(n924) );
  SDFFX1 \fifo_reg[4][6]  ( .D(n1484), .SI(\fifo[4][5] ), .SE(test_se), .CLK(
        n23), .Q(\fifo[4][6] ), .QN(n925) );
  SDFFX1 \fifo_reg[4][5]  ( .D(n1485), .SI(\fifo[4][4] ), .SE(test_se), .CLK(
        n23), .Q(\fifo[4][5] ), .QN(n926) );
  SDFFX1 \fifo_reg[4][4]  ( .D(n1486), .SI(\fifo[4][3] ), .SE(test_se), .CLK(
        n22), .Q(\fifo[4][4] ), .QN(n927) );
  SDFFX1 \fifo_reg[4][3]  ( .D(n1487), .SI(\fifo[4][2] ), .SE(test_se), .CLK(
        n22), .Q(\fifo[4][3] ), .QN(n928) );
  SDFFX1 \fifo_reg[4][2]  ( .D(n1488), .SI(\fifo[4][1] ), .SE(test_se), .CLK(
        n22), .Q(\fifo[4][2] ), .QN(n929) );
  SDFFX1 \fifo_reg[4][1]  ( .D(n1489), .SI(\fifo[4][0] ), .SE(test_se), .CLK(
        n22), .Q(\fifo[4][1] ), .QN(n930) );
  SDFFX1 \fifo_reg[4][0]  ( .D(n1490), .SI(\fifo[3][31] ), .SE(test_se), .CLK(
        n22), .Q(\fifo[4][0] ), .QN(n931) );
  SDFFX1 \fifo_reg[5][31]  ( .D(n1491), .SI(\fifo[5][30] ), .SE(test_se), 
        .CLK(n8), .Q(\fifo[5][31] ), .QN(n932) );
  SDFFX1 \fifo_reg[5][30]  ( .D(n1492), .SI(\fifo[5][29] ), .SE(test_se), 
        .CLK(n7), .Q(\fifo[5][30] ), .QN(n933) );
  SDFFX1 \fifo_reg[5][29]  ( .D(n1493), .SI(\fifo[5][28] ), .SE(test_se), 
        .CLK(n7), .Q(\fifo[5][29] ), .QN(n934) );
  SDFFX1 \fifo_reg[5][28]  ( .D(n1494), .SI(\fifo[5][27] ), .SE(test_se), 
        .CLK(n7), .Q(\fifo[5][28] ), .QN(n935) );
  SDFFX1 \fifo_reg[5][27]  ( .D(n1495), .SI(\fifo[5][26] ), .SE(test_se), 
        .CLK(n7), .Q(\fifo[5][27] ), .QN(n936) );
  SDFFX1 \fifo_reg[5][26]  ( .D(n1496), .SI(\fifo[5][25] ), .SE(test_se), 
        .CLK(n7), .Q(\fifo[5][26] ), .QN(n937) );
  SDFFX1 \fifo_reg[5][25]  ( .D(n1497), .SI(\fifo[5][24] ), .SE(test_se), 
        .CLK(n8), .Q(\fifo[5][25] ), .QN(n938) );
  SDFFX1 \fifo_reg[5][24]  ( .D(n1498), .SI(\fifo[5][23] ), .SE(test_se), 
        .CLK(n7), .Q(\fifo[5][24] ), .QN(n939) );
  SDFFX1 \fifo_reg[5][23]  ( .D(n1499), .SI(\fifo[5][22] ), .SE(test_se), 
        .CLK(n7), .Q(\fifo[5][23] ), .QN(n940) );
  SDFFX1 \fifo_reg[5][22]  ( .D(n1500), .SI(\fifo[5][21] ), .SE(test_se), 
        .CLK(n6), .Q(\fifo[5][22] ), .QN(n941) );
  SDFFX1 \fifo_reg[5][21]  ( .D(n1501), .SI(\fifo[5][20] ), .SE(test_se), 
        .CLK(n7), .Q(\fifo[5][21] ), .QN(n942) );
  SDFFX1 \fifo_reg[5][20]  ( .D(n1502), .SI(\fifo[5][19] ), .SE(test_se), 
        .CLK(n6), .Q(\fifo[5][20] ), .QN(n943) );
  SDFFX1 \fifo_reg[5][19]  ( .D(n1503), .SI(\fifo[5][18] ), .SE(test_se), 
        .CLK(n7), .Q(\fifo[5][19] ), .QN(n944) );
  SDFFX1 \fifo_reg[5][18]  ( .D(n1504), .SI(\fifo[5][17] ), .SE(test_se), 
        .CLK(n6), .Q(\fifo[5][18] ), .QN(n945) );
  SDFFX1 \fifo_reg[5][17]  ( .D(n1505), .SI(\fifo[5][16] ), .SE(test_se), 
        .CLK(n7), .Q(\fifo[5][17] ), .QN(n946) );
  SDFFX1 \fifo_reg[5][16]  ( .D(n1506), .SI(\fifo[5][15] ), .SE(test_se), 
        .CLK(n6), .Q(\fifo[5][16] ), .QN(n947) );
  SDFFX1 \fifo_reg[5][15]  ( .D(n1507), .SI(\fifo[5][14] ), .SE(test_se), 
        .CLK(n6), .Q(\fifo[5][15] ), .QN(n948) );
  SDFFX1 \fifo_reg[5][14]  ( .D(n1508), .SI(\fifo[5][13] ), .SE(test_se), 
        .CLK(n6), .Q(\fifo[5][14] ), .QN(n949) );
  SDFFX1 \fifo_reg[5][13]  ( .D(n1509), .SI(\fifo[5][12] ), .SE(test_se), 
        .CLK(n7), .Q(\fifo[5][13] ), .QN(n950) );
  SDFFX1 \fifo_reg[5][12]  ( .D(n1510), .SI(\fifo[5][11] ), .SE(test_se), 
        .CLK(n6), .Q(\fifo[5][12] ), .QN(n951) );
  SDFFX1 \fifo_reg[5][11]  ( .D(n1511), .SI(\fifo[5][10] ), .SE(test_se), 
        .CLK(n6), .Q(\fifo[5][11] ), .QN(n952) );
  SDFFX1 \fifo_reg[5][10]  ( .D(n1512), .SI(\fifo[5][9] ), .SE(test_se), .CLK(
        n6), .Q(\fifo[5][10] ), .QN(n953) );
  SDFFX1 \fifo_reg[5][9]  ( .D(n1513), .SI(\fifo[5][8] ), .SE(test_se), .CLK(
        n6), .Q(\fifo[5][9] ), .QN(n954) );
  SDFFX1 \fifo_reg[5][8]  ( .D(n1514), .SI(\fifo[5][7] ), .SE(test_se), .CLK(
        n6), .Q(\fifo[5][8] ), .QN(n955) );
  SDFFX1 \fifo_reg[5][7]  ( .D(n1515), .SI(\fifo[5][6] ), .SE(test_se), .CLK(
        n7), .Q(\fifo[5][7] ), .QN(n956) );
  SDFFX1 \fifo_reg[5][6]  ( .D(n1516), .SI(\fifo[5][5] ), .SE(test_se), .CLK(
        n6), .Q(\fifo[5][6] ), .QN(n957) );
  SDFFX1 \fifo_reg[5][5]  ( .D(n1517), .SI(\fifo[5][4] ), .SE(test_se), .CLK(
        n25), .Q(\fifo[5][5] ), .QN(n958) );
  SDFFX1 \fifo_reg[5][4]  ( .D(n1518), .SI(\fifo[5][3] ), .SE(test_se), .CLK(
        n25), .Q(\fifo[5][4] ), .QN(n959) );
  SDFFX1 \fifo_reg[5][3]  ( .D(n1519), .SI(\fifo[5][2] ), .SE(test_se), .CLK(
        n25), .Q(\fifo[5][3] ), .QN(n960) );
  SDFFX1 \fifo_reg[5][2]  ( .D(n1520), .SI(\fifo[5][1] ), .SE(test_se), .CLK(
        n25), .Q(\fifo[5][2] ), .QN(n961) );
  SDFFX1 \fifo_reg[5][1]  ( .D(n1521), .SI(\fifo[5][0] ), .SE(test_se), .CLK(
        n25), .Q(\fifo[5][1] ), .QN(n962) );
  SDFFX1 \fifo_reg[5][0]  ( .D(n1522), .SI(\fifo[4][31] ), .SE(test_se), .CLK(
        n24), .Q(\fifo[5][0] ), .QN(n963) );
  SDFFX1 \fifo_reg[6][31]  ( .D(n1523), .SI(\fifo[6][30] ), .SE(test_se), 
        .CLK(n10), .Q(\fifo[6][31] ), .QN(n964) );
  SDFFX1 \fifo_reg[6][30]  ( .D(n1524), .SI(\fifo[6][29] ), .SE(test_se), 
        .CLK(n9), .Q(\fifo[6][30] ), .QN(n965) );
  SDFFX1 \fifo_reg[6][29]  ( .D(n1525), .SI(\fifo[6][28] ), .SE(test_se), 
        .CLK(n10), .Q(\fifo[6][29] ), .QN(n966) );
  SDFFX1 \fifo_reg[6][28]  ( .D(n1526), .SI(\fifo[6][27] ), .SE(test_se), 
        .CLK(n9), .Q(\fifo[6][28] ), .QN(n967) );
  SDFFX1 \fifo_reg[6][27]  ( .D(n1527), .SI(\fifo[6][26] ), .SE(test_se), 
        .CLK(n9), .Q(\fifo[6][27] ), .QN(n968) );
  SDFFX1 \fifo_reg[6][26]  ( .D(n1528), .SI(\fifo[6][25] ), .SE(test_se), 
        .CLK(n9), .Q(\fifo[6][26] ), .QN(n969) );
  SDFFX1 \fifo_reg[6][25]  ( .D(n1529), .SI(\fifo[6][24] ), .SE(test_se), 
        .CLK(n9), .Q(\fifo[6][25] ), .QN(n970) );
  SDFFX1 \fifo_reg[6][24]  ( .D(n1530), .SI(\fifo[6][23] ), .SE(test_se), 
        .CLK(n9), .Q(\fifo[6][24] ), .QN(n971) );
  SDFFX1 \fifo_reg[6][23]  ( .D(n1531), .SI(\fifo[6][22] ), .SE(test_se), 
        .CLK(n10), .Q(\fifo[6][23] ), .QN(n972) );
  SDFFX1 \fifo_reg[6][22]  ( .D(n1532), .SI(\fifo[6][21] ), .SE(test_se), 
        .CLK(n9), .Q(\fifo[6][22] ), .QN(n973) );
  SDFFX1 \fifo_reg[6][21]  ( .D(n1533), .SI(\fifo[6][20] ), .SE(test_se), 
        .CLK(n9), .Q(\fifo[6][21] ), .QN(n974) );
  SDFFX1 \fifo_reg[6][20]  ( .D(n1534), .SI(\fifo[6][19] ), .SE(test_se), 
        .CLK(n9), .Q(\fifo[6][20] ), .QN(n975) );
  SDFFX1 \fifo_reg[6][19]  ( .D(n1535), .SI(\fifo[6][18] ), .SE(test_se), 
        .CLK(n9), .Q(\fifo[6][19] ), .QN(n976) );
  SDFFX1 \fifo_reg[6][18]  ( .D(n1536), .SI(\fifo[6][17] ), .SE(test_se), 
        .CLK(n8), .Q(\fifo[6][18] ), .QN(n977) );
  SDFFX1 \fifo_reg[6][17]  ( .D(n1537), .SI(\fifo[6][16] ), .SE(test_se), 
        .CLK(n9), .Q(\fifo[6][17] ), .QN(n978) );
  SDFFX1 \fifo_reg[6][16]  ( .D(n1538), .SI(\fifo[6][15] ), .SE(test_se), 
        .CLK(n8), .Q(\fifo[6][16] ), .QN(n979) );
  SDFFX1 \fifo_reg[6][15]  ( .D(n1539), .SI(\fifo[6][14] ), .SE(test_se), 
        .CLK(n9), .Q(\fifo[6][15] ), .QN(n980) );
  SDFFX1 \fifo_reg[6][14]  ( .D(n1540), .SI(\fifo[6][13] ), .SE(test_se), 
        .CLK(n8), .Q(\fifo[6][14] ), .QN(n981) );
  SDFFX1 \fifo_reg[6][13]  ( .D(n1541), .SI(\fifo[6][12] ), .SE(test_se), 
        .CLK(n8), .Q(\fifo[6][13] ), .QN(n982) );
  SDFFX1 \fifo_reg[6][12]  ( .D(n1542), .SI(\fifo[6][11] ), .SE(test_se), 
        .CLK(n8), .Q(\fifo[6][12] ), .QN(n983) );
  SDFFX1 \fifo_reg[6][11]  ( .D(n1543), .SI(\fifo[6][10] ), .SE(test_se), 
        .CLK(n9), .Q(\fifo[6][11] ), .QN(n984) );
  SDFFX1 \fifo_reg[6][10]  ( .D(n1544), .SI(\fifo[6][9] ), .SE(test_se), .CLK(
        n8), .Q(\fifo[6][10] ), .QN(n985) );
  SDFFX1 \fifo_reg[6][9]  ( .D(n1545), .SI(\fifo[6][8] ), .SE(test_se), .CLK(
        n10), .Q(\fifo[6][9] ), .QN(n986) );
  SDFFX1 \fifo_reg[6][8]  ( .D(n1546), .SI(\fifo[6][7] ), .SE(test_se), .CLK(
        n8), .Q(\fifo[6][8] ), .QN(n987) );
  SDFFX1 \fifo_reg[6][7]  ( .D(n1547), .SI(\fifo[6][6] ), .SE(test_se), .CLK(
        n8), .Q(\fifo[6][7] ), .QN(n988) );
  SDFFX1 \fifo_reg[6][6]  ( .D(n1548), .SI(\fifo[6][5] ), .SE(test_se), .CLK(
        n8), .Q(\fifo[6][6] ), .QN(n989) );
  SDFFX1 \fifo_reg[6][5]  ( .D(n1549), .SI(\fifo[6][4] ), .SE(test_se), .CLK(
        n8), .Q(\fifo[6][5] ), .QN(n990) );
  SDFFX1 \fifo_reg[6][4]  ( .D(n1550), .SI(\fifo[6][3] ), .SE(test_se), .CLK(
        n7), .Q(\fifo[6][4] ), .QN(n991) );
  SDFFX1 \fifo_reg[6][3]  ( .D(n1551), .SI(\fifo[6][2] ), .SE(test_se), .CLK(
        n8), .Q(\fifo[6][3] ), .QN(n992) );
  SDFFX1 \fifo_reg[6][2]  ( .D(n1552), .SI(\fifo[6][1] ), .SE(test_se), .CLK(
        n9), .Q(\fifo[6][2] ), .QN(n993) );
  SDFFX1 \fifo_reg[6][1]  ( .D(n1553), .SI(\fifo[6][0] ), .SE(test_se), .CLK(
        n8), .Q(\fifo[6][1] ), .QN(n994) );
  SDFFX1 \fifo_reg[6][0]  ( .D(n1554), .SI(\fifo[5][31] ), .SE(test_se), .CLK(
        n7), .Q(\fifo[6][0] ), .QN(n995) );
  SDFFX1 \fifo_reg[7][31]  ( .D(n1555), .SI(\fifo[7][30] ), .SE(test_se), 
        .CLK(n12), .Q(\fifo[7][31] ), .QN(n996) );
  SDFFX1 \fifo_reg[7][30]  ( .D(n1556), .SI(\fifo[7][29] ), .SE(test_se), 
        .CLK(n12), .Q(\fifo[7][30] ), .QN(n997) );
  SDFFX1 \fifo_reg[7][29]  ( .D(n1557), .SI(\fifo[7][28] ), .SE(test_se), 
        .CLK(n12), .Q(\fifo[7][29] ), .QN(n998) );
  SDFFX1 \fifo_reg[7][28]  ( .D(n1558), .SI(\fifo[7][27] ), .SE(test_se), 
        .CLK(n12), .Q(\fifo[7][28] ), .QN(n999) );
  SDFFX1 \fifo_reg[7][27]  ( .D(n1559), .SI(\fifo[7][26] ), .SE(test_se), 
        .CLK(n12), .Q(\fifo[7][27] ), .QN(n1000) );
  SDFFX1 \fifo_reg[7][26]  ( .D(n1560), .SI(\fifo[7][25] ), .SE(test_se), 
        .CLK(n12), .Q(\fifo[7][26] ), .QN(n1001) );
  SDFFX1 \fifo_reg[7][25]  ( .D(n1561), .SI(\fifo[7][24] ), .SE(test_se), 
        .CLK(n12), .Q(\fifo[7][25] ), .QN(n1002) );
  SDFFX1 \fifo_reg[7][24]  ( .D(n1562), .SI(\fifo[7][23] ), .SE(test_se), 
        .CLK(n12), .Q(\fifo[7][24] ), .QN(n1003) );
  SDFFX1 \fifo_reg[7][23]  ( .D(n1563), .SI(\fifo[7][22] ), .SE(test_se), 
        .CLK(n11), .Q(\fifo[7][23] ), .QN(n1004) );
  SDFFX1 \fifo_reg[7][22]  ( .D(n1564), .SI(\fifo[7][21] ), .SE(test_se), 
        .CLK(n11), .Q(\fifo[7][22] ), .QN(n1005) );
  SDFFX1 \fifo_reg[7][21]  ( .D(n1565), .SI(\fifo[7][20] ), .SE(test_se), 
        .CLK(n11), .Q(\fifo[7][21] ), .QN(n1006) );
  SDFFX1 \fifo_reg[7][20]  ( .D(n1566), .SI(\fifo[7][19] ), .SE(test_se), 
        .CLK(n11), .Q(\fifo[7][20] ), .QN(n1007) );
  SDFFX1 \fifo_reg[7][19]  ( .D(n1567), .SI(\fifo[7][18] ), .SE(test_se), 
        .CLK(n11), .Q(\fifo[7][19] ), .QN(n1008) );
  SDFFX1 \fifo_reg[7][18]  ( .D(n1568), .SI(\fifo[7][17] ), .SE(test_se), 
        .CLK(n11), .Q(\fifo[7][18] ), .QN(n1009) );
  SDFFX1 \fifo_reg[7][17]  ( .D(n1569), .SI(\fifo[7][16] ), .SE(test_se), 
        .CLK(n11), .Q(\fifo[7][17] ), .QN(n1010) );
  SDFFX1 \fifo_reg[7][16]  ( .D(n1570), .SI(\fifo[7][15] ), .SE(test_se), 
        .CLK(n11), .Q(\fifo[7][16] ), .QN(n1011) );
  SDFFX1 \fifo_reg[7][15]  ( .D(n1571), .SI(\fifo[7][14] ), .SE(test_se), 
        .CLK(n11), .Q(\fifo[7][15] ), .QN(n1012) );
  SDFFX1 \fifo_reg[7][14]  ( .D(n1572), .SI(\fifo[7][13] ), .SE(test_se), 
        .CLK(n11), .Q(\fifo[7][14] ), .QN(n1013) );
  SDFFX1 \fifo_reg[7][13]  ( .D(n1573), .SI(\fifo[7][12] ), .SE(test_se), 
        .CLK(n11), .Q(\fifo[7][13] ), .QN(n1014) );
  SDFFX1 \fifo_reg[7][12]  ( .D(n1574), .SI(\fifo[7][11] ), .SE(test_se), 
        .CLK(n11), .Q(\fifo[7][12] ), .QN(n1015) );
  SDFFX1 \fifo_reg[7][11]  ( .D(n1575), .SI(\fifo[7][10] ), .SE(test_se), 
        .CLK(n11), .Q(\fifo[7][11] ), .QN(n1016) );
  SDFFX1 \fifo_reg[7][10]  ( .D(n1576), .SI(\fifo[7][9] ), .SE(test_se), .CLK(
        n11), .Q(\fifo[7][10] ), .QN(n1017) );
  SDFFX1 \fifo_reg[7][9]  ( .D(n1577), .SI(\fifo[7][8] ), .SE(test_se), .CLK(
        n10), .Q(\fifo[7][9] ), .QN(n1018) );
  SDFFX1 \fifo_reg[7][8]  ( .D(n1578), .SI(\fifo[7][7] ), .SE(test_se), .CLK(
        n10), .Q(\fifo[7][8] ), .QN(n1019) );
  SDFFX1 \fifo_reg[7][7]  ( .D(n1579), .SI(\fifo[7][6] ), .SE(test_se), .CLK(
        n10), .Q(\fifo[7][7] ), .QN(n1020) );
  SDFFX1 \fifo_reg[7][6]  ( .D(n1580), .SI(\fifo[7][5] ), .SE(test_se), .CLK(
        n10), .Q(\fifo[7][6] ), .QN(n1021) );
  SDFFX1 \fifo_reg[7][5]  ( .D(n1581), .SI(\fifo[7][4] ), .SE(test_se), .CLK(
        n10), .Q(\fifo[7][5] ), .QN(n1022) );
  SDFFX1 \fifo_reg[7][4]  ( .D(n1582), .SI(\fifo[7][3] ), .SE(test_se), .CLK(
        n10), .Q(\fifo[7][4] ), .QN(n1023) );
  SDFFX1 \fifo_reg[7][3]  ( .D(n1583), .SI(\fifo[7][2] ), .SE(test_se), .CLK(
        n10), .Q(\fifo[7][3] ), .QN(n1024) );
  SDFFX1 \fifo_reg[7][2]  ( .D(n1584), .SI(\fifo[7][1] ), .SE(test_se), .CLK(
        n10), .Q(\fifo[7][2] ), .QN(n1025) );
  SDFFX1 \fifo_reg[7][1]  ( .D(n1585), .SI(\fifo[7][0] ), .SE(test_se), .CLK(
        n10), .Q(\fifo[7][1] ), .QN(n1026) );
  SDFFX1 \fifo_reg[7][0]  ( .D(n1586), .SI(\fifo[6][31] ), .SE(test_se), .CLK(
        n10), .Q(\fifo[7][0] ), .QN(n1027) );
  SDFFX1 \fifo_reg[8][31]  ( .D(n1587), .SI(\fifo[8][30] ), .SE(test_se), 
        .CLK(n14), .Q(\fifo[8][31] ), .QN(n1028) );
  SDFFX1 \fifo_reg[8][30]  ( .D(n1588), .SI(\fifo[8][29] ), .SE(test_se), 
        .CLK(n14), .Q(\fifo[8][30] ), .QN(n1029) );
  SDFFX1 \fifo_reg[8][29]  ( .D(n1589), .SI(\fifo[8][28] ), .SE(test_se), 
        .CLK(n14), .Q(\fifo[8][29] ), .QN(n1030) );
  SDFFX1 \fifo_reg[8][28]  ( .D(n1590), .SI(\fifo[8][27] ), .SE(test_se), 
        .CLK(n14), .Q(\fifo[8][28] ), .QN(n1031) );
  SDFFX1 \fifo_reg[8][27]  ( .D(n1591), .SI(\fifo[8][26] ), .SE(test_se), 
        .CLK(n14), .Q(\fifo[8][27] ), .QN(n1032) );
  SDFFX1 \fifo_reg[8][26]  ( .D(n1592), .SI(\fifo[8][25] ), .SE(test_se), 
        .CLK(n14), .Q(\fifo[8][26] ), .QN(n1033) );
  SDFFX1 \fifo_reg[8][25]  ( .D(n1593), .SI(\fifo[8][24] ), .SE(test_se), 
        .CLK(n14), .Q(\fifo[8][25] ), .QN(n1034) );
  SDFFX1 \fifo_reg[8][24]  ( .D(n1594), .SI(\fifo[8][23] ), .SE(test_se), 
        .CLK(n14), .Q(\fifo[8][24] ), .QN(n1035) );
  SDFFX1 \fifo_reg[8][23]  ( .D(n1595), .SI(\fifo[8][22] ), .SE(test_se), 
        .CLK(n14), .Q(\fifo[8][23] ), .QN(n1036) );
  SDFFX1 \fifo_reg[8][22]  ( .D(n1596), .SI(\fifo[8][21] ), .SE(test_se), 
        .CLK(n14), .Q(\fifo[8][22] ), .QN(n1037) );
  SDFFX1 \fifo_reg[8][21]  ( .D(n1597), .SI(\fifo[8][20] ), .SE(test_se), 
        .CLK(n14), .Q(\fifo[8][21] ), .QN(n1038) );
  SDFFX1 \fifo_reg[8][20]  ( .D(n1598), .SI(\fifo[8][19] ), .SE(test_se), 
        .CLK(n14), .Q(\fifo[8][20] ), .QN(n1039) );
  SDFFX1 \fifo_reg[8][19]  ( .D(n1599), .SI(\fifo[8][18] ), .SE(test_se), 
        .CLK(n13), .Q(\fifo[8][19] ), .QN(n1040) );
  SDFFX1 \fifo_reg[8][18]  ( .D(n1600), .SI(\fifo[8][17] ), .SE(test_se), 
        .CLK(n13), .Q(\fifo[8][18] ), .QN(n1041) );
  SDFFX1 \fifo_reg[8][17]  ( .D(n1601), .SI(\fifo[8][16] ), .SE(test_se), 
        .CLK(n13), .Q(\fifo[8][17] ), .QN(n1042) );
  SDFFX1 \fifo_reg[8][16]  ( .D(n1602), .SI(\fifo[8][15] ), .SE(test_se), 
        .CLK(n13), .Q(\fifo[8][16] ), .QN(n1043) );
  SDFFX1 \fifo_reg[8][15]  ( .D(n1603), .SI(\fifo[8][14] ), .SE(test_se), 
        .CLK(n13), .Q(\fifo[8][15] ), .QN(n1044) );
  SDFFX1 \fifo_reg[8][14]  ( .D(n1604), .SI(\fifo[8][13] ), .SE(test_se), 
        .CLK(n13), .Q(\fifo[8][14] ), .QN(n1045) );
  SDFFX1 \fifo_reg[8][13]  ( .D(n1605), .SI(\fifo[8][12] ), .SE(test_se), 
        .CLK(n13), .Q(\fifo[8][13] ), .QN(n1046) );
  SDFFX1 \fifo_reg[8][12]  ( .D(n1606), .SI(\fifo[8][11] ), .SE(test_se), 
        .CLK(n13), .Q(\fifo[8][12] ), .QN(n1047) );
  SDFFX1 \fifo_reg[8][11]  ( .D(n1607), .SI(\fifo[8][10] ), .SE(test_se), 
        .CLK(n13), .Q(\fifo[8][11] ), .QN(n1048) );
  SDFFX1 \fifo_reg[8][10]  ( .D(n1608), .SI(\fifo[8][9] ), .SE(test_se), .CLK(
        n13), .Q(\fifo[8][10] ), .QN(n1049) );
  SDFFX1 \fifo_reg[8][9]  ( .D(n1609), .SI(\fifo[8][8] ), .SE(test_se), .CLK(
        n13), .Q(\fifo[8][9] ), .QN(n1050) );
  SDFFX1 \fifo_reg[8][8]  ( .D(n1610), .SI(\fifo[8][7] ), .SE(test_se), .CLK(
        n13), .Q(\fifo[8][8] ), .QN(n1051) );
  SDFFX1 \fifo_reg[8][7]  ( .D(n1611), .SI(\fifo[8][6] ), .SE(test_se), .CLK(
        n13), .Q(\fifo[8][7] ), .QN(n1052) );
  SDFFX1 \fifo_reg[8][6]  ( .D(n1612), .SI(\fifo[8][5] ), .SE(test_se), .CLK(
        n13), .Q(\fifo[8][6] ), .QN(n1053) );
  SDFFX1 \fifo_reg[8][5]  ( .D(n1613), .SI(\fifo[8][4] ), .SE(test_se), .CLK(
        n12), .Q(\fifo[8][5] ), .QN(n1054) );
  SDFFX1 \fifo_reg[8][4]  ( .D(n1614), .SI(\fifo[8][3] ), .SE(test_se), .CLK(
        n12), .Q(\fifo[8][4] ), .QN(n1055) );
  SDFFX1 \fifo_reg[8][3]  ( .D(n1615), .SI(\fifo[8][2] ), .SE(test_se), .CLK(
        n12), .Q(\fifo[8][3] ), .QN(n1056) );
  SDFFX1 \fifo_reg[8][2]  ( .D(n1616), .SI(\fifo[8][1] ), .SE(test_se), .CLK(
        n12), .Q(\fifo[8][2] ), .QN(n1057) );
  SDFFX1 \fifo_reg[8][1]  ( .D(n1617), .SI(\fifo[8][0] ), .SE(test_se), .CLK(
        n12), .Q(\fifo[8][1] ), .QN(n1058) );
  SDFFX1 \fifo_reg[8][0]  ( .D(n1618), .SI(\fifo[7][31] ), .SE(test_se), .CLK(
        n12), .Q(\fifo[8][0] ), .QN(n1059) );
  SDFFX1 \fifo_reg[9][31]  ( .D(n1619), .SI(\fifo[9][30] ), .SE(test_se), 
        .CLK(n36), .Q(\fifo[9][31] ), .QN(n1060) );
  SDFFX1 \fifo_reg[9][30]  ( .D(n1620), .SI(\fifo[9][29] ), .SE(test_se), 
        .CLK(n36), .Q(\fifo[9][30] ), .QN(n1061) );
  SDFFX1 \fifo_reg[9][29]  ( .D(n1621), .SI(\fifo[9][28] ), .SE(test_se), 
        .CLK(n36), .Q(\fifo[9][29] ), .QN(n1062) );
  SDFFX1 \fifo_reg[9][28]  ( .D(n1622), .SI(\fifo[9][27] ), .SE(test_se), 
        .CLK(n36), .Q(\fifo[9][28] ), .QN(n1063) );
  SDFFX1 \fifo_reg[9][27]  ( .D(n1623), .SI(\fifo[9][26] ), .SE(test_se), 
        .CLK(n36), .Q(\fifo[9][27] ), .QN(n1064) );
  SDFFX1 \fifo_reg[9][26]  ( .D(n1624), .SI(\fifo[9][25] ), .SE(test_se), 
        .CLK(n36), .Q(\fifo[9][26] ), .QN(n1065) );
  SDFFX1 \fifo_reg[9][25]  ( .D(n1625), .SI(\fifo[9][24] ), .SE(test_se), 
        .CLK(n36), .Q(\fifo[9][25] ), .QN(n1066) );
  SDFFX1 \fifo_reg[9][24]  ( .D(n1626), .SI(\fifo[9][23] ), .SE(test_se), 
        .CLK(n35), .Q(\fifo[9][24] ), .QN(n1067) );
  SDFFX1 \fifo_reg[9][23]  ( .D(n1627), .SI(\fifo[9][22] ), .SE(test_se), 
        .CLK(n35), .Q(\fifo[9][23] ), .QN(n1068) );
  SDFFX1 \fifo_reg[9][22]  ( .D(n1628), .SI(\fifo[9][21] ), .SE(test_se), 
        .CLK(n35), .Q(\fifo[9][22] ), .QN(n1069) );
  SDFFX1 \fifo_reg[9][21]  ( .D(n1629), .SI(\fifo[9][20] ), .SE(test_se), 
        .CLK(n35), .Q(\fifo[9][21] ), .QN(n1070) );
  SDFFX1 \fifo_reg[9][20]  ( .D(n1630), .SI(\fifo[9][19] ), .SE(test_se), 
        .CLK(n35), .Q(\fifo[9][20] ), .QN(n1071) );
  SDFFX1 \fifo_reg[9][19]  ( .D(n1631), .SI(\fifo[9][18] ), .SE(test_se), 
        .CLK(n35), .Q(\fifo[9][19] ), .QN(n1072) );
  SDFFX1 \fifo_reg[9][18]  ( .D(n1632), .SI(\fifo[9][17] ), .SE(test_se), 
        .CLK(n35), .Q(\fifo[9][18] ), .QN(n1073) );
  SDFFX1 \fifo_reg[9][17]  ( .D(n1633), .SI(\fifo[9][16] ), .SE(test_se), 
        .CLK(n35), .Q(\fifo[9][17] ), .QN(n1074) );
  SDFFX1 \fifo_reg[9][16]  ( .D(n1634), .SI(\fifo[9][15] ), .SE(test_se), 
        .CLK(n35), .Q(\fifo[9][16] ), .QN(n1075) );
  SDFFX1 \fifo_reg[9][15]  ( .D(n1635), .SI(\fifo[9][14] ), .SE(test_se), 
        .CLK(n35), .Q(\fifo[9][15] ), .QN(n1076) );
  SDFFX1 \fifo_reg[9][14]  ( .D(n1636), .SI(\fifo[9][13] ), .SE(test_se), 
        .CLK(n35), .Q(\fifo[9][14] ), .QN(n1077) );
  SDFFX1 \fifo_reg[9][13]  ( .D(n1637), .SI(\fifo[9][12] ), .SE(test_se), 
        .CLK(n35), .Q(\fifo[9][13] ), .QN(n1078) );
  SDFFX1 \fifo_reg[9][12]  ( .D(n1638), .SI(\fifo[9][11] ), .SE(test_se), 
        .CLK(n40), .Q(\fifo[9][12] ), .QN(n1079) );
  SDFFX1 \fifo_reg[9][11]  ( .D(n1639), .SI(\fifo[9][10] ), .SE(test_se), 
        .CLK(n15), .Q(\fifo[9][11] ), .QN(n1080) );
  SDFFX1 \fifo_reg[9][10]  ( .D(n1640), .SI(\fifo[9][9] ), .SE(test_se), .CLK(
        n15), .Q(\fifo[9][10] ), .QN(n1081) );
  SDFFX1 \fifo_reg[9][9]  ( .D(n1641), .SI(\fifo[9][8] ), .SE(test_se), .CLK(
        n15), .Q(\fifo[9][9] ), .QN(n1082) );
  SDFFX1 \fifo_reg[9][8]  ( .D(n1642), .SI(\fifo[9][7] ), .SE(test_se), .CLK(
        n15), .Q(\fifo[9][8] ), .QN(n1083) );
  SDFFX1 \fifo_reg[9][7]  ( .D(n1643), .SI(\fifo[9][6] ), .SE(test_se), .CLK(
        n15), .Q(\fifo[9][7] ), .QN(n1084) );
  SDFFX1 \fifo_reg[9][6]  ( .D(n1644), .SI(\fifo[9][5] ), .SE(test_se), .CLK(
        n15), .Q(\fifo[9][6] ), .QN(n1085) );
  SDFFX1 \fifo_reg[9][5]  ( .D(n1645), .SI(\fifo[9][4] ), .SE(test_se), .CLK(
        n15), .Q(\fifo[9][5] ), .QN(n1086) );
  SDFFX1 \fifo_reg[9][4]  ( .D(n1646), .SI(\fifo[9][3] ), .SE(test_se), .CLK(
        n15), .Q(\fifo[9][4] ), .QN(n1087) );
  SDFFX1 \fifo_reg[9][3]  ( .D(n1647), .SI(\fifo[9][2] ), .SE(test_se), .CLK(
        n15), .Q(\fifo[9][3] ), .QN(n1088) );
  SDFFX1 \fifo_reg[9][2]  ( .D(n1648), .SI(\fifo[9][1] ), .SE(test_se), .CLK(
        n15), .Q(\fifo[9][2] ), .QN(n1089) );
  SDFFX1 \fifo_reg[9][1]  ( .D(n1649), .SI(\fifo[9][0] ), .SE(test_se), .CLK(
        n14), .Q(\fifo[9][1] ), .QN(n1090) );
  SDFFX1 \fifo_reg[9][0]  ( .D(n1650), .SI(\fifo[8][31] ), .SE(test_se), .CLK(
        n14), .Q(\fifo[9][0] ), .QN(n1091) );
  SDFFX1 \fifo_reg[10][31]  ( .D(n1651), .SI(\fifo[10][30] ), .SE(test_se), 
        .CLK(n38), .Q(\fifo[10][31] ), .QN(n1092) );
  SDFFX1 \fifo_reg[10][30]  ( .D(n1652), .SI(\fifo[10][29] ), .SE(test_se), 
        .CLK(n38), .Q(\fifo[10][30] ), .QN(n1093) );
  SDFFX1 \fifo_reg[10][29]  ( .D(n1653), .SI(\fifo[10][28] ), .SE(test_se), 
        .CLK(n38), .Q(\fifo[10][29] ), .QN(n1094) );
  SDFFX1 \fifo_reg[10][28]  ( .D(n1654), .SI(\fifo[10][27] ), .SE(test_se), 
        .CLK(n38), .Q(\fifo[10][28] ), .QN(n1095) );
  SDFFX1 \fifo_reg[10][27]  ( .D(n1655), .SI(\fifo[10][26] ), .SE(test_se), 
        .CLK(n38), .Q(\fifo[10][27] ), .QN(n1096) );
  SDFFX1 \fifo_reg[10][26]  ( .D(n1656), .SI(\fifo[10][25] ), .SE(test_se), 
        .CLK(n38), .Q(\fifo[10][26] ), .QN(n1097) );
  SDFFX1 \fifo_reg[10][25]  ( .D(n1657), .SI(\fifo[10][24] ), .SE(test_se), 
        .CLK(n38), .Q(\fifo[10][25] ), .QN(n1098) );
  SDFFX1 \fifo_reg[10][24]  ( .D(n1658), .SI(\fifo[10][23] ), .SE(test_se), 
        .CLK(n38), .Q(\fifo[10][24] ), .QN(n1099) );
  SDFFX1 \fifo_reg[10][23]  ( .D(n1659), .SI(\fifo[10][22] ), .SE(test_se), 
        .CLK(n38), .Q(\fifo[10][23] ), .QN(n1100) );
  SDFFX1 \fifo_reg[10][22]  ( .D(n1660), .SI(\fifo[10][21] ), .SE(test_se), 
        .CLK(n38), .Q(\fifo[10][22] ), .QN(n1101) );
  SDFFX1 \fifo_reg[10][21]  ( .D(n1661), .SI(\fifo[10][20] ), .SE(test_se), 
        .CLK(n38), .Q(\fifo[10][21] ), .QN(n1102) );
  SDFFX1 \fifo_reg[10][20]  ( .D(n1662), .SI(\fifo[10][19] ), .SE(test_se), 
        .CLK(n37), .Q(\fifo[10][20] ), .QN(n1103) );
  SDFFX1 \fifo_reg[10][19]  ( .D(n1663), .SI(\fifo[10][18] ), .SE(test_se), 
        .CLK(n37), .Q(\fifo[10][19] ), .QN(n1104) );
  SDFFX1 \fifo_reg[10][18]  ( .D(n1664), .SI(\fifo[10][17] ), .SE(test_se), 
        .CLK(n37), .Q(\fifo[10][18] ), .QN(n1105) );
  SDFFX1 \fifo_reg[10][17]  ( .D(n1665), .SI(\fifo[10][16] ), .SE(test_se), 
        .CLK(n37), .Q(\fifo[10][17] ), .QN(n1106) );
  SDFFX1 \fifo_reg[10][16]  ( .D(n1666), .SI(\fifo[10][15] ), .SE(test_se), 
        .CLK(n37), .Q(\fifo[10][16] ), .QN(n1107) );
  SDFFX1 \fifo_reg[10][15]  ( .D(n1667), .SI(\fifo[10][14] ), .SE(test_se), 
        .CLK(n37), .Q(\fifo[10][15] ), .QN(n1108) );
  SDFFX1 \fifo_reg[10][14]  ( .D(n1668), .SI(\fifo[10][13] ), .SE(test_se), 
        .CLK(n37), .Q(\fifo[10][14] ), .QN(n1109) );
  SDFFX1 \fifo_reg[10][13]  ( .D(n1669), .SI(\fifo[10][12] ), .SE(test_se), 
        .CLK(n37), .Q(\fifo[10][13] ), .QN(n1110) );
  SDFFX1 \fifo_reg[10][12]  ( .D(n1670), .SI(\fifo[10][11] ), .SE(test_se), 
        .CLK(n37), .Q(\fifo[10][12] ), .QN(n1111) );
  SDFFX1 \fifo_reg[10][11]  ( .D(n1671), .SI(\fifo[10][10] ), .SE(test_se), 
        .CLK(n37), .Q(\fifo[10][11] ), .QN(n1112) );
  SDFFX1 \fifo_reg[10][10]  ( .D(n1672), .SI(\fifo[10][9] ), .SE(test_se), 
        .CLK(n37), .Q(\fifo[10][10] ), .QN(n1113) );
  SDFFX1 \fifo_reg[10][9]  ( .D(n1673), .SI(\fifo[10][8] ), .SE(test_se), 
        .CLK(n37), .Q(\fifo[10][9] ), .QN(n1114) );
  SDFFX1 \fifo_reg[10][8]  ( .D(n1674), .SI(\fifo[10][7] ), .SE(test_se), 
        .CLK(n37), .Q(\fifo[10][8] ), .QN(n1115) );
  SDFFX1 \fifo_reg[10][7]  ( .D(n1675), .SI(\fifo[10][6] ), .SE(test_se), 
        .CLK(n37), .Q(\fifo[10][7] ), .QN(n1116) );
  SDFFX1 \fifo_reg[10][6]  ( .D(n1676), .SI(\fifo[10][5] ), .SE(test_se), 
        .CLK(n36), .Q(\fifo[10][6] ), .QN(n1117) );
  SDFFX1 \fifo_reg[10][5]  ( .D(n1677), .SI(\fifo[10][4] ), .SE(test_se), 
        .CLK(n36), .Q(\fifo[10][5] ), .QN(n1118) );
  SDFFX1 \fifo_reg[10][4]  ( .D(n1678), .SI(\fifo[10][3] ), .SE(test_se), 
        .CLK(n36), .Q(\fifo[10][4] ), .QN(n1119) );
  SDFFX1 \fifo_reg[10][3]  ( .D(n1679), .SI(\fifo[10][2] ), .SE(test_se), 
        .CLK(n36), .Q(\fifo[10][3] ), .QN(n1120) );
  SDFFX1 \fifo_reg[10][2]  ( .D(n1680), .SI(\fifo[10][1] ), .SE(test_se), 
        .CLK(n36), .Q(\fifo[10][2] ), .QN(n1121) );
  SDFFX1 \fifo_reg[10][1]  ( .D(n1681), .SI(\fifo[10][0] ), .SE(test_se), 
        .CLK(n36), .Q(\fifo[10][1] ), .QN(n1122) );
  SDFFX1 \fifo_reg[10][0]  ( .D(n1682), .SI(\fifo[9][31] ), .SE(test_se), 
        .CLK(n36), .Q(\fifo[10][0] ), .QN(n1123) );
  SDFFX1 \fifo_reg[11][31]  ( .D(n1683), .SI(\fifo[11][30] ), .SE(test_se), 
        .CLK(n41), .Q(\fifo[11][31] ), .QN(n1124) );
  SDFFX1 \fifo_reg[11][30]  ( .D(n1684), .SI(\fifo[11][29] ), .SE(test_se), 
        .CLK(n41), .Q(\fifo[11][30] ), .QN(n1125) );
  SDFFX1 \fifo_reg[11][29]  ( .D(n1685), .SI(\fifo[11][28] ), .SE(test_se), 
        .CLK(n40), .Q(\fifo[11][29] ), .QN(n1126) );
  SDFFX1 \fifo_reg[11][28]  ( .D(n1686), .SI(\fifo[11][27] ), .SE(test_se), 
        .CLK(n40), .Q(\fifo[11][28] ), .QN(n1127) );
  SDFFX1 \fifo_reg[11][27]  ( .D(n1687), .SI(\fifo[11][26] ), .SE(test_se), 
        .CLK(n40), .Q(\fifo[11][27] ), .QN(n1128) );
  SDFFX1 \fifo_reg[11][26]  ( .D(n1688), .SI(\fifo[11][25] ), .SE(test_se), 
        .CLK(n40), .Q(\fifo[11][26] ), .QN(n1129) );
  SDFFX1 \fifo_reg[11][25]  ( .D(n1689), .SI(\fifo[11][24] ), .SE(test_se), 
        .CLK(n40), .Q(\fifo[11][25] ), .QN(n1130) );
  SDFFX1 \fifo_reg[11][24]  ( .D(n1690), .SI(\fifo[11][23] ), .SE(test_se), 
        .CLK(n40), .Q(\fifo[11][24] ), .QN(n1131) );
  SDFFX1 \fifo_reg[11][23]  ( .D(n1691), .SI(\fifo[11][22] ), .SE(test_se), 
        .CLK(n40), .Q(\fifo[11][23] ), .QN(n1132) );
  SDFFX1 \fifo_reg[11][22]  ( .D(n1692), .SI(\fifo[11][21] ), .SE(test_se), 
        .CLK(n40), .Q(\fifo[11][22] ), .QN(n1133) );
  SDFFX1 \fifo_reg[11][21]  ( .D(n1693), .SI(\fifo[11][20] ), .SE(test_se), 
        .CLK(n40), .Q(\fifo[11][21] ), .QN(n1134) );
  SDFFX1 \fifo_reg[11][20]  ( .D(n1694), .SI(\fifo[11][19] ), .SE(test_se), 
        .CLK(n40), .Q(\fifo[11][20] ), .QN(n1135) );
  SDFFX1 \fifo_reg[11][19]  ( .D(n1695), .SI(\fifo[11][18] ), .SE(test_se), 
        .CLK(n40), .Q(\fifo[11][19] ), .QN(n1136) );
  SDFFX1 \fifo_reg[11][18]  ( .D(n1696), .SI(\fifo[11][17] ), .SE(test_se), 
        .CLK(n40), .Q(\fifo[11][18] ), .QN(n1137) );
  SDFFX1 \fifo_reg[11][17]  ( .D(n1697), .SI(\fifo[11][16] ), .SE(test_se), 
        .CLK(n40), .Q(\fifo[11][17] ), .QN(n1138) );
  SDFFX1 \fifo_reg[11][16]  ( .D(n1698), .SI(\fifo[11][15] ), .SE(test_se), 
        .CLK(n39), .Q(\fifo[11][16] ), .QN(n1139) );
  SDFFX1 \fifo_reg[11][15]  ( .D(n1699), .SI(\fifo[11][14] ), .SE(test_se), 
        .CLK(n39), .Q(\fifo[11][15] ), .QN(n1140) );
  SDFFX1 \fifo_reg[11][14]  ( .D(n1700), .SI(\fifo[11][13] ), .SE(test_se), 
        .CLK(n39), .Q(\fifo[11][14] ), .QN(n1141) );
  SDFFX1 \fifo_reg[11][13]  ( .D(n1701), .SI(\fifo[11][12] ), .SE(test_se), 
        .CLK(n39), .Q(\fifo[11][13] ), .QN(n1142) );
  SDFFX1 \fifo_reg[11][12]  ( .D(n1702), .SI(\fifo[11][11] ), .SE(test_se), 
        .CLK(n39), .Q(\fifo[11][12] ), .QN(n1143) );
  SDFFX1 \fifo_reg[11][11]  ( .D(n1703), .SI(\fifo[11][10] ), .SE(test_se), 
        .CLK(n39), .Q(\fifo[11][11] ), .QN(n1144) );
  SDFFX1 \fifo_reg[11][10]  ( .D(n1704), .SI(\fifo[11][9] ), .SE(test_se), 
        .CLK(n39), .Q(\fifo[11][10] ), .QN(n1145) );
  SDFFX1 \fifo_reg[11][9]  ( .D(n1705), .SI(\fifo[11][8] ), .SE(test_se), 
        .CLK(n39), .Q(\fifo[11][9] ), .QN(n1146) );
  SDFFX1 \fifo_reg[11][8]  ( .D(n1706), .SI(\fifo[11][7] ), .SE(test_se), 
        .CLK(n39), .Q(\fifo[11][8] ), .QN(n1147) );
  SDFFX1 \fifo_reg[11][7]  ( .D(n1707), .SI(\fifo[11][6] ), .SE(test_se), 
        .CLK(n39), .Q(\fifo[11][7] ), .QN(n1148) );
  SDFFX1 \fifo_reg[11][6]  ( .D(n1708), .SI(\fifo[11][5] ), .SE(test_se), 
        .CLK(n39), .Q(\fifo[11][6] ), .QN(n1149) );
  SDFFX1 \fifo_reg[11][5]  ( .D(n1709), .SI(\fifo[11][4] ), .SE(test_se), 
        .CLK(n39), .Q(\fifo[11][5] ), .QN(n1150) );
  SDFFX1 \fifo_reg[11][4]  ( .D(n1710), .SI(\fifo[11][3] ), .SE(test_se), 
        .CLK(n39), .Q(\fifo[11][4] ), .QN(n1151) );
  SDFFX1 \fifo_reg[11][3]  ( .D(n1711), .SI(\fifo[11][2] ), .SE(test_se), 
        .CLK(n39), .Q(\fifo[11][3] ), .QN(n1152) );
  SDFFX1 \fifo_reg[11][2]  ( .D(n1712), .SI(\fifo[11][1] ), .SE(test_se), 
        .CLK(n38), .Q(\fifo[11][2] ), .QN(n1153) );
  SDFFX1 \fifo_reg[11][1]  ( .D(n1713), .SI(\fifo[11][0] ), .SE(test_se), 
        .CLK(n38), .Q(\fifo[11][1] ), .QN(n1154) );
  SDFFX1 \fifo_reg[11][0]  ( .D(n1714), .SI(\fifo[10][31] ), .SE(test_se), 
        .CLK(n38), .Q(\fifo[11][0] ), .QN(n1155) );
  SDFFX1 \fifo_reg[12][31]  ( .D(n1715), .SI(\fifo[12][30] ), .SE(test_se), 
        .CLK(n43), .Q(\fifo[12][31] ), .QN(n1156) );
  SDFFX1 \fifo_reg[12][30]  ( .D(n1716), .SI(\fifo[12][29] ), .SE(test_se), 
        .CLK(n43), .Q(\fifo[12][30] ), .QN(n1157) );
  SDFFX1 \fifo_reg[12][29]  ( .D(n1717), .SI(\fifo[12][28] ), .SE(test_se), 
        .CLK(n43), .Q(\fifo[12][29] ), .QN(n1158) );
  SDFFX1 \fifo_reg[12][28]  ( .D(n1718), .SI(\fifo[12][27] ), .SE(test_se), 
        .CLK(n43), .Q(\fifo[12][28] ), .QN(n1159) );
  SDFFX1 \fifo_reg[12][27]  ( .D(n1719), .SI(\fifo[12][26] ), .SE(test_se), 
        .CLK(n43), .Q(\fifo[12][27] ), .QN(n1160) );
  SDFFX1 \fifo_reg[12][26]  ( .D(n1720), .SI(\fifo[12][25] ), .SE(test_se), 
        .CLK(n43), .Q(\fifo[12][26] ), .QN(n1161) );
  SDFFX1 \fifo_reg[12][25]  ( .D(n1721), .SI(\fifo[12][24] ), .SE(test_se), 
        .CLK(n42), .Q(\fifo[12][25] ), .QN(n1162) );
  SDFFX1 \fifo_reg[12][24]  ( .D(n1722), .SI(\fifo[12][23] ), .SE(test_se), 
        .CLK(n42), .Q(\fifo[12][24] ), .QN(n1163) );
  SDFFX1 \fifo_reg[12][23]  ( .D(n1723), .SI(\fifo[12][22] ), .SE(test_se), 
        .CLK(n42), .Q(\fifo[12][23] ), .QN(n1164) );
  SDFFX1 \fifo_reg[12][22]  ( .D(n1724), .SI(\fifo[12][21] ), .SE(test_se), 
        .CLK(n42), .Q(\fifo[12][22] ), .QN(n1165) );
  SDFFX1 \fifo_reg[12][21]  ( .D(n1725), .SI(\fifo[12][20] ), .SE(test_se), 
        .CLK(n42), .Q(\fifo[12][21] ), .QN(n1166) );
  SDFFX1 \fifo_reg[12][20]  ( .D(n1726), .SI(\fifo[12][19] ), .SE(test_se), 
        .CLK(n42), .Q(\fifo[12][20] ), .QN(n1167) );
  SDFFX1 \fifo_reg[12][19]  ( .D(n1727), .SI(\fifo[12][18] ), .SE(test_se), 
        .CLK(n42), .Q(\fifo[12][19] ), .QN(n1168) );
  SDFFX1 \fifo_reg[12][18]  ( .D(n1728), .SI(\fifo[12][17] ), .SE(test_se), 
        .CLK(n42), .Q(\fifo[12][18] ), .QN(n1169) );
  SDFFX1 \fifo_reg[12][17]  ( .D(n1729), .SI(\fifo[12][16] ), .SE(test_se), 
        .CLK(n42), .Q(\fifo[12][17] ), .QN(n1170) );
  SDFFX1 \fifo_reg[12][16]  ( .D(n1730), .SI(\fifo[12][15] ), .SE(test_se), 
        .CLK(n42), .Q(\fifo[12][16] ), .QN(n1171) );
  SDFFX1 \fifo_reg[12][15]  ( .D(n1731), .SI(\fifo[12][14] ), .SE(test_se), 
        .CLK(n42), .Q(\fifo[12][15] ), .QN(n1172) );
  SDFFX1 \fifo_reg[12][14]  ( .D(n1732), .SI(\fifo[12][13] ), .SE(test_se), 
        .CLK(n42), .Q(\fifo[12][14] ), .QN(n1173) );
  SDFFX1 \fifo_reg[12][13]  ( .D(n1733), .SI(\fifo[12][12] ), .SE(test_se), 
        .CLK(n42), .Q(\fifo[12][13] ), .QN(n1174) );
  SDFFX1 \fifo_reg[12][12]  ( .D(n1734), .SI(\fifo[12][11] ), .SE(test_se), 
        .CLK(n42), .Q(\fifo[12][12] ), .QN(n1175) );
  SDFFX1 \fifo_reg[12][11]  ( .D(n1735), .SI(\fifo[12][10] ), .SE(test_se), 
        .CLK(n41), .Q(\fifo[12][11] ), .QN(n1176) );
  SDFFX1 \fifo_reg[12][10]  ( .D(n1736), .SI(\fifo[12][9] ), .SE(test_se), 
        .CLK(n41), .Q(\fifo[12][10] ), .QN(n1177) );
  SDFFX1 \fifo_reg[12][9]  ( .D(n1737), .SI(\fifo[12][8] ), .SE(test_se), 
        .CLK(n41), .Q(\fifo[12][9] ), .QN(n1178) );
  SDFFX1 \fifo_reg[12][8]  ( .D(n1738), .SI(\fifo[12][7] ), .SE(test_se), 
        .CLK(n41), .Q(\fifo[12][8] ), .QN(n1179) );
  SDFFX1 \fifo_reg[12][7]  ( .D(n1739), .SI(\fifo[12][6] ), .SE(test_se), 
        .CLK(n41), .Q(\fifo[12][7] ), .QN(n1180) );
  SDFFX1 \fifo_reg[12][6]  ( .D(n1740), .SI(\fifo[12][5] ), .SE(test_se), 
        .CLK(n41), .Q(\fifo[12][6] ), .QN(n1181) );
  SDFFX1 \fifo_reg[12][5]  ( .D(n1741), .SI(\fifo[12][4] ), .SE(test_se), 
        .CLK(n41), .Q(\fifo[12][5] ), .QN(n1182) );
  SDFFX1 \fifo_reg[12][4]  ( .D(n1742), .SI(\fifo[12][3] ), .SE(test_se), 
        .CLK(n41), .Q(\fifo[12][4] ), .QN(n1183) );
  SDFFX1 \fifo_reg[12][3]  ( .D(n1743), .SI(\fifo[12][2] ), .SE(test_se), 
        .CLK(n41), .Q(\fifo[12][3] ), .QN(n1184) );
  SDFFX1 \fifo_reg[12][2]  ( .D(n1744), .SI(\fifo[12][1] ), .SE(test_se), 
        .CLK(n41), .Q(\fifo[12][2] ), .QN(n1185) );
  SDFFX1 \fifo_reg[12][1]  ( .D(n1745), .SI(\fifo[12][0] ), .SE(test_se), 
        .CLK(n41), .Q(\fifo[12][1] ), .QN(n1186) );
  SDFFX1 \fifo_reg[12][0]  ( .D(n1746), .SI(\fifo[11][31] ), .SE(test_se), 
        .CLK(n41), .Q(\fifo[12][0] ), .QN(n1187) );
  SDFFX1 \fifo_reg[13][31]  ( .D(n1747), .SI(\fifo[13][30] ), .SE(test_se), 
        .CLK(n26), .Q(\fifo[13][31] ), .QN(n1188) );
  SDFFX1 \fifo_reg[13][30]  ( .D(n1748), .SI(\fifo[13][29] ), .SE(test_se), 
        .CLK(n25), .Q(\fifo[13][30] ), .QN(n1189) );
  SDFFX1 \fifo_reg[13][29]  ( .D(n1749), .SI(\fifo[13][28] ), .SE(test_se), 
        .CLK(n25), .Q(\fifo[13][29] ), .QN(n1190) );
  SDFFX1 \fifo_reg[13][28]  ( .D(n1750), .SI(\fifo[13][27] ), .SE(test_se), 
        .CLK(n25), .Q(\fifo[13][28] ), .QN(n1191) );
  SDFFX1 \fifo_reg[13][27]  ( .D(n1751), .SI(\fifo[13][26] ), .SE(test_se), 
        .CLK(n25), .Q(\fifo[13][27] ), .QN(n1192) );
  SDFFX1 \fifo_reg[13][26]  ( .D(n1752), .SI(\fifo[13][25] ), .SE(test_se), 
        .CLK(n25), .Q(\fifo[13][26] ), .QN(n1193) );
  SDFFX1 \fifo_reg[13][25]  ( .D(n1753), .SI(\fifo[13][24] ), .SE(test_se), 
        .CLK(n25), .Q(\fifo[13][25] ), .QN(n1194) );
  SDFFX1 \fifo_reg[13][24]  ( .D(n1754), .SI(\fifo[13][23] ), .SE(test_se), 
        .CLK(n25), .Q(\fifo[13][24] ), .QN(n1195) );
  SDFFX1 \fifo_reg[13][23]  ( .D(n1755), .SI(\fifo[13][22] ), .SE(test_se), 
        .CLK(n25), .Q(\fifo[13][23] ), .QN(n1196) );
  SDFFX1 \fifo_reg[13][22]  ( .D(n1756), .SI(\fifo[13][21] ), .SE(test_se), 
        .CLK(n25), .Q(\fifo[13][22] ), .QN(n1197) );
  SDFFX1 \fifo_reg[13][21]  ( .D(n1757), .SI(\fifo[13][20] ), .SE(test_se), 
        .CLK(n30), .Q(\fifo[13][21] ), .QN(n1198) );
  SDFFX1 \fifo_reg[13][20]  ( .D(n1758), .SI(\fifo[13][19] ), .SE(test_se), 
        .CLK(n44), .Q(\fifo[13][20] ), .QN(n1199) );
  SDFFX1 \fifo_reg[13][19]  ( .D(n1759), .SI(\fifo[13][18] ), .SE(test_se), 
        .CLK(n44), .Q(\fifo[13][19] ), .QN(n1200) );
  SDFFX1 \fifo_reg[13][18]  ( .D(n1760), .SI(\fifo[13][17] ), .SE(test_se), 
        .CLK(n44), .Q(\fifo[13][18] ), .QN(n1201) );
  SDFFX1 \fifo_reg[13][17]  ( .D(n1761), .SI(\fifo[13][16] ), .SE(test_se), 
        .CLK(n44), .Q(\fifo[13][17] ), .QN(n1202) );
  SDFFX1 \fifo_reg[13][16]  ( .D(n1762), .SI(\fifo[13][15] ), .SE(test_se), 
        .CLK(n44), .Q(\fifo[13][16] ), .QN(n1203) );
  SDFFX1 \fifo_reg[13][15]  ( .D(n1763), .SI(\fifo[13][14] ), .SE(test_se), 
        .CLK(n44), .Q(\fifo[13][15] ), .QN(n1204) );
  SDFFX1 \fifo_reg[13][14]  ( .D(n1764), .SI(\fifo[13][13] ), .SE(test_se), 
        .CLK(n44), .Q(\fifo[13][14] ), .QN(n1205) );
  SDFFX1 \fifo_reg[13][13]  ( .D(n1765), .SI(\fifo[13][12] ), .SE(test_se), 
        .CLK(n44), .Q(\fifo[13][13] ), .QN(n1206) );
  SDFFX1 \fifo_reg[13][12]  ( .D(n1766), .SI(\fifo[13][11] ), .SE(test_se), 
        .CLK(n44), .Q(\fifo[13][12] ), .QN(n1207) );
  SDFFX1 \fifo_reg[13][11]  ( .D(n1767), .SI(\fifo[13][10] ), .SE(test_se), 
        .CLK(n44), .Q(\fifo[13][11] ), .QN(n1208) );
  SDFFX1 \fifo_reg[13][10]  ( .D(n1768), .SI(\fifo[13][9] ), .SE(test_se), 
        .CLK(n44), .Q(\fifo[13][10] ), .QN(n1209) );
  SDFFX1 \fifo_reg[13][9]  ( .D(n1769), .SI(\fifo[13][8] ), .SE(test_se), 
        .CLK(n44), .Q(\fifo[13][9] ), .QN(n1210) );
  SDFFX1 \fifo_reg[13][8]  ( .D(n1770), .SI(\fifo[13][7] ), .SE(test_se), 
        .CLK(n44), .Q(\fifo[13][8] ), .QN(n1211) );
  SDFFX1 \fifo_reg[13][7]  ( .D(n1771), .SI(\fifo[13][6] ), .SE(test_se), 
        .CLK(n43), .Q(\fifo[13][7] ), .QN(n1212) );
  SDFFX1 \fifo_reg[13][6]  ( .D(n1772), .SI(\fifo[13][5] ), .SE(test_se), 
        .CLK(n43), .Q(\fifo[13][6] ), .QN(n1213) );
  SDFFX1 \fifo_reg[13][5]  ( .D(n1773), .SI(\fifo[13][4] ), .SE(test_se), 
        .CLK(n43), .Q(\fifo[13][5] ), .QN(n1214) );
  SDFFX1 \fifo_reg[13][4]  ( .D(n1774), .SI(\fifo[13][3] ), .SE(test_se), 
        .CLK(n43), .Q(\fifo[13][4] ), .QN(n1215) );
  SDFFX1 \fifo_reg[13][3]  ( .D(n1775), .SI(\fifo[13][2] ), .SE(test_se), 
        .CLK(n43), .Q(\fifo[13][3] ), .QN(n1216) );
  SDFFX1 \fifo_reg[13][2]  ( .D(n1776), .SI(\fifo[13][1] ), .SE(test_se), 
        .CLK(n43), .Q(\fifo[13][2] ), .QN(n1217) );
  SDFFX1 \fifo_reg[13][1]  ( .D(n1777), .SI(\fifo[13][0] ), .SE(test_se), 
        .CLK(n43), .Q(\fifo[13][1] ), .QN(n1218) );
  SDFFX1 \fifo_reg[13][0]  ( .D(n1778), .SI(\fifo[12][31] ), .SE(test_se), 
        .CLK(n43), .Q(\fifo[13][0] ), .QN(n1219) );
  SDFFX1 \fifo_reg[14][31]  ( .D(n1779), .SI(\fifo[14][30] ), .SE(test_se), 
        .CLK(n28), .Q(\fifo[14][31] ), .QN(n1220) );
  SDFFX1 \fifo_reg[14][30]  ( .D(n1780), .SI(\fifo[14][29] ), .SE(test_se), 
        .CLK(n28), .Q(\fifo[14][30] ), .QN(n1221) );
  SDFFX1 \fifo_reg[14][29]  ( .D(n1781), .SI(\fifo[14][28] ), .SE(test_se), 
        .CLK(n28), .Q(\fifo[14][29] ), .QN(n1222) );
  SDFFX1 \fifo_reg[14][28]  ( .D(n1782), .SI(\fifo[14][27] ), .SE(test_se), 
        .CLK(n28), .Q(\fifo[14][28] ), .QN(n1223) );
  SDFFX1 \fifo_reg[14][27]  ( .D(n1783), .SI(\fifo[14][26] ), .SE(test_se), 
        .CLK(n28), .Q(\fifo[14][27] ), .QN(n1224) );
  SDFFX1 \fifo_reg[14][26]  ( .D(n1784), .SI(\fifo[14][25] ), .SE(test_se), 
        .CLK(n27), .Q(\fifo[14][26] ), .QN(n1225) );
  SDFFX1 \fifo_reg[14][25]  ( .D(n1785), .SI(\fifo[14][24] ), .SE(test_se), 
        .CLK(n27), .Q(\fifo[14][25] ), .QN(n1226) );
  SDFFX1 \fifo_reg[14][24]  ( .D(n1786), .SI(\fifo[14][23] ), .SE(test_se), 
        .CLK(n27), .Q(\fifo[14][24] ), .QN(n1227) );
  SDFFX1 \fifo_reg[14][23]  ( .D(n1787), .SI(\fifo[14][22] ), .SE(test_se), 
        .CLK(n27), .Q(\fifo[14][23] ), .QN(n1228) );
  SDFFX1 \fifo_reg[14][22]  ( .D(n1788), .SI(\fifo[14][21] ), .SE(test_se), 
        .CLK(n27), .Q(\fifo[14][22] ), .QN(n1229) );
  SDFFX1 \fifo_reg[14][21]  ( .D(n1789), .SI(\fifo[14][20] ), .SE(test_se), 
        .CLK(n27), .Q(\fifo[14][21] ), .QN(n1230) );
  SDFFX1 \fifo_reg[14][20]  ( .D(n1790), .SI(\fifo[14][19] ), .SE(test_se), 
        .CLK(n27), .Q(\fifo[14][20] ), .QN(n1231) );
  SDFFX1 \fifo_reg[14][19]  ( .D(n1791), .SI(\fifo[14][18] ), .SE(test_se), 
        .CLK(n27), .Q(\fifo[14][19] ), .QN(n1232) );
  SDFFX1 \fifo_reg[14][18]  ( .D(n1792), .SI(\fifo[14][17] ), .SE(test_se), 
        .CLK(n27), .Q(\fifo[14][18] ), .QN(n1233) );
  SDFFX1 \fifo_reg[14][17]  ( .D(n1793), .SI(\fifo[14][16] ), .SE(test_se), 
        .CLK(n27), .Q(\fifo[14][17] ), .QN(n1234) );
  SDFFX1 \fifo_reg[14][16]  ( .D(n1794), .SI(\fifo[14][15] ), .SE(test_se), 
        .CLK(n27), .Q(\fifo[14][16] ), .QN(n1235) );
  SDFFX1 \fifo_reg[14][15]  ( .D(n1795), .SI(\fifo[14][14] ), .SE(test_se), 
        .CLK(n27), .Q(\fifo[14][15] ), .QN(n1236) );
  SDFFX1 \fifo_reg[14][14]  ( .D(n1796), .SI(\fifo[14][13] ), .SE(test_se), 
        .CLK(n27), .Q(\fifo[14][14] ), .QN(n1237) );
  SDFFX1 \fifo_reg[14][13]  ( .D(n1797), .SI(\fifo[14][12] ), .SE(test_se), 
        .CLK(n27), .Q(\fifo[14][13] ), .QN(n1238) );
  SDFFX1 \fifo_reg[14][12]  ( .D(n1798), .SI(\fifo[14][11] ), .SE(test_se), 
        .CLK(n26), .Q(\fifo[14][12] ), .QN(n1239) );
  SDFFX1 \fifo_reg[14][11]  ( .D(n1799), .SI(\fifo[14][10] ), .SE(test_se), 
        .CLK(n26), .Q(\fifo[14][11] ), .QN(n1240) );
  SDFFX1 \fifo_reg[14][10]  ( .D(n1800), .SI(\fifo[14][9] ), .SE(test_se), 
        .CLK(n26), .Q(\fifo[14][10] ), .QN(n1241) );
  SDFFX1 \fifo_reg[14][9]  ( .D(n1801), .SI(\fifo[14][8] ), .SE(test_se), 
        .CLK(n26), .Q(\fifo[14][9] ), .QN(n1242) );
  SDFFX1 \fifo_reg[14][8]  ( .D(n1802), .SI(\fifo[14][7] ), .SE(test_se), 
        .CLK(n26), .Q(\fifo[14][8] ), .QN(n1243) );
  SDFFX1 \fifo_reg[14][7]  ( .D(n1803), .SI(\fifo[14][6] ), .SE(test_se), 
        .CLK(n26), .Q(\fifo[14][7] ), .QN(n1244) );
  SDFFX1 \fifo_reg[14][6]  ( .D(n1804), .SI(\fifo[14][5] ), .SE(test_se), 
        .CLK(n26), .Q(\fifo[14][6] ), .QN(n1245) );
  SDFFX1 \fifo_reg[14][5]  ( .D(n1805), .SI(\fifo[14][4] ), .SE(test_se), 
        .CLK(n26), .Q(\fifo[14][5] ), .QN(n1246) );
  SDFFX1 \fifo_reg[14][4]  ( .D(n1806), .SI(\fifo[14][3] ), .SE(test_se), 
        .CLK(n26), .Q(\fifo[14][4] ), .QN(n1247) );
  SDFFX1 \fifo_reg[14][3]  ( .D(n1807), .SI(\fifo[14][2] ), .SE(test_se), 
        .CLK(n26), .Q(\fifo[14][3] ), .QN(n1248) );
  SDFFX1 \fifo_reg[14][2]  ( .D(n1808), .SI(\fifo[14][1] ), .SE(test_se), 
        .CLK(n26), .Q(\fifo[14][2] ), .QN(n1249) );
  SDFFX1 \fifo_reg[14][1]  ( .D(n1809), .SI(\fifo[14][0] ), .SE(test_se), 
        .CLK(n26), .Q(\fifo[14][1] ), .QN(n1250) );
  SDFFX1 \fifo_reg[14][0]  ( .D(n1810), .SI(\fifo[13][31] ), .SE(test_se), 
        .CLK(n26), .Q(\fifo[14][0] ), .QN(n1251) );
  SDFFX1 \fifo_reg[15][31]  ( .D(n1811), .SI(\fifo[15][30] ), .SE(test_se), 
        .CLK(n30), .Q(\fifo[15][31] ), .QN(n1252) );
  SDFFX1 \fifo_reg[15][30]  ( .D(n1812), .SI(\fifo[15][29] ), .SE(test_se), 
        .CLK(n30), .Q(\fifo[15][30] ), .QN(n1253) );
  SDFFX1 \fifo_reg[15][29]  ( .D(n1813), .SI(\fifo[15][28] ), .SE(test_se), 
        .CLK(n30), .Q(\fifo[15][29] ), .QN(n1254) );
  SDFFX1 \fifo_reg[15][28]  ( .D(n1814), .SI(\fifo[15][27] ), .SE(test_se), 
        .CLK(n30), .Q(\fifo[15][28] ), .QN(n1255) );
  SDFFX1 \fifo_reg[15][27]  ( .D(n1815), .SI(\fifo[15][26] ), .SE(test_se), 
        .CLK(n30), .Q(\fifo[15][27] ), .QN(n1256) );
  SDFFX1 \fifo_reg[15][26]  ( .D(n1816), .SI(\fifo[15][25] ), .SE(test_se), 
        .CLK(n30), .Q(\fifo[15][26] ), .QN(n1257) );
  SDFFX1 \fifo_reg[15][25]  ( .D(n1817), .SI(\fifo[15][24] ), .SE(test_se), 
        .CLK(n30), .Q(\fifo[15][25] ), .QN(n1258) );
  SDFFX1 \fifo_reg[15][24]  ( .D(n1818), .SI(\fifo[15][23] ), .SE(test_se), 
        .CLK(n30), .Q(\fifo[15][24] ), .QN(n1259) );
  SDFFX1 \fifo_reg[15][23]  ( .D(n1819), .SI(\fifo[15][22] ), .SE(test_se), 
        .CLK(n30), .Q(\fifo[15][23] ), .QN(n1260) );
  SDFFX1 \fifo_reg[15][22]  ( .D(n1820), .SI(\fifo[15][21] ), .SE(test_se), 
        .CLK(n29), .Q(\fifo[15][22] ), .QN(n1261) );
  SDFFX1 \fifo_reg[15][21]  ( .D(n1821), .SI(\fifo[15][20] ), .SE(test_se), 
        .CLK(n29), .Q(\fifo[15][21] ), .QN(n1262) );
  SDFFX1 \fifo_reg[15][20]  ( .D(n1822), .SI(\fifo[15][19] ), .SE(test_se), 
        .CLK(n29), .Q(\fifo[15][20] ), .QN(n1263) );
  SDFFX1 \fifo_reg[15][19]  ( .D(n1823), .SI(\fifo[15][18] ), .SE(test_se), 
        .CLK(n29), .Q(\fifo[15][19] ), .QN(n1264) );
  SDFFX1 \fifo_reg[15][18]  ( .D(n1824), .SI(\fifo[15][17] ), .SE(test_se), 
        .CLK(n29), .Q(\fifo[15][18] ), .QN(n1265) );
  SDFFX1 \fifo_reg[15][17]  ( .D(n1825), .SI(\fifo[15][16] ), .SE(test_se), 
        .CLK(n29), .Q(\fifo[15][17] ), .QN(n1266) );
  SDFFX1 \fifo_reg[15][16]  ( .D(n1826), .SI(\fifo[15][15] ), .SE(test_se), 
        .CLK(n29), .Q(\fifo[15][16] ), .QN(n1267) );
  SDFFX1 \fifo_reg[15][15]  ( .D(n1827), .SI(\fifo[15][14] ), .SE(test_se), 
        .CLK(n29), .Q(\fifo[15][15] ), .QN(n1268) );
  SDFFX1 \fifo_reg[15][14]  ( .D(n1828), .SI(\fifo[15][13] ), .SE(test_se), 
        .CLK(n29), .Q(\fifo[15][14] ), .QN(n1269) );
  SDFFX1 \fifo_reg[15][13]  ( .D(n1829), .SI(\fifo[15][12] ), .SE(test_se), 
        .CLK(n29), .Q(\fifo[15][13] ), .QN(n1270) );
  SDFFX1 \fifo_reg[15][12]  ( .D(n1830), .SI(\fifo[15][11] ), .SE(test_se), 
        .CLK(n29), .Q(\fifo[15][12] ), .QN(n1271) );
  SDFFX1 \fifo_reg[15][11]  ( .D(n1831), .SI(\fifo[15][10] ), .SE(test_se), 
        .CLK(n29), .Q(\fifo[15][11] ), .QN(n1272) );
  SDFFX1 \fifo_reg[15][10]  ( .D(n1832), .SI(\fifo[15][9] ), .SE(test_se), 
        .CLK(n29), .Q(\fifo[15][10] ), .QN(n1273) );
  SDFFX1 \fifo_reg[15][9]  ( .D(n1833), .SI(\fifo[15][8] ), .SE(test_se), 
        .CLK(n29), .Q(\fifo[15][9] ), .QN(n1274) );
  SDFFX1 \fifo_reg[15][8]  ( .D(n1834), .SI(\fifo[15][7] ), .SE(test_se), 
        .CLK(n28), .Q(\fifo[15][8] ), .QN(n1275) );
  SDFFX1 \fifo_reg[15][7]  ( .D(n1835), .SI(\fifo[15][6] ), .SE(test_se), 
        .CLK(n28), .Q(\fifo[15][7] ), .QN(n1276) );
  SDFFX1 \fifo_reg[15][6]  ( .D(n1836), .SI(\fifo[15][5] ), .SE(test_se), 
        .CLK(n28), .Q(\fifo[15][6] ), .QN(n1277) );
  SDFFX1 \fifo_reg[15][5]  ( .D(n1837), .SI(\fifo[15][4] ), .SE(test_se), 
        .CLK(n28), .Q(\fifo[15][5] ), .QN(n1278) );
  SDFFX1 \fifo_reg[15][4]  ( .D(n1838), .SI(\fifo[15][3] ), .SE(test_se), 
        .CLK(n28), .Q(\fifo[15][4] ), .QN(n1279) );
  SDFFX1 \fifo_reg[15][3]  ( .D(n1839), .SI(\fifo[15][2] ), .SE(test_se), 
        .CLK(n28), .Q(\fifo[15][3] ), .QN(n1280) );
  SDFFX1 \fifo_reg[15][2]  ( .D(n1840), .SI(\fifo[15][1] ), .SE(test_se), 
        .CLK(n28), .Q(\fifo[15][2] ), .QN(n1281) );
  SDFFX1 \fifo_reg[15][1]  ( .D(n1841), .SI(\fifo[15][0] ), .SE(test_se), 
        .CLK(n28), .Q(\fifo[15][1] ), .QN(n1282) );
  SDFFX1 \fifo_reg[15][0]  ( .D(n1842), .SI(\fifo[14][31] ), .SE(test_se), 
        .CLK(n28), .Q(\fifo[15][0] ), .QN(n1283) );
  SDFFX1 \data_out_reg[31]  ( .D(N155), .SI(test_si2), .SE(test_se), .CLK(n6), 
        .Q(data_out[31]) );
  SDFFX1 \data_out_reg[30]  ( .D(N154), .SI(data_out[29]), .SE(test_se), .CLK(
        n32), .Q(data_out[30]) );
  SDFFX1 \data_out_reg[29]  ( .D(N153), .SI(data_out[28]), .SE(test_se), .CLK(
        n32), .Q(data_out[29]) );
  SDFFX1 \data_out_reg[28]  ( .D(N152), .SI(data_out[27]), .SE(test_se), .CLK(
        n32), .Q(data_out[28]) );
  SDFFX1 \data_out_reg[27]  ( .D(N151), .SI(data_out[26]), .SE(test_se), .CLK(
        n32), .Q(data_out[27]) );
  SDFFX1 \data_out_reg[26]  ( .D(N150), .SI(data_out[25]), .SE(test_se), .CLK(
        n32), .Q(data_out[26]) );
  SDFFX1 \data_out_reg[25]  ( .D(N149), .SI(data_out[24]), .SE(test_se), .CLK(
        n32), .Q(data_out[25]) );
  SDFFX1 \data_out_reg[24]  ( .D(N148), .SI(data_out[23]), .SE(test_se), .CLK(
        n32), .Q(data_out[24]) );
  SDFFX1 \data_out_reg[23]  ( .D(N147), .SI(data_out[22]), .SE(test_se), .CLK(
        n32), .Q(data_out[23]) );
  SDFFX1 \data_out_reg[22]  ( .D(N146), .SI(data_out[21]), .SE(test_se), .CLK(
        n32), .Q(data_out[22]) );
  SDFFX1 \data_out_reg[21]  ( .D(N145), .SI(data_out[20]), .SE(test_se), .CLK(
        n32), .Q(data_out[21]) );
  SDFFX1 \data_out_reg[20]  ( .D(N144), .SI(data_out[19]), .SE(test_se), .CLK(
        n32), .Q(data_out[20]) );
  SDFFX1 \data_out_reg[19]  ( .D(N143), .SI(data_out[18]), .SE(test_se), .CLK(
        n32), .Q(data_out[19]) );
  SDFFX1 \data_out_reg[18]  ( .D(N142), .SI(data_out[17]), .SE(test_se), .CLK(
        n32), .Q(data_out[18]) );
  SDFFX1 \data_out_reg[17]  ( .D(N141), .SI(data_out[16]), .SE(test_se), .CLK(
        n31), .Q(data_out[17]) );
  SDFFX1 \data_out_reg[16]  ( .D(N140), .SI(data_out[15]), .SE(test_se), .CLK(
        n31), .Q(data_out[16]) );
  SDFFX1 \data_out_reg[15]  ( .D(N139), .SI(data_out[14]), .SE(test_se), .CLK(
        n31), .Q(data_out[15]) );
  SDFFX1 \data_out_reg[14]  ( .D(N138), .SI(data_out[13]), .SE(test_se), .CLK(
        n31), .Q(data_out[14]) );
  SDFFX1 \data_out_reg[13]  ( .D(N137), .SI(data_out[12]), .SE(test_se), .CLK(
        n31), .Q(data_out[13]) );
  SDFFX1 \data_out_reg[12]  ( .D(N136), .SI(data_out[11]), .SE(test_se), .CLK(
        n31), .Q(data_out[12]) );
  SDFFX1 \data_out_reg[11]  ( .D(N135), .SI(data_out[10]), .SE(test_se), .CLK(
        n31), .Q(data_out[11]) );
  SDFFX1 \data_out_reg[10]  ( .D(N134), .SI(data_out[9]), .SE(test_se), .CLK(
        n31), .Q(data_out[10]) );
  SDFFX1 \data_out_reg[9]  ( .D(N133), .SI(data_out[8]), .SE(test_se), .CLK(
        n31), .Q(data_out[9]) );
  SDFFX1 \data_out_reg[8]  ( .D(N132), .SI(data_out[7]), .SE(test_se), .CLK(
        n31), .Q(data_out[8]) );
  SDFFX1 \data_out_reg[7]  ( .D(N131), .SI(data_out[6]), .SE(test_se), .CLK(
        n31), .Q(data_out[7]) );
  SDFFX1 \data_out_reg[6]  ( .D(N130), .SI(data_out[5]), .SE(test_se), .CLK(
        n31), .Q(data_out[6]) );
  SDFFX1 \data_out_reg[5]  ( .D(N129), .SI(data_out[4]), .SE(test_se), .CLK(
        n31), .Q(data_out[5]) );
  SDFFX1 \data_out_reg[4]  ( .D(N128), .SI(data_out[3]), .SE(test_se), .CLK(
        n31), .Q(data_out[4]) );
  SDFFX1 \data_out_reg[3]  ( .D(N127), .SI(data_out[2]), .SE(test_se), .CLK(
        n30), .Q(data_out[3]) );
  SDFFX1 \data_out_reg[2]  ( .D(N126), .SI(data_out[1]), .SE(test_se), .CLK(
        n30), .Q(data_out[2]) );
  SDFFX1 \data_out_reg[1]  ( .D(N125), .SI(data_out[0]), .SE(test_se), .CLK(
        n30), .Q(data_out[1]) );
  SDFFX1 \data_out_reg[0]  ( .D(N124), .SI(cnt[4]), .SE(test_se), .CLK(n30), 
        .Q(data_out[0]) );
  NBUFFX2 U3 ( .INP(clk), .Z(n6) );
  NBUFFX2 U4 ( .INP(clk), .Z(n31) );
  NBUFFX2 U5 ( .INP(clk), .Z(n29) );
  NBUFFX2 U6 ( .INP(clk), .Z(n27) );
  NBUFFX2 U7 ( .INP(clk), .Z(n28) );
  NBUFFX2 U8 ( .INP(clk), .Z(n30) );
  NBUFFX2 U9 ( .INP(clk), .Z(n26) );
  NBUFFX2 U10 ( .INP(clk), .Z(n42) );
  NBUFFX2 U11 ( .INP(clk), .Z(n43) );
  NBUFFX2 U12 ( .INP(clk), .Z(n39) );
  NBUFFX2 U13 ( .INP(clk), .Z(n41) );
  NBUFFX2 U14 ( .INP(clk), .Z(n37) );
  NBUFFX2 U15 ( .INP(clk), .Z(n38) );
  NBUFFX2 U16 ( .INP(clk), .Z(n40) );
  NBUFFX2 U17 ( .INP(clk), .Z(n36) );
  NBUFFX2 U18 ( .INP(clk), .Z(n13) );
  NBUFFX2 U19 ( .INP(clk), .Z(n14) );
  NBUFFX2 U20 ( .INP(clk), .Z(n11) );
  NBUFFX2 U21 ( .INP(clk), .Z(n12) );
  NBUFFX2 U22 ( .INP(clk), .Z(n9) );
  NBUFFX2 U23 ( .INP(clk), .Z(n10) );
  NBUFFX2 U24 ( .INP(clk), .Z(n25) );
  NBUFFX2 U25 ( .INP(clk), .Z(n7) );
  NBUFFX2 U26 ( .INP(clk), .Z(n8) );
  NBUFFX2 U27 ( .INP(clk), .Z(n23) );
  NBUFFX2 U28 ( .INP(clk), .Z(n24) );
  NBUFFX2 U29 ( .INP(clk), .Z(n21) );
  NBUFFX2 U30 ( .INP(clk), .Z(n22) );
  NBUFFX2 U31 ( .INP(clk), .Z(n18) );
  NBUFFX2 U32 ( .INP(clk), .Z(n19) );
  NBUFFX2 U33 ( .INP(clk), .Z(n15) );
  NBUFFX2 U34 ( .INP(clk), .Z(n16) );
  NBUFFX2 U35 ( .INP(clk), .Z(n17) );
  NBUFFX2 U36 ( .INP(clk), .Z(n32) );
  NBUFFX2 U37 ( .INP(clk), .Z(n33) );
  NBUFFX2 U38 ( .INP(clk), .Z(n34) );
  NBUFFX2 U39 ( .INP(clk), .Z(n35) );
  NBUFFX2 U40 ( .INP(clk), .Z(n20) );
  NBUFFX2 U41 ( .INP(clk), .Z(n5) );
  NBUFFX2 U42 ( .INP(clk), .Z(n44) );
  INVX0 U43 ( .INP(n45), .ZN(full) );
  INVX0 U44 ( .INP(eth_top_test_point_11887_in), .ZN(n428) );
  MUX21X1 U45 ( .IN1(\fifo[15][0] ), .IN2(data_in[0]), .S(n46), .Q(n1842) );
  MUX21X1 U46 ( .IN1(\fifo[15][1] ), .IN2(data_in[1]), .S(n46), .Q(n1841) );
  MUX21X1 U47 ( .IN1(\fifo[15][2] ), .IN2(data_in[2]), .S(n46), .Q(n1840) );
  MUX21X1 U48 ( .IN1(\fifo[15][3] ), .IN2(data_in[3]), .S(n46), .Q(n1839) );
  MUX21X1 U49 ( .IN1(\fifo[15][4] ), .IN2(data_in[4]), .S(n46), .Q(n1838) );
  MUX21X1 U50 ( .IN1(\fifo[15][5] ), .IN2(data_in[5]), .S(n46), .Q(n1837) );
  MUX21X1 U51 ( .IN1(\fifo[15][6] ), .IN2(data_in[6]), .S(n46), .Q(n1836) );
  MUX21X1 U52 ( .IN1(\fifo[15][7] ), .IN2(data_in[7]), .S(n46), .Q(n1835) );
  MUX21X1 U53 ( .IN1(\fifo[15][8] ), .IN2(data_in[8]), .S(n46), .Q(n1834) );
  MUX21X1 U54 ( .IN1(\fifo[15][9] ), .IN2(data_in[9]), .S(n46), .Q(n1833) );
  MUX21X1 U55 ( .IN1(\fifo[15][10] ), .IN2(data_in[10]), .S(n46), .Q(n1832) );
  MUX21X1 U56 ( .IN1(\fifo[15][11] ), .IN2(data_in[11]), .S(n46), .Q(n1831) );
  MUX21X1 U57 ( .IN1(\fifo[15][12] ), .IN2(data_in[12]), .S(n46), .Q(n1830) );
  MUX21X1 U58 ( .IN1(\fifo[15][13] ), .IN2(data_in[13]), .S(n46), .Q(n1829) );
  MUX21X1 U59 ( .IN1(\fifo[15][14] ), .IN2(data_in[14]), .S(n46), .Q(n1828) );
  MUX21X1 U60 ( .IN1(\fifo[15][15] ), .IN2(data_in[15]), .S(n46), .Q(n1827) );
  MUX21X1 U61 ( .IN1(\fifo[15][16] ), .IN2(data_in[16]), .S(n46), .Q(n1826) );
  MUX21X1 U62 ( .IN1(\fifo[15][17] ), .IN2(data_in[17]), .S(n46), .Q(n1825) );
  MUX21X1 U63 ( .IN1(\fifo[15][18] ), .IN2(data_in[18]), .S(n46), .Q(n1824) );
  MUX21X1 U64 ( .IN1(\fifo[15][19] ), .IN2(data_in[19]), .S(n46), .Q(n1823) );
  MUX21X1 U65 ( .IN1(\fifo[15][20] ), .IN2(data_in[20]), .S(n46), .Q(n1822) );
  MUX21X1 U66 ( .IN1(\fifo[15][21] ), .IN2(data_in[21]), .S(n46), .Q(n1821) );
  MUX21X1 U67 ( .IN1(\fifo[15][22] ), .IN2(data_in[22]), .S(n46), .Q(n1820) );
  MUX21X1 U68 ( .IN1(\fifo[15][23] ), .IN2(data_in[23]), .S(n46), .Q(n1819) );
  MUX21X1 U69 ( .IN1(\fifo[15][24] ), .IN2(data_in[24]), .S(n46), .Q(n1818) );
  MUX21X1 U70 ( .IN1(\fifo[15][25] ), .IN2(data_in[25]), .S(n46), .Q(n1817) );
  MUX21X1 U71 ( .IN1(\fifo[15][26] ), .IN2(data_in[26]), .S(n46), .Q(n1816) );
  MUX21X1 U72 ( .IN1(\fifo[15][27] ), .IN2(data_in[27]), .S(n46), .Q(n1815) );
  MUX21X1 U73 ( .IN1(\fifo[15][28] ), .IN2(data_in[28]), .S(n46), .Q(n1814) );
  MUX21X1 U74 ( .IN1(\fifo[15][29] ), .IN2(data_in[29]), .S(n46), .Q(n1813) );
  MUX21X1 U75 ( .IN1(\fifo[15][30] ), .IN2(data_in[30]), .S(n46), .Q(n1812) );
  MUX21X1 U76 ( .IN1(\fifo[15][31] ), .IN2(data_in[31]), .S(n46), .Q(n1811) );
  AND2X1 U77 ( .IN1(n47), .IN2(n48), .Q(n46) );
  MUX21X1 U78 ( .IN1(\fifo[14][0] ), .IN2(data_in[0]), .S(n49), .Q(n1810) );
  MUX21X1 U79 ( .IN1(\fifo[14][1] ), .IN2(data_in[1]), .S(n49), .Q(n1809) );
  MUX21X1 U80 ( .IN1(\fifo[14][2] ), .IN2(data_in[2]), .S(n49), .Q(n1808) );
  MUX21X1 U81 ( .IN1(\fifo[14][3] ), .IN2(data_in[3]), .S(n49), .Q(n1807) );
  MUX21X1 U82 ( .IN1(\fifo[14][4] ), .IN2(data_in[4]), .S(n49), .Q(n1806) );
  MUX21X1 U83 ( .IN1(\fifo[14][5] ), .IN2(data_in[5]), .S(n49), .Q(n1805) );
  MUX21X1 U84 ( .IN1(\fifo[14][6] ), .IN2(data_in[6]), .S(n49), .Q(n1804) );
  MUX21X1 U85 ( .IN1(\fifo[14][7] ), .IN2(data_in[7]), .S(n49), .Q(n1803) );
  MUX21X1 U86 ( .IN1(\fifo[14][8] ), .IN2(data_in[8]), .S(n49), .Q(n1802) );
  MUX21X1 U87 ( .IN1(\fifo[14][9] ), .IN2(data_in[9]), .S(n49), .Q(n1801) );
  MUX21X1 U88 ( .IN1(\fifo[14][10] ), .IN2(data_in[10]), .S(n49), .Q(n1800) );
  MUX21X1 U89 ( .IN1(\fifo[14][11] ), .IN2(data_in[11]), .S(n49), .Q(n1799) );
  MUX21X1 U90 ( .IN1(\fifo[14][12] ), .IN2(data_in[12]), .S(n49), .Q(n1798) );
  MUX21X1 U91 ( .IN1(\fifo[14][13] ), .IN2(data_in[13]), .S(n49), .Q(n1797) );
  MUX21X1 U92 ( .IN1(\fifo[14][14] ), .IN2(data_in[14]), .S(n49), .Q(n1796) );
  MUX21X1 U93 ( .IN1(\fifo[14][15] ), .IN2(data_in[15]), .S(n49), .Q(n1795) );
  MUX21X1 U94 ( .IN1(\fifo[14][16] ), .IN2(data_in[16]), .S(n49), .Q(n1794) );
  MUX21X1 U95 ( .IN1(\fifo[14][17] ), .IN2(data_in[17]), .S(n49), .Q(n1793) );
  MUX21X1 U96 ( .IN1(\fifo[14][18] ), .IN2(data_in[18]), .S(n49), .Q(n1792) );
  MUX21X1 U97 ( .IN1(\fifo[14][19] ), .IN2(data_in[19]), .S(n49), .Q(n1791) );
  MUX21X1 U98 ( .IN1(\fifo[14][20] ), .IN2(data_in[20]), .S(n49), .Q(n1790) );
  MUX21X1 U99 ( .IN1(\fifo[14][21] ), .IN2(data_in[21]), .S(n49), .Q(n1789) );
  MUX21X1 U100 ( .IN1(\fifo[14][22] ), .IN2(data_in[22]), .S(n49), .Q(n1788)
         );
  MUX21X1 U101 ( .IN1(\fifo[14][23] ), .IN2(data_in[23]), .S(n49), .Q(n1787)
         );
  MUX21X1 U102 ( .IN1(\fifo[14][24] ), .IN2(data_in[24]), .S(n49), .Q(n1786)
         );
  MUX21X1 U103 ( .IN1(\fifo[14][25] ), .IN2(data_in[25]), .S(n49), .Q(n1785)
         );
  MUX21X1 U104 ( .IN1(\fifo[14][26] ), .IN2(data_in[26]), .S(n49), .Q(n1784)
         );
  MUX21X1 U105 ( .IN1(\fifo[14][27] ), .IN2(data_in[27]), .S(n49), .Q(n1783)
         );
  MUX21X1 U106 ( .IN1(\fifo[14][28] ), .IN2(data_in[28]), .S(n49), .Q(n1782)
         );
  MUX21X1 U107 ( .IN1(\fifo[14][29] ), .IN2(data_in[29]), .S(n49), .Q(n1781)
         );
  MUX21X1 U108 ( .IN1(\fifo[14][30] ), .IN2(data_in[30]), .S(n49), .Q(n1780)
         );
  MUX21X1 U109 ( .IN1(\fifo[14][31] ), .IN2(data_in[31]), .S(n49), .Q(n1779)
         );
  AND2X1 U110 ( .IN1(n50), .IN2(n48), .Q(n49) );
  MUX21X1 U111 ( .IN1(\fifo[13][0] ), .IN2(data_in[0]), .S(n51), .Q(n1778) );
  MUX21X1 U112 ( .IN1(\fifo[13][1] ), .IN2(data_in[1]), .S(n51), .Q(n1777) );
  MUX21X1 U113 ( .IN1(\fifo[13][2] ), .IN2(data_in[2]), .S(n51), .Q(n1776) );
  MUX21X1 U114 ( .IN1(\fifo[13][3] ), .IN2(data_in[3]), .S(n51), .Q(n1775) );
  MUX21X1 U115 ( .IN1(\fifo[13][4] ), .IN2(data_in[4]), .S(n51), .Q(n1774) );
  MUX21X1 U116 ( .IN1(\fifo[13][5] ), .IN2(data_in[5]), .S(n51), .Q(n1773) );
  MUX21X1 U117 ( .IN1(\fifo[13][6] ), .IN2(data_in[6]), .S(n51), .Q(n1772) );
  MUX21X1 U118 ( .IN1(\fifo[13][7] ), .IN2(data_in[7]), .S(n51), .Q(n1771) );
  MUX21X1 U119 ( .IN1(\fifo[13][8] ), .IN2(data_in[8]), .S(n51), .Q(n1770) );
  MUX21X1 U120 ( .IN1(\fifo[13][9] ), .IN2(data_in[9]), .S(n51), .Q(n1769) );
  MUX21X1 U121 ( .IN1(\fifo[13][10] ), .IN2(data_in[10]), .S(n51), .Q(n1768)
         );
  MUX21X1 U122 ( .IN1(\fifo[13][11] ), .IN2(data_in[11]), .S(n51), .Q(n1767)
         );
  MUX21X1 U123 ( .IN1(\fifo[13][12] ), .IN2(data_in[12]), .S(n51), .Q(n1766)
         );
  MUX21X1 U124 ( .IN1(\fifo[13][13] ), .IN2(data_in[13]), .S(n51), .Q(n1765)
         );
  MUX21X1 U125 ( .IN1(\fifo[13][14] ), .IN2(data_in[14]), .S(n51), .Q(n1764)
         );
  MUX21X1 U126 ( .IN1(\fifo[13][15] ), .IN2(data_in[15]), .S(n51), .Q(n1763)
         );
  MUX21X1 U127 ( .IN1(\fifo[13][16] ), .IN2(data_in[16]), .S(n51), .Q(n1762)
         );
  MUX21X1 U128 ( .IN1(\fifo[13][17] ), .IN2(data_in[17]), .S(n51), .Q(n1761)
         );
  MUX21X1 U129 ( .IN1(\fifo[13][18] ), .IN2(data_in[18]), .S(n51), .Q(n1760)
         );
  MUX21X1 U130 ( .IN1(\fifo[13][19] ), .IN2(data_in[19]), .S(n51), .Q(n1759)
         );
  MUX21X1 U131 ( .IN1(\fifo[13][20] ), .IN2(data_in[20]), .S(n51), .Q(n1758)
         );
  MUX21X1 U132 ( .IN1(\fifo[13][21] ), .IN2(data_in[21]), .S(n51), .Q(n1757)
         );
  MUX21X1 U133 ( .IN1(\fifo[13][22] ), .IN2(data_in[22]), .S(n51), .Q(n1756)
         );
  MUX21X1 U134 ( .IN1(\fifo[13][23] ), .IN2(data_in[23]), .S(n51), .Q(n1755)
         );
  MUX21X1 U135 ( .IN1(\fifo[13][24] ), .IN2(data_in[24]), .S(n51), .Q(n1754)
         );
  MUX21X1 U136 ( .IN1(\fifo[13][25] ), .IN2(data_in[25]), .S(n51), .Q(n1753)
         );
  MUX21X1 U137 ( .IN1(\fifo[13][26] ), .IN2(data_in[26]), .S(n51), .Q(n1752)
         );
  MUX21X1 U138 ( .IN1(\fifo[13][27] ), .IN2(data_in[27]), .S(n51), .Q(n1751)
         );
  MUX21X1 U139 ( .IN1(\fifo[13][28] ), .IN2(data_in[28]), .S(n51), .Q(n1750)
         );
  MUX21X1 U140 ( .IN1(\fifo[13][29] ), .IN2(data_in[29]), .S(n51), .Q(n1749)
         );
  MUX21X1 U141 ( .IN1(\fifo[13][30] ), .IN2(data_in[30]), .S(n51), .Q(n1748)
         );
  MUX21X1 U142 ( .IN1(\fifo[13][31] ), .IN2(data_in[31]), .S(n51), .Q(n1747)
         );
  AND2X1 U143 ( .IN1(n52), .IN2(n48), .Q(n51) );
  MUX21X1 U144 ( .IN1(\fifo[12][0] ), .IN2(data_in[0]), .S(n53), .Q(n1746) );
  MUX21X1 U145 ( .IN1(\fifo[12][1] ), .IN2(data_in[1]), .S(n53), .Q(n1745) );
  MUX21X1 U146 ( .IN1(\fifo[12][2] ), .IN2(data_in[2]), .S(n53), .Q(n1744) );
  MUX21X1 U147 ( .IN1(\fifo[12][3] ), .IN2(data_in[3]), .S(n53), .Q(n1743) );
  MUX21X1 U148 ( .IN1(\fifo[12][4] ), .IN2(data_in[4]), .S(n53), .Q(n1742) );
  MUX21X1 U149 ( .IN1(\fifo[12][5] ), .IN2(data_in[5]), .S(n53), .Q(n1741) );
  MUX21X1 U150 ( .IN1(\fifo[12][6] ), .IN2(data_in[6]), .S(n53), .Q(n1740) );
  MUX21X1 U151 ( .IN1(\fifo[12][7] ), .IN2(data_in[7]), .S(n53), .Q(n1739) );
  MUX21X1 U152 ( .IN1(\fifo[12][8] ), .IN2(data_in[8]), .S(n53), .Q(n1738) );
  MUX21X1 U153 ( .IN1(\fifo[12][9] ), .IN2(data_in[9]), .S(n53), .Q(n1737) );
  MUX21X1 U154 ( .IN1(\fifo[12][10] ), .IN2(data_in[10]), .S(n53), .Q(n1736)
         );
  MUX21X1 U155 ( .IN1(\fifo[12][11] ), .IN2(data_in[11]), .S(n53), .Q(n1735)
         );
  MUX21X1 U156 ( .IN1(\fifo[12][12] ), .IN2(data_in[12]), .S(n53), .Q(n1734)
         );
  MUX21X1 U157 ( .IN1(\fifo[12][13] ), .IN2(data_in[13]), .S(n53), .Q(n1733)
         );
  MUX21X1 U158 ( .IN1(\fifo[12][14] ), .IN2(data_in[14]), .S(n53), .Q(n1732)
         );
  MUX21X1 U159 ( .IN1(\fifo[12][15] ), .IN2(data_in[15]), .S(n53), .Q(n1731)
         );
  MUX21X1 U160 ( .IN1(\fifo[12][16] ), .IN2(data_in[16]), .S(n53), .Q(n1730)
         );
  MUX21X1 U161 ( .IN1(\fifo[12][17] ), .IN2(data_in[17]), .S(n53), .Q(n1729)
         );
  MUX21X1 U162 ( .IN1(\fifo[12][18] ), .IN2(data_in[18]), .S(n53), .Q(n1728)
         );
  MUX21X1 U163 ( .IN1(\fifo[12][19] ), .IN2(data_in[19]), .S(n53), .Q(n1727)
         );
  MUX21X1 U164 ( .IN1(\fifo[12][20] ), .IN2(data_in[20]), .S(n53), .Q(n1726)
         );
  MUX21X1 U165 ( .IN1(\fifo[12][21] ), .IN2(data_in[21]), .S(n53), .Q(n1725)
         );
  MUX21X1 U166 ( .IN1(\fifo[12][22] ), .IN2(data_in[22]), .S(n53), .Q(n1724)
         );
  MUX21X1 U167 ( .IN1(\fifo[12][23] ), .IN2(data_in[23]), .S(n53), .Q(n1723)
         );
  MUX21X1 U168 ( .IN1(\fifo[12][24] ), .IN2(data_in[24]), .S(n53), .Q(n1722)
         );
  MUX21X1 U169 ( .IN1(\fifo[12][25] ), .IN2(data_in[25]), .S(n53), .Q(n1721)
         );
  MUX21X1 U170 ( .IN1(\fifo[12][26] ), .IN2(data_in[26]), .S(n53), .Q(n1720)
         );
  MUX21X1 U171 ( .IN1(\fifo[12][27] ), .IN2(data_in[27]), .S(n53), .Q(n1719)
         );
  MUX21X1 U172 ( .IN1(\fifo[12][28] ), .IN2(data_in[28]), .S(n53), .Q(n1718)
         );
  MUX21X1 U173 ( .IN1(\fifo[12][29] ), .IN2(data_in[29]), .S(n53), .Q(n1717)
         );
  MUX21X1 U174 ( .IN1(\fifo[12][30] ), .IN2(data_in[30]), .S(n53), .Q(n1716)
         );
  MUX21X1 U175 ( .IN1(\fifo[12][31] ), .IN2(data_in[31]), .S(n53), .Q(n1715)
         );
  AND2X1 U176 ( .IN1(n54), .IN2(n48), .Q(n53) );
  NOR2X0 U177 ( .IN1(n3), .IN2(n1), .QN(n48) );
  MUX21X1 U178 ( .IN1(\fifo[11][0] ), .IN2(data_in[0]), .S(n55), .Q(n1714) );
  MUX21X1 U179 ( .IN1(\fifo[11][1] ), .IN2(data_in[1]), .S(n55), .Q(n1713) );
  MUX21X1 U180 ( .IN1(\fifo[11][2] ), .IN2(data_in[2]), .S(n55), .Q(n1712) );
  MUX21X1 U181 ( .IN1(\fifo[11][3] ), .IN2(data_in[3]), .S(n55), .Q(n1711) );
  MUX21X1 U182 ( .IN1(\fifo[11][4] ), .IN2(data_in[4]), .S(n55), .Q(n1710) );
  MUX21X1 U183 ( .IN1(\fifo[11][5] ), .IN2(data_in[5]), .S(n55), .Q(n1709) );
  MUX21X1 U184 ( .IN1(\fifo[11][6] ), .IN2(data_in[6]), .S(n55), .Q(n1708) );
  MUX21X1 U185 ( .IN1(\fifo[11][7] ), .IN2(data_in[7]), .S(n55), .Q(n1707) );
  MUX21X1 U186 ( .IN1(\fifo[11][8] ), .IN2(data_in[8]), .S(n55), .Q(n1706) );
  MUX21X1 U187 ( .IN1(\fifo[11][9] ), .IN2(data_in[9]), .S(n55), .Q(n1705) );
  MUX21X1 U188 ( .IN1(\fifo[11][10] ), .IN2(data_in[10]), .S(n55), .Q(n1704)
         );
  MUX21X1 U189 ( .IN1(\fifo[11][11] ), .IN2(data_in[11]), .S(n55), .Q(n1703)
         );
  MUX21X1 U190 ( .IN1(\fifo[11][12] ), .IN2(data_in[12]), .S(n55), .Q(n1702)
         );
  MUX21X1 U191 ( .IN1(\fifo[11][13] ), .IN2(data_in[13]), .S(n55), .Q(n1701)
         );
  MUX21X1 U192 ( .IN1(\fifo[11][14] ), .IN2(data_in[14]), .S(n55), .Q(n1700)
         );
  MUX21X1 U193 ( .IN1(\fifo[11][15] ), .IN2(data_in[15]), .S(n55), .Q(n1699)
         );
  MUX21X1 U194 ( .IN1(\fifo[11][16] ), .IN2(data_in[16]), .S(n55), .Q(n1698)
         );
  MUX21X1 U195 ( .IN1(\fifo[11][17] ), .IN2(data_in[17]), .S(n55), .Q(n1697)
         );
  MUX21X1 U196 ( .IN1(\fifo[11][18] ), .IN2(data_in[18]), .S(n55), .Q(n1696)
         );
  MUX21X1 U197 ( .IN1(\fifo[11][19] ), .IN2(data_in[19]), .S(n55), .Q(n1695)
         );
  MUX21X1 U198 ( .IN1(\fifo[11][20] ), .IN2(data_in[20]), .S(n55), .Q(n1694)
         );
  MUX21X1 U199 ( .IN1(\fifo[11][21] ), .IN2(data_in[21]), .S(n55), .Q(n1693)
         );
  MUX21X1 U200 ( .IN1(\fifo[11][22] ), .IN2(data_in[22]), .S(n55), .Q(n1692)
         );
  MUX21X1 U201 ( .IN1(\fifo[11][23] ), .IN2(data_in[23]), .S(n55), .Q(n1691)
         );
  MUX21X1 U202 ( .IN1(\fifo[11][24] ), .IN2(data_in[24]), .S(n55), .Q(n1690)
         );
  MUX21X1 U203 ( .IN1(\fifo[11][25] ), .IN2(data_in[25]), .S(n55), .Q(n1689)
         );
  MUX21X1 U204 ( .IN1(\fifo[11][26] ), .IN2(data_in[26]), .S(n55), .Q(n1688)
         );
  MUX21X1 U205 ( .IN1(\fifo[11][27] ), .IN2(data_in[27]), .S(n55), .Q(n1687)
         );
  MUX21X1 U206 ( .IN1(\fifo[11][28] ), .IN2(data_in[28]), .S(n55), .Q(n1686)
         );
  MUX21X1 U207 ( .IN1(\fifo[11][29] ), .IN2(data_in[29]), .S(n55), .Q(n1685)
         );
  MUX21X1 U208 ( .IN1(\fifo[11][30] ), .IN2(data_in[30]), .S(n55), .Q(n1684)
         );
  MUX21X1 U209 ( .IN1(\fifo[11][31] ), .IN2(data_in[31]), .S(n55), .Q(n1683)
         );
  AND2X1 U210 ( .IN1(n56), .IN2(n47), .Q(n55) );
  MUX21X1 U211 ( .IN1(\fifo[10][0] ), .IN2(data_in[0]), .S(n57), .Q(n1682) );
  MUX21X1 U212 ( .IN1(\fifo[10][1] ), .IN2(data_in[1]), .S(n57), .Q(n1681) );
  MUX21X1 U213 ( .IN1(\fifo[10][2] ), .IN2(data_in[2]), .S(n57), .Q(n1680) );
  MUX21X1 U214 ( .IN1(\fifo[10][3] ), .IN2(data_in[3]), .S(n57), .Q(n1679) );
  MUX21X1 U215 ( .IN1(\fifo[10][4] ), .IN2(data_in[4]), .S(n57), .Q(n1678) );
  MUX21X1 U216 ( .IN1(\fifo[10][5] ), .IN2(data_in[5]), .S(n57), .Q(n1677) );
  MUX21X1 U217 ( .IN1(\fifo[10][6] ), .IN2(data_in[6]), .S(n57), .Q(n1676) );
  MUX21X1 U218 ( .IN1(\fifo[10][7] ), .IN2(data_in[7]), .S(n57), .Q(n1675) );
  MUX21X1 U219 ( .IN1(\fifo[10][8] ), .IN2(data_in[8]), .S(n57), .Q(n1674) );
  MUX21X1 U220 ( .IN1(\fifo[10][9] ), .IN2(data_in[9]), .S(n57), .Q(n1673) );
  MUX21X1 U221 ( .IN1(\fifo[10][10] ), .IN2(data_in[10]), .S(n57), .Q(n1672)
         );
  MUX21X1 U222 ( .IN1(\fifo[10][11] ), .IN2(data_in[11]), .S(n57), .Q(n1671)
         );
  MUX21X1 U223 ( .IN1(\fifo[10][12] ), .IN2(data_in[12]), .S(n57), .Q(n1670)
         );
  MUX21X1 U224 ( .IN1(\fifo[10][13] ), .IN2(data_in[13]), .S(n57), .Q(n1669)
         );
  MUX21X1 U225 ( .IN1(\fifo[10][14] ), .IN2(data_in[14]), .S(n57), .Q(n1668)
         );
  MUX21X1 U226 ( .IN1(\fifo[10][15] ), .IN2(data_in[15]), .S(n57), .Q(n1667)
         );
  MUX21X1 U227 ( .IN1(\fifo[10][16] ), .IN2(data_in[16]), .S(n57), .Q(n1666)
         );
  MUX21X1 U228 ( .IN1(\fifo[10][17] ), .IN2(data_in[17]), .S(n57), .Q(n1665)
         );
  MUX21X1 U229 ( .IN1(\fifo[10][18] ), .IN2(data_in[18]), .S(n57), .Q(n1664)
         );
  MUX21X1 U230 ( .IN1(\fifo[10][19] ), .IN2(data_in[19]), .S(n57), .Q(n1663)
         );
  MUX21X1 U231 ( .IN1(\fifo[10][20] ), .IN2(data_in[20]), .S(n57), .Q(n1662)
         );
  MUX21X1 U232 ( .IN1(\fifo[10][21] ), .IN2(data_in[21]), .S(n57), .Q(n1661)
         );
  MUX21X1 U233 ( .IN1(\fifo[10][22] ), .IN2(data_in[22]), .S(n57), .Q(n1660)
         );
  MUX21X1 U234 ( .IN1(\fifo[10][23] ), .IN2(data_in[23]), .S(n57), .Q(n1659)
         );
  MUX21X1 U235 ( .IN1(\fifo[10][24] ), .IN2(data_in[24]), .S(n57), .Q(n1658)
         );
  MUX21X1 U236 ( .IN1(\fifo[10][25] ), .IN2(data_in[25]), .S(n57), .Q(n1657)
         );
  MUX21X1 U237 ( .IN1(\fifo[10][26] ), .IN2(data_in[26]), .S(n57), .Q(n1656)
         );
  MUX21X1 U238 ( .IN1(\fifo[10][27] ), .IN2(data_in[27]), .S(n57), .Q(n1655)
         );
  MUX21X1 U239 ( .IN1(\fifo[10][28] ), .IN2(data_in[28]), .S(n57), .Q(n1654)
         );
  MUX21X1 U240 ( .IN1(\fifo[10][29] ), .IN2(data_in[29]), .S(n57), .Q(n1653)
         );
  MUX21X1 U241 ( .IN1(\fifo[10][30] ), .IN2(data_in[30]), .S(n57), .Q(n1652)
         );
  MUX21X1 U242 ( .IN1(\fifo[10][31] ), .IN2(data_in[31]), .S(n57), .Q(n1651)
         );
  AND2X1 U243 ( .IN1(n56), .IN2(n50), .Q(n57) );
  MUX21X1 U244 ( .IN1(\fifo[9][0] ), .IN2(data_in[0]), .S(n58), .Q(n1650) );
  MUX21X1 U245 ( .IN1(\fifo[9][1] ), .IN2(data_in[1]), .S(n58), .Q(n1649) );
  MUX21X1 U246 ( .IN1(\fifo[9][2] ), .IN2(data_in[2]), .S(n58), .Q(n1648) );
  MUX21X1 U247 ( .IN1(\fifo[9][3] ), .IN2(data_in[3]), .S(n58), .Q(n1647) );
  MUX21X1 U248 ( .IN1(\fifo[9][4] ), .IN2(data_in[4]), .S(n58), .Q(n1646) );
  MUX21X1 U249 ( .IN1(\fifo[9][5] ), .IN2(data_in[5]), .S(n58), .Q(n1645) );
  MUX21X1 U250 ( .IN1(\fifo[9][6] ), .IN2(data_in[6]), .S(n58), .Q(n1644) );
  MUX21X1 U251 ( .IN1(\fifo[9][7] ), .IN2(data_in[7]), .S(n58), .Q(n1643) );
  MUX21X1 U252 ( .IN1(\fifo[9][8] ), .IN2(data_in[8]), .S(n58), .Q(n1642) );
  MUX21X1 U253 ( .IN1(\fifo[9][9] ), .IN2(data_in[9]), .S(n58), .Q(n1641) );
  MUX21X1 U254 ( .IN1(\fifo[9][10] ), .IN2(data_in[10]), .S(n58), .Q(n1640) );
  MUX21X1 U255 ( .IN1(\fifo[9][11] ), .IN2(data_in[11]), .S(n58), .Q(n1639) );
  MUX21X1 U256 ( .IN1(\fifo[9][12] ), .IN2(data_in[12]), .S(n58), .Q(n1638) );
  MUX21X1 U257 ( .IN1(\fifo[9][13] ), .IN2(data_in[13]), .S(n58), .Q(n1637) );
  MUX21X1 U258 ( .IN1(\fifo[9][14] ), .IN2(data_in[14]), .S(n58), .Q(n1636) );
  MUX21X1 U259 ( .IN1(\fifo[9][15] ), .IN2(data_in[15]), .S(n58), .Q(n1635) );
  MUX21X1 U260 ( .IN1(\fifo[9][16] ), .IN2(data_in[16]), .S(n58), .Q(n1634) );
  MUX21X1 U261 ( .IN1(\fifo[9][17] ), .IN2(data_in[17]), .S(n58), .Q(n1633) );
  MUX21X1 U262 ( .IN1(\fifo[9][18] ), .IN2(data_in[18]), .S(n58), .Q(n1632) );
  MUX21X1 U263 ( .IN1(\fifo[9][19] ), .IN2(data_in[19]), .S(n58), .Q(n1631) );
  MUX21X1 U264 ( .IN1(\fifo[9][20] ), .IN2(data_in[20]), .S(n58), .Q(n1630) );
  MUX21X1 U265 ( .IN1(\fifo[9][21] ), .IN2(data_in[21]), .S(n58), .Q(n1629) );
  MUX21X1 U266 ( .IN1(\fifo[9][22] ), .IN2(data_in[22]), .S(n58), .Q(n1628) );
  MUX21X1 U267 ( .IN1(\fifo[9][23] ), .IN2(data_in[23]), .S(n58), .Q(n1627) );
  MUX21X1 U268 ( .IN1(\fifo[9][24] ), .IN2(data_in[24]), .S(n58), .Q(n1626) );
  MUX21X1 U269 ( .IN1(\fifo[9][25] ), .IN2(data_in[25]), .S(n58), .Q(n1625) );
  MUX21X1 U270 ( .IN1(\fifo[9][26] ), .IN2(data_in[26]), .S(n58), .Q(n1624) );
  MUX21X1 U271 ( .IN1(\fifo[9][27] ), .IN2(data_in[27]), .S(n58), .Q(n1623) );
  MUX21X1 U272 ( .IN1(\fifo[9][28] ), .IN2(data_in[28]), .S(n58), .Q(n1622) );
  MUX21X1 U273 ( .IN1(\fifo[9][29] ), .IN2(data_in[29]), .S(n58), .Q(n1621) );
  MUX21X1 U274 ( .IN1(\fifo[9][30] ), .IN2(data_in[30]), .S(n58), .Q(n1620) );
  MUX21X1 U275 ( .IN1(\fifo[9][31] ), .IN2(data_in[31]), .S(n58), .Q(n1619) );
  AND2X1 U276 ( .IN1(n56), .IN2(n52), .Q(n58) );
  MUX21X1 U277 ( .IN1(\fifo[8][0] ), .IN2(data_in[0]), .S(n59), .Q(n1618) );
  MUX21X1 U278 ( .IN1(\fifo[8][1] ), .IN2(data_in[1]), .S(n59), .Q(n1617) );
  MUX21X1 U279 ( .IN1(\fifo[8][2] ), .IN2(data_in[2]), .S(n59), .Q(n1616) );
  MUX21X1 U280 ( .IN1(\fifo[8][3] ), .IN2(data_in[3]), .S(n59), .Q(n1615) );
  MUX21X1 U281 ( .IN1(\fifo[8][4] ), .IN2(data_in[4]), .S(n59), .Q(n1614) );
  MUX21X1 U282 ( .IN1(\fifo[8][5] ), .IN2(data_in[5]), .S(n59), .Q(n1613) );
  MUX21X1 U283 ( .IN1(\fifo[8][6] ), .IN2(data_in[6]), .S(n59), .Q(n1612) );
  MUX21X1 U284 ( .IN1(\fifo[8][7] ), .IN2(data_in[7]), .S(n59), .Q(n1611) );
  MUX21X1 U285 ( .IN1(\fifo[8][8] ), .IN2(data_in[8]), .S(n59), .Q(n1610) );
  MUX21X1 U286 ( .IN1(\fifo[8][9] ), .IN2(data_in[9]), .S(n59), .Q(n1609) );
  MUX21X1 U287 ( .IN1(\fifo[8][10] ), .IN2(data_in[10]), .S(n59), .Q(n1608) );
  MUX21X1 U288 ( .IN1(\fifo[8][11] ), .IN2(data_in[11]), .S(n59), .Q(n1607) );
  MUX21X1 U289 ( .IN1(\fifo[8][12] ), .IN2(data_in[12]), .S(n59), .Q(n1606) );
  MUX21X1 U290 ( .IN1(\fifo[8][13] ), .IN2(data_in[13]), .S(n59), .Q(n1605) );
  MUX21X1 U291 ( .IN1(\fifo[8][14] ), .IN2(data_in[14]), .S(n59), .Q(n1604) );
  MUX21X1 U292 ( .IN1(\fifo[8][15] ), .IN2(data_in[15]), .S(n59), .Q(n1603) );
  MUX21X1 U293 ( .IN1(\fifo[8][16] ), .IN2(data_in[16]), .S(n59), .Q(n1602) );
  MUX21X1 U294 ( .IN1(\fifo[8][17] ), .IN2(data_in[17]), .S(n59), .Q(n1601) );
  MUX21X1 U295 ( .IN1(\fifo[8][18] ), .IN2(data_in[18]), .S(n59), .Q(n1600) );
  MUX21X1 U296 ( .IN1(\fifo[8][19] ), .IN2(data_in[19]), .S(n59), .Q(n1599) );
  MUX21X1 U297 ( .IN1(\fifo[8][20] ), .IN2(data_in[20]), .S(n59), .Q(n1598) );
  MUX21X1 U298 ( .IN1(\fifo[8][21] ), .IN2(data_in[21]), .S(n59), .Q(n1597) );
  MUX21X1 U299 ( .IN1(\fifo[8][22] ), .IN2(data_in[22]), .S(n59), .Q(n1596) );
  MUX21X1 U300 ( .IN1(\fifo[8][23] ), .IN2(data_in[23]), .S(n59), .Q(n1595) );
  MUX21X1 U301 ( .IN1(\fifo[8][24] ), .IN2(data_in[24]), .S(n59), .Q(n1594) );
  MUX21X1 U302 ( .IN1(\fifo[8][25] ), .IN2(data_in[25]), .S(n59), .Q(n1593) );
  MUX21X1 U303 ( .IN1(\fifo[8][26] ), .IN2(data_in[26]), .S(n59), .Q(n1592) );
  MUX21X1 U304 ( .IN1(\fifo[8][27] ), .IN2(data_in[27]), .S(n59), .Q(n1591) );
  MUX21X1 U305 ( .IN1(\fifo[8][28] ), .IN2(data_in[28]), .S(n59), .Q(n1590) );
  MUX21X1 U306 ( .IN1(\fifo[8][29] ), .IN2(data_in[29]), .S(n59), .Q(n1589) );
  MUX21X1 U307 ( .IN1(\fifo[8][30] ), .IN2(data_in[30]), .S(n59), .Q(n1588) );
  MUX21X1 U308 ( .IN1(\fifo[8][31] ), .IN2(data_in[31]), .S(n59), .Q(n1587) );
  AND2X1 U309 ( .IN1(n56), .IN2(n54), .Q(n59) );
  MUX21X1 U310 ( .IN1(\fifo[7][0] ), .IN2(data_in[0]), .S(n60), .Q(n1586) );
  MUX21X1 U311 ( .IN1(\fifo[7][1] ), .IN2(data_in[1]), .S(n60), .Q(n1585) );
  MUX21X1 U312 ( .IN1(\fifo[7][2] ), .IN2(data_in[2]), .S(n60), .Q(n1584) );
  MUX21X1 U313 ( .IN1(\fifo[7][3] ), .IN2(data_in[3]), .S(n60), .Q(n1583) );
  MUX21X1 U314 ( .IN1(\fifo[7][4] ), .IN2(data_in[4]), .S(n60), .Q(n1582) );
  MUX21X1 U315 ( .IN1(\fifo[7][5] ), .IN2(data_in[5]), .S(n60), .Q(n1581) );
  MUX21X1 U316 ( .IN1(\fifo[7][6] ), .IN2(data_in[6]), .S(n60), .Q(n1580) );
  MUX21X1 U317 ( .IN1(\fifo[7][7] ), .IN2(data_in[7]), .S(n60), .Q(n1579) );
  MUX21X1 U318 ( .IN1(\fifo[7][8] ), .IN2(data_in[8]), .S(n60), .Q(n1578) );
  MUX21X1 U319 ( .IN1(\fifo[7][9] ), .IN2(data_in[9]), .S(n60), .Q(n1577) );
  MUX21X1 U320 ( .IN1(\fifo[7][10] ), .IN2(data_in[10]), .S(n60), .Q(n1576) );
  MUX21X1 U321 ( .IN1(\fifo[7][11] ), .IN2(data_in[11]), .S(n60), .Q(n1575) );
  MUX21X1 U322 ( .IN1(\fifo[7][12] ), .IN2(data_in[12]), .S(n60), .Q(n1574) );
  MUX21X1 U323 ( .IN1(\fifo[7][13] ), .IN2(data_in[13]), .S(n60), .Q(n1573) );
  MUX21X1 U324 ( .IN1(\fifo[7][14] ), .IN2(data_in[14]), .S(n60), .Q(n1572) );
  MUX21X1 U325 ( .IN1(\fifo[7][15] ), .IN2(data_in[15]), .S(n60), .Q(n1571) );
  MUX21X1 U326 ( .IN1(\fifo[7][16] ), .IN2(data_in[16]), .S(n60), .Q(n1570) );
  MUX21X1 U327 ( .IN1(\fifo[7][17] ), .IN2(data_in[17]), .S(n60), .Q(n1569) );
  MUX21X1 U328 ( .IN1(\fifo[7][18] ), .IN2(data_in[18]), .S(n60), .Q(n1568) );
  MUX21X1 U329 ( .IN1(\fifo[7][19] ), .IN2(data_in[19]), .S(n60), .Q(n1567) );
  MUX21X1 U330 ( .IN1(\fifo[7][20] ), .IN2(data_in[20]), .S(n60), .Q(n1566) );
  MUX21X1 U331 ( .IN1(\fifo[7][21] ), .IN2(data_in[21]), .S(n60), .Q(n1565) );
  MUX21X1 U332 ( .IN1(\fifo[7][22] ), .IN2(data_in[22]), .S(n60), .Q(n1564) );
  MUX21X1 U333 ( .IN1(\fifo[7][23] ), .IN2(data_in[23]), .S(n60), .Q(n1563) );
  MUX21X1 U334 ( .IN1(\fifo[7][24] ), .IN2(data_in[24]), .S(n60), .Q(n1562) );
  MUX21X1 U335 ( .IN1(\fifo[7][25] ), .IN2(data_in[25]), .S(n60), .Q(n1561) );
  MUX21X1 U336 ( .IN1(\fifo[7][26] ), .IN2(data_in[26]), .S(n60), .Q(n1560) );
  MUX21X1 U337 ( .IN1(\fifo[7][27] ), .IN2(data_in[27]), .S(n60), .Q(n1559) );
  MUX21X1 U338 ( .IN1(\fifo[7][28] ), .IN2(data_in[28]), .S(n60), .Q(n1558) );
  MUX21X1 U339 ( .IN1(\fifo[7][29] ), .IN2(data_in[29]), .S(n60), .Q(n1557) );
  MUX21X1 U340 ( .IN1(\fifo[7][30] ), .IN2(data_in[30]), .S(n60), .Q(n1556) );
  MUX21X1 U341 ( .IN1(\fifo[7][31] ), .IN2(data_in[31]), .S(n60), .Q(n1555) );
  MUX21X1 U342 ( .IN1(\fifo[6][0] ), .IN2(data_in[0]), .S(n61), .Q(n1554) );
  MUX21X1 U343 ( .IN1(\fifo[6][1] ), .IN2(data_in[1]), .S(n61), .Q(n1553) );
  MUX21X1 U344 ( .IN1(\fifo[6][2] ), .IN2(data_in[2]), .S(n61), .Q(n1552) );
  MUX21X1 U345 ( .IN1(\fifo[6][3] ), .IN2(data_in[3]), .S(n61), .Q(n1551) );
  MUX21X1 U346 ( .IN1(\fifo[6][4] ), .IN2(data_in[4]), .S(n61), .Q(n1550) );
  MUX21X1 U347 ( .IN1(\fifo[6][5] ), .IN2(data_in[5]), .S(n61), .Q(n1549) );
  MUX21X1 U348 ( .IN1(\fifo[6][6] ), .IN2(data_in[6]), .S(n61), .Q(n1548) );
  MUX21X1 U349 ( .IN1(\fifo[6][7] ), .IN2(data_in[7]), .S(n61), .Q(n1547) );
  MUX21X1 U350 ( .IN1(\fifo[6][8] ), .IN2(data_in[8]), .S(n61), .Q(n1546) );
  MUX21X1 U351 ( .IN1(\fifo[6][9] ), .IN2(data_in[9]), .S(n61), .Q(n1545) );
  MUX21X1 U352 ( .IN1(\fifo[6][10] ), .IN2(data_in[10]), .S(n61), .Q(n1544) );
  MUX21X1 U353 ( .IN1(\fifo[6][11] ), .IN2(data_in[11]), .S(n61), .Q(n1543) );
  MUX21X1 U354 ( .IN1(\fifo[6][12] ), .IN2(data_in[12]), .S(n61), .Q(n1542) );
  MUX21X1 U355 ( .IN1(\fifo[6][13] ), .IN2(data_in[13]), .S(n61), .Q(n1541) );
  MUX21X1 U356 ( .IN1(\fifo[6][14] ), .IN2(data_in[14]), .S(n61), .Q(n1540) );
  MUX21X1 U357 ( .IN1(\fifo[6][15] ), .IN2(data_in[15]), .S(n61), .Q(n1539) );
  MUX21X1 U358 ( .IN1(\fifo[6][16] ), .IN2(data_in[16]), .S(n61), .Q(n1538) );
  MUX21X1 U359 ( .IN1(\fifo[6][17] ), .IN2(data_in[17]), .S(n61), .Q(n1537) );
  MUX21X1 U360 ( .IN1(\fifo[6][18] ), .IN2(data_in[18]), .S(n61), .Q(n1536) );
  MUX21X1 U361 ( .IN1(\fifo[6][19] ), .IN2(data_in[19]), .S(n61), .Q(n1535) );
  MUX21X1 U362 ( .IN1(\fifo[6][20] ), .IN2(data_in[20]), .S(n61), .Q(n1534) );
  MUX21X1 U363 ( .IN1(\fifo[6][21] ), .IN2(data_in[21]), .S(n61), .Q(n1533) );
  MUX21X1 U364 ( .IN1(\fifo[6][22] ), .IN2(data_in[22]), .S(n61), .Q(n1532) );
  MUX21X1 U365 ( .IN1(\fifo[6][23] ), .IN2(data_in[23]), .S(n61), .Q(n1531) );
  MUX21X1 U366 ( .IN1(\fifo[6][24] ), .IN2(data_in[24]), .S(n61), .Q(n1530) );
  MUX21X1 U367 ( .IN1(\fifo[6][25] ), .IN2(data_in[25]), .S(n61), .Q(n1529) );
  MUX21X1 U368 ( .IN1(\fifo[6][26] ), .IN2(data_in[26]), .S(n61), .Q(n1528) );
  MUX21X1 U369 ( .IN1(\fifo[6][27] ), .IN2(data_in[27]), .S(n61), .Q(n1527) );
  MUX21X1 U370 ( .IN1(\fifo[6][28] ), .IN2(data_in[28]), .S(n61), .Q(n1526) );
  MUX21X1 U371 ( .IN1(\fifo[6][29] ), .IN2(data_in[29]), .S(n61), .Q(n1525) );
  MUX21X1 U372 ( .IN1(\fifo[6][30] ), .IN2(data_in[30]), .S(n61), .Q(n1524) );
  MUX21X1 U373 ( .IN1(\fifo[6][31] ), .IN2(data_in[31]), .S(n61), .Q(n1523) );
  AND2X1 U374 ( .IN1(n62), .IN2(n50), .Q(n61) );
  MUX21X1 U375 ( .IN1(\fifo[5][0] ), .IN2(data_in[0]), .S(n63), .Q(n1522) );
  MUX21X1 U376 ( .IN1(\fifo[5][1] ), .IN2(data_in[1]), .S(n63), .Q(n1521) );
  MUX21X1 U377 ( .IN1(\fifo[5][2] ), .IN2(data_in[2]), .S(n63), .Q(n1520) );
  MUX21X1 U378 ( .IN1(\fifo[5][3] ), .IN2(data_in[3]), .S(n63), .Q(n1519) );
  MUX21X1 U379 ( .IN1(\fifo[5][4] ), .IN2(data_in[4]), .S(n63), .Q(n1518) );
  MUX21X1 U380 ( .IN1(\fifo[5][5] ), .IN2(data_in[5]), .S(n63), .Q(n1517) );
  MUX21X1 U381 ( .IN1(\fifo[5][6] ), .IN2(data_in[6]), .S(n63), .Q(n1516) );
  MUX21X1 U382 ( .IN1(\fifo[5][7] ), .IN2(data_in[7]), .S(n63), .Q(n1515) );
  MUX21X1 U383 ( .IN1(\fifo[5][8] ), .IN2(data_in[8]), .S(n63), .Q(n1514) );
  MUX21X1 U384 ( .IN1(\fifo[5][9] ), .IN2(data_in[9]), .S(n63), .Q(n1513) );
  MUX21X1 U385 ( .IN1(\fifo[5][10] ), .IN2(data_in[10]), .S(n63), .Q(n1512) );
  MUX21X1 U386 ( .IN1(\fifo[5][11] ), .IN2(data_in[11]), .S(n63), .Q(n1511) );
  MUX21X1 U387 ( .IN1(\fifo[5][12] ), .IN2(data_in[12]), .S(n63), .Q(n1510) );
  MUX21X1 U388 ( .IN1(\fifo[5][13] ), .IN2(data_in[13]), .S(n63), .Q(n1509) );
  MUX21X1 U389 ( .IN1(\fifo[5][14] ), .IN2(data_in[14]), .S(n63), .Q(n1508) );
  MUX21X1 U390 ( .IN1(\fifo[5][15] ), .IN2(data_in[15]), .S(n63), .Q(n1507) );
  MUX21X1 U391 ( .IN1(\fifo[5][16] ), .IN2(data_in[16]), .S(n63), .Q(n1506) );
  MUX21X1 U392 ( .IN1(\fifo[5][17] ), .IN2(data_in[17]), .S(n63), .Q(n1505) );
  MUX21X1 U393 ( .IN1(\fifo[5][18] ), .IN2(data_in[18]), .S(n63), .Q(n1504) );
  MUX21X1 U394 ( .IN1(\fifo[5][19] ), .IN2(data_in[19]), .S(n63), .Q(n1503) );
  MUX21X1 U395 ( .IN1(\fifo[5][20] ), .IN2(data_in[20]), .S(n63), .Q(n1502) );
  MUX21X1 U396 ( .IN1(\fifo[5][21] ), .IN2(data_in[21]), .S(n63), .Q(n1501) );
  MUX21X1 U397 ( .IN1(\fifo[5][22] ), .IN2(data_in[22]), .S(n63), .Q(n1500) );
  MUX21X1 U398 ( .IN1(\fifo[5][23] ), .IN2(data_in[23]), .S(n63), .Q(n1499) );
  MUX21X1 U399 ( .IN1(\fifo[5][24] ), .IN2(data_in[24]), .S(n63), .Q(n1498) );
  MUX21X1 U400 ( .IN1(\fifo[5][25] ), .IN2(data_in[25]), .S(n63), .Q(n1497) );
  MUX21X1 U401 ( .IN1(\fifo[5][26] ), .IN2(data_in[26]), .S(n63), .Q(n1496) );
  MUX21X1 U402 ( .IN1(\fifo[5][27] ), .IN2(data_in[27]), .S(n63), .Q(n1495) );
  MUX21X1 U403 ( .IN1(\fifo[5][28] ), .IN2(data_in[28]), .S(n63), .Q(n1494) );
  MUX21X1 U404 ( .IN1(\fifo[5][29] ), .IN2(data_in[29]), .S(n63), .Q(n1493) );
  MUX21X1 U405 ( .IN1(\fifo[5][30] ), .IN2(data_in[30]), .S(n63), .Q(n1492) );
  MUX21X1 U406 ( .IN1(\fifo[5][31] ), .IN2(data_in[31]), .S(n63), .Q(n1491) );
  AND2X1 U407 ( .IN1(n62), .IN2(n52), .Q(n63) );
  MUX21X1 U408 ( .IN1(\fifo[4][0] ), .IN2(data_in[0]), .S(n64), .Q(n1490) );
  MUX21X1 U409 ( .IN1(\fifo[4][1] ), .IN2(data_in[1]), .S(n64), .Q(n1489) );
  MUX21X1 U410 ( .IN1(\fifo[4][2] ), .IN2(data_in[2]), .S(n64), .Q(n1488) );
  MUX21X1 U411 ( .IN1(\fifo[4][3] ), .IN2(data_in[3]), .S(n64), .Q(n1487) );
  MUX21X1 U412 ( .IN1(\fifo[4][4] ), .IN2(data_in[4]), .S(n64), .Q(n1486) );
  MUX21X1 U413 ( .IN1(\fifo[4][5] ), .IN2(data_in[5]), .S(n64), .Q(n1485) );
  MUX21X1 U414 ( .IN1(\fifo[4][6] ), .IN2(data_in[6]), .S(n64), .Q(n1484) );
  MUX21X1 U415 ( .IN1(\fifo[4][7] ), .IN2(data_in[7]), .S(n64), .Q(n1483) );
  MUX21X1 U416 ( .IN1(\fifo[4][8] ), .IN2(data_in[8]), .S(n64), .Q(n1482) );
  MUX21X1 U417 ( .IN1(\fifo[4][9] ), .IN2(data_in[9]), .S(n64), .Q(n1481) );
  MUX21X1 U418 ( .IN1(\fifo[4][10] ), .IN2(data_in[10]), .S(n64), .Q(n1480) );
  MUX21X1 U419 ( .IN1(\fifo[4][11] ), .IN2(data_in[11]), .S(n64), .Q(n1479) );
  MUX21X1 U420 ( .IN1(\fifo[4][12] ), .IN2(data_in[12]), .S(n64), .Q(n1478) );
  MUX21X1 U421 ( .IN1(\fifo[4][13] ), .IN2(data_in[13]), .S(n64), .Q(n1477) );
  MUX21X1 U422 ( .IN1(\fifo[4][14] ), .IN2(data_in[14]), .S(n64), .Q(n1476) );
  MUX21X1 U423 ( .IN1(\fifo[4][15] ), .IN2(data_in[15]), .S(n64), .Q(n1475) );
  MUX21X1 U424 ( .IN1(\fifo[4][16] ), .IN2(data_in[16]), .S(n64), .Q(n1474) );
  MUX21X1 U425 ( .IN1(\fifo[4][17] ), .IN2(data_in[17]), .S(n64), .Q(n1473) );
  MUX21X1 U426 ( .IN1(\fifo[4][18] ), .IN2(data_in[18]), .S(n64), .Q(n1472) );
  MUX21X1 U427 ( .IN1(\fifo[4][19] ), .IN2(data_in[19]), .S(n64), .Q(n1471) );
  MUX21X1 U428 ( .IN1(\fifo[4][20] ), .IN2(data_in[20]), .S(n64), .Q(n1470) );
  MUX21X1 U429 ( .IN1(\fifo[4][21] ), .IN2(data_in[21]), .S(n64), .Q(n1469) );
  MUX21X1 U430 ( .IN1(\fifo[4][22] ), .IN2(data_in[22]), .S(n64), .Q(n1468) );
  MUX21X1 U431 ( .IN1(\fifo[4][23] ), .IN2(data_in[23]), .S(n64), .Q(n1467) );
  MUX21X1 U432 ( .IN1(\fifo[4][24] ), .IN2(data_in[24]), .S(n64), .Q(n1466) );
  MUX21X1 U433 ( .IN1(\fifo[4][25] ), .IN2(data_in[25]), .S(n64), .Q(n1465) );
  MUX21X1 U434 ( .IN1(\fifo[4][26] ), .IN2(data_in[26]), .S(n64), .Q(n1464) );
  MUX21X1 U435 ( .IN1(\fifo[4][27] ), .IN2(data_in[27]), .S(n64), .Q(n1463) );
  MUX21X1 U436 ( .IN1(\fifo[4][28] ), .IN2(data_in[28]), .S(n64), .Q(n1462) );
  MUX21X1 U437 ( .IN1(\fifo[4][29] ), .IN2(data_in[29]), .S(n64), .Q(n1461) );
  MUX21X1 U438 ( .IN1(\fifo[4][30] ), .IN2(data_in[30]), .S(n64), .Q(n1460) );
  MUX21X1 U439 ( .IN1(\fifo[4][31] ), .IN2(data_in[31]), .S(n64), .Q(n1459) );
  AND2X1 U440 ( .IN1(n62), .IN2(n54), .Q(n64) );
  MUX21X1 U441 ( .IN1(\fifo[3][0] ), .IN2(data_in[0]), .S(n65), .Q(n1458) );
  MUX21X1 U442 ( .IN1(\fifo[3][1] ), .IN2(data_in[1]), .S(n65), .Q(n1457) );
  MUX21X1 U443 ( .IN1(\fifo[3][2] ), .IN2(data_in[2]), .S(n65), .Q(n1456) );
  MUX21X1 U444 ( .IN1(\fifo[3][3] ), .IN2(data_in[3]), .S(n65), .Q(n1455) );
  MUX21X1 U445 ( .IN1(\fifo[3][4] ), .IN2(data_in[4]), .S(n65), .Q(n1454) );
  MUX21X1 U446 ( .IN1(\fifo[3][5] ), .IN2(data_in[5]), .S(n65), .Q(n1453) );
  MUX21X1 U447 ( .IN1(\fifo[3][6] ), .IN2(data_in[6]), .S(n65), .Q(n1452) );
  MUX21X1 U448 ( .IN1(\fifo[3][7] ), .IN2(data_in[7]), .S(n65), .Q(n1451) );
  MUX21X1 U449 ( .IN1(\fifo[3][8] ), .IN2(data_in[8]), .S(n65), .Q(n1450) );
  MUX21X1 U450 ( .IN1(\fifo[3][9] ), .IN2(data_in[9]), .S(n65), .Q(n1449) );
  MUX21X1 U451 ( .IN1(\fifo[3][10] ), .IN2(data_in[10]), .S(n65), .Q(n1448) );
  MUX21X1 U452 ( .IN1(\fifo[3][11] ), .IN2(data_in[11]), .S(n65), .Q(n1447) );
  MUX21X1 U453 ( .IN1(\fifo[3][12] ), .IN2(data_in[12]), .S(n65), .Q(n1446) );
  MUX21X1 U454 ( .IN1(\fifo[3][13] ), .IN2(data_in[13]), .S(n65), .Q(n1445) );
  MUX21X1 U455 ( .IN1(\fifo[3][14] ), .IN2(data_in[14]), .S(n65), .Q(n1444) );
  MUX21X1 U456 ( .IN1(\fifo[3][15] ), .IN2(data_in[15]), .S(n65), .Q(n1443) );
  MUX21X1 U457 ( .IN1(\fifo[3][16] ), .IN2(data_in[16]), .S(n65), .Q(n1442) );
  MUX21X1 U458 ( .IN1(\fifo[3][17] ), .IN2(data_in[17]), .S(n65), .Q(n1441) );
  MUX21X1 U459 ( .IN1(\fifo[3][18] ), .IN2(data_in[18]), .S(n65), .Q(n1440) );
  MUX21X1 U460 ( .IN1(\fifo[3][19] ), .IN2(data_in[19]), .S(n65), .Q(n1439) );
  MUX21X1 U461 ( .IN1(\fifo[3][20] ), .IN2(data_in[20]), .S(n65), .Q(n1438) );
  MUX21X1 U462 ( .IN1(\fifo[3][21] ), .IN2(data_in[21]), .S(n65), .Q(n1437) );
  MUX21X1 U463 ( .IN1(\fifo[3][22] ), .IN2(data_in[22]), .S(n65), .Q(n1436) );
  MUX21X1 U464 ( .IN1(\fifo[3][23] ), .IN2(data_in[23]), .S(n65), .Q(n1435) );
  MUX21X1 U465 ( .IN1(\fifo[3][24] ), .IN2(data_in[24]), .S(n65), .Q(n1434) );
  MUX21X1 U466 ( .IN1(\fifo[3][25] ), .IN2(data_in[25]), .S(n65), .Q(n1433) );
  MUX21X1 U467 ( .IN1(\fifo[3][26] ), .IN2(data_in[26]), .S(n65), .Q(n1432) );
  MUX21X1 U468 ( .IN1(\fifo[3][27] ), .IN2(data_in[27]), .S(n65), .Q(n1431) );
  MUX21X1 U469 ( .IN1(\fifo[3][28] ), .IN2(data_in[28]), .S(n65), .Q(n1430) );
  MUX21X1 U470 ( .IN1(\fifo[3][29] ), .IN2(data_in[29]), .S(n65), .Q(n1429) );
  MUX21X1 U471 ( .IN1(\fifo[3][30] ), .IN2(data_in[30]), .S(n65), .Q(n1428) );
  MUX21X1 U472 ( .IN1(\fifo[3][31] ), .IN2(data_in[31]), .S(n65), .Q(n1427) );
  AND2X1 U473 ( .IN1(n66), .IN2(n47), .Q(n65) );
  MUX21X1 U474 ( .IN1(\fifo[2][0] ), .IN2(data_in[0]), .S(n67), .Q(n1426) );
  MUX21X1 U475 ( .IN1(\fifo[2][1] ), .IN2(data_in[1]), .S(n67), .Q(n1425) );
  MUX21X1 U476 ( .IN1(\fifo[2][2] ), .IN2(data_in[2]), .S(n67), .Q(n1424) );
  MUX21X1 U477 ( .IN1(\fifo[2][3] ), .IN2(data_in[3]), .S(n67), .Q(n1423) );
  MUX21X1 U478 ( .IN1(\fifo[2][4] ), .IN2(data_in[4]), .S(n67), .Q(n1422) );
  MUX21X1 U479 ( .IN1(\fifo[2][5] ), .IN2(data_in[5]), .S(n67), .Q(n1421) );
  MUX21X1 U480 ( .IN1(\fifo[2][6] ), .IN2(data_in[6]), .S(n67), .Q(n1420) );
  MUX21X1 U481 ( .IN1(\fifo[2][7] ), .IN2(data_in[7]), .S(n67), .Q(n1419) );
  MUX21X1 U482 ( .IN1(\fifo[2][8] ), .IN2(data_in[8]), .S(n67), .Q(n1418) );
  MUX21X1 U483 ( .IN1(\fifo[2][9] ), .IN2(data_in[9]), .S(n67), .Q(n1417) );
  MUX21X1 U484 ( .IN1(\fifo[2][10] ), .IN2(data_in[10]), .S(n67), .Q(n1416) );
  MUX21X1 U485 ( .IN1(\fifo[2][11] ), .IN2(data_in[11]), .S(n67), .Q(n1415) );
  MUX21X1 U486 ( .IN1(\fifo[2][12] ), .IN2(data_in[12]), .S(n67), .Q(n1414) );
  MUX21X1 U487 ( .IN1(\fifo[2][13] ), .IN2(data_in[13]), .S(n67), .Q(n1413) );
  MUX21X1 U488 ( .IN1(\fifo[2][14] ), .IN2(data_in[14]), .S(n67), .Q(n1412) );
  MUX21X1 U489 ( .IN1(\fifo[2][15] ), .IN2(data_in[15]), .S(n67), .Q(n1411) );
  MUX21X1 U490 ( .IN1(\fifo[2][16] ), .IN2(data_in[16]), .S(n67), .Q(n1410) );
  MUX21X1 U491 ( .IN1(\fifo[2][17] ), .IN2(data_in[17]), .S(n67), .Q(n1409) );
  MUX21X1 U492 ( .IN1(\fifo[2][18] ), .IN2(data_in[18]), .S(n67), .Q(n1408) );
  MUX21X1 U493 ( .IN1(\fifo[2][19] ), .IN2(data_in[19]), .S(n67), .Q(n1407) );
  MUX21X1 U494 ( .IN1(\fifo[2][20] ), .IN2(data_in[20]), .S(n67), .Q(n1406) );
  MUX21X1 U495 ( .IN1(\fifo[2][21] ), .IN2(data_in[21]), .S(n67), .Q(n1405) );
  MUX21X1 U496 ( .IN1(\fifo[2][22] ), .IN2(data_in[22]), .S(n67), .Q(n1404) );
  MUX21X1 U497 ( .IN1(\fifo[2][23] ), .IN2(data_in[23]), .S(n67), .Q(n1403) );
  MUX21X1 U498 ( .IN1(\fifo[2][24] ), .IN2(data_in[24]), .S(n67), .Q(n1402) );
  MUX21X1 U499 ( .IN1(\fifo[2][25] ), .IN2(data_in[25]), .S(n67), .Q(n1401) );
  MUX21X1 U500 ( .IN1(\fifo[2][26] ), .IN2(data_in[26]), .S(n67), .Q(n1400) );
  MUX21X1 U501 ( .IN1(\fifo[2][27] ), .IN2(data_in[27]), .S(n67), .Q(n1399) );
  MUX21X1 U502 ( .IN1(\fifo[2][28] ), .IN2(data_in[28]), .S(n67), .Q(n1398) );
  MUX21X1 U503 ( .IN1(\fifo[2][29] ), .IN2(data_in[29]), .S(n67), .Q(n1397) );
  MUX21X1 U504 ( .IN1(\fifo[2][30] ), .IN2(data_in[30]), .S(n67), .Q(n1396) );
  MUX21X1 U505 ( .IN1(\fifo[2][31] ), .IN2(data_in[31]), .S(n67), .Q(n1395) );
  AND2X1 U506 ( .IN1(n66), .IN2(n50), .Q(n67) );
  INVX0 U507 ( .INP(n68), .ZN(n50) );
  MUX21X1 U508 ( .IN1(\fifo[1][0] ), .IN2(data_in[0]), .S(n69), .Q(n1394) );
  MUX21X1 U509 ( .IN1(\fifo[1][1] ), .IN2(data_in[1]), .S(n69), .Q(n1393) );
  MUX21X1 U510 ( .IN1(\fifo[1][2] ), .IN2(data_in[2]), .S(n69), .Q(n1392) );
  MUX21X1 U511 ( .IN1(\fifo[1][3] ), .IN2(data_in[3]), .S(n69), .Q(n1391) );
  MUX21X1 U512 ( .IN1(\fifo[1][4] ), .IN2(data_in[4]), .S(n69), .Q(n1390) );
  MUX21X1 U513 ( .IN1(\fifo[1][5] ), .IN2(data_in[5]), .S(n69), .Q(n1389) );
  MUX21X1 U514 ( .IN1(\fifo[1][6] ), .IN2(data_in[6]), .S(n69), .Q(n1388) );
  MUX21X1 U515 ( .IN1(\fifo[1][7] ), .IN2(data_in[7]), .S(n69), .Q(n1387) );
  MUX21X1 U516 ( .IN1(\fifo[1][8] ), .IN2(data_in[8]), .S(n69), .Q(n1386) );
  MUX21X1 U517 ( .IN1(\fifo[1][9] ), .IN2(data_in[9]), .S(n69), .Q(n1385) );
  MUX21X1 U518 ( .IN1(\fifo[1][10] ), .IN2(data_in[10]), .S(n69), .Q(n1384) );
  MUX21X1 U519 ( .IN1(\fifo[1][11] ), .IN2(data_in[11]), .S(n69), .Q(n1383) );
  MUX21X1 U520 ( .IN1(\fifo[1][12] ), .IN2(data_in[12]), .S(n69), .Q(n1382) );
  MUX21X1 U521 ( .IN1(\fifo[1][13] ), .IN2(data_in[13]), .S(n69), .Q(n1381) );
  MUX21X1 U522 ( .IN1(\fifo[1][14] ), .IN2(data_in[14]), .S(n69), .Q(n1380) );
  MUX21X1 U523 ( .IN1(\fifo[1][15] ), .IN2(data_in[15]), .S(n69), .Q(n1379) );
  MUX21X1 U524 ( .IN1(\fifo[1][16] ), .IN2(data_in[16]), .S(n69), .Q(n1378) );
  MUX21X1 U525 ( .IN1(\fifo[1][17] ), .IN2(data_in[17]), .S(n69), .Q(n1377) );
  MUX21X1 U526 ( .IN1(\fifo[1][18] ), .IN2(data_in[18]), .S(n69), .Q(n1376) );
  MUX21X1 U527 ( .IN1(\fifo[1][19] ), .IN2(data_in[19]), .S(n69), .Q(n1375) );
  MUX21X1 U528 ( .IN1(\fifo[1][20] ), .IN2(data_in[20]), .S(n69), .Q(n1374) );
  MUX21X1 U529 ( .IN1(\fifo[1][21] ), .IN2(data_in[21]), .S(n69), .Q(n1373) );
  MUX21X1 U530 ( .IN1(\fifo[1][22] ), .IN2(data_in[22]), .S(n69), .Q(n1372) );
  MUX21X1 U531 ( .IN1(\fifo[1][23] ), .IN2(data_in[23]), .S(n69), .Q(n1371) );
  MUX21X1 U532 ( .IN1(\fifo[1][24] ), .IN2(data_in[24]), .S(n69), .Q(n1370) );
  MUX21X1 U533 ( .IN1(\fifo[1][25] ), .IN2(data_in[25]), .S(n69), .Q(n1369) );
  MUX21X1 U534 ( .IN1(\fifo[1][26] ), .IN2(data_in[26]), .S(n69), .Q(n1368) );
  MUX21X1 U535 ( .IN1(\fifo[1][27] ), .IN2(data_in[27]), .S(n69), .Q(n1367) );
  MUX21X1 U536 ( .IN1(\fifo[1][28] ), .IN2(data_in[28]), .S(n69), .Q(n1366) );
  MUX21X1 U537 ( .IN1(\fifo[1][29] ), .IN2(data_in[29]), .S(n69), .Q(n1365) );
  MUX21X1 U538 ( .IN1(\fifo[1][30] ), .IN2(data_in[30]), .S(n69), .Q(n1364) );
  MUX21X1 U539 ( .IN1(\fifo[1][31] ), .IN2(data_in[31]), .S(n69), .Q(n1363) );
  AND2X1 U540 ( .IN1(n66), .IN2(n52), .Q(n69) );
  INVX0 U541 ( .INP(n70), .ZN(n52) );
  MUX21X1 U542 ( .IN1(data_in[0]), .IN2(\fifo[0][0] ), .S(n71), .Q(n1362) );
  MUX21X1 U543 ( .IN1(data_in[1]), .IN2(\fifo[0][1] ), .S(n71), .Q(n1361) );
  MUX21X1 U544 ( .IN1(data_in[2]), .IN2(\fifo[0][2] ), .S(n71), .Q(n1360) );
  MUX21X1 U545 ( .IN1(data_in[3]), .IN2(\fifo[0][3] ), .S(n71), .Q(n1359) );
  MUX21X1 U546 ( .IN1(data_in[4]), .IN2(\fifo[0][4] ), .S(n71), .Q(n1358) );
  MUX21X1 U547 ( .IN1(data_in[5]), .IN2(\fifo[0][5] ), .S(n71), .Q(n1357) );
  MUX21X1 U548 ( .IN1(data_in[6]), .IN2(\fifo[0][6] ), .S(n71), .Q(n1356) );
  MUX21X1 U549 ( .IN1(data_in[7]), .IN2(\fifo[0][7] ), .S(n71), .Q(n1355) );
  MUX21X1 U550 ( .IN1(data_in[8]), .IN2(\fifo[0][8] ), .S(n71), .Q(n1354) );
  MUX21X1 U551 ( .IN1(data_in[9]), .IN2(\fifo[0][9] ), .S(n71), .Q(n1353) );
  MUX21X1 U552 ( .IN1(data_in[10]), .IN2(\fifo[0][10] ), .S(n71), .Q(n1352) );
  MUX21X1 U553 ( .IN1(data_in[11]), .IN2(\fifo[0][11] ), .S(n71), .Q(n1351) );
  MUX21X1 U554 ( .IN1(data_in[12]), .IN2(\fifo[0][12] ), .S(n71), .Q(n1350) );
  MUX21X1 U555 ( .IN1(data_in[13]), .IN2(\fifo[0][13] ), .S(n71), .Q(n1349) );
  MUX21X1 U556 ( .IN1(data_in[14]), .IN2(\fifo[0][14] ), .S(n71), .Q(n1348) );
  MUX21X1 U557 ( .IN1(data_in[15]), .IN2(\fifo[0][15] ), .S(n71), .Q(n1347) );
  MUX21X1 U558 ( .IN1(data_in[16]), .IN2(\fifo[0][16] ), .S(n71), .Q(n1346) );
  MUX21X1 U559 ( .IN1(data_in[17]), .IN2(\fifo[0][17] ), .S(n71), .Q(n1345) );
  MUX21X1 U560 ( .IN1(data_in[18]), .IN2(\fifo[0][18] ), .S(n71), .Q(n1344) );
  MUX21X1 U561 ( .IN1(data_in[19]), .IN2(\fifo[0][19] ), .S(n71), .Q(n1343) );
  MUX21X1 U562 ( .IN1(data_in[20]), .IN2(\fifo[0][20] ), .S(n71), .Q(n1342) );
  MUX21X1 U563 ( .IN1(data_in[21]), .IN2(\fifo[0][21] ), .S(n71), .Q(n1341) );
  MUX21X1 U564 ( .IN1(data_in[22]), .IN2(\fifo[0][22] ), .S(n71), .Q(n1340) );
  MUX21X1 U565 ( .IN1(data_in[23]), .IN2(\fifo[0][23] ), .S(n71), .Q(n1339) );
  MUX21X1 U566 ( .IN1(data_in[24]), .IN2(\fifo[0][24] ), .S(n71), .Q(n1338) );
  MUX21X1 U567 ( .IN1(data_in[25]), .IN2(\fifo[0][25] ), .S(n71), .Q(n1337) );
  MUX21X1 U568 ( .IN1(data_in[26]), .IN2(\fifo[0][26] ), .S(n71), .Q(n1336) );
  MUX21X1 U569 ( .IN1(data_in[27]), .IN2(\fifo[0][27] ), .S(n71), .Q(n1335) );
  MUX21X1 U570 ( .IN1(data_in[28]), .IN2(\fifo[0][28] ), .S(n71), .Q(n1334) );
  MUX21X1 U571 ( .IN1(data_in[29]), .IN2(\fifo[0][29] ), .S(n71), .Q(n1333) );
  MUX21X1 U572 ( .IN1(data_in[30]), .IN2(\fifo[0][30] ), .S(n71), .Q(n1332) );
  MUX21X1 U573 ( .IN1(data_in[31]), .IN2(\fifo[0][31] ), .S(n71), .Q(n1331) );
  AOI22X1 U574 ( .IN1(clear), .IN2(write), .IN3(n66), .IN4(n54), .QN(n71) );
  NOR2X0 U575 ( .IN1(n72), .IN2(write_pointer[1]), .QN(n54) );
  NOR2X0 U576 ( .IN1(write_pointer[3]), .IN2(write_pointer[2]), .QN(n66) );
  AO221X1 U577 ( .IN1(n56), .IN2(n73), .IN3(write_pointer[3]), .IN4(n74), 
        .IN5(n60), .Q(n1330) );
  AND2X1 U578 ( .IN1(n62), .IN2(n47), .Q(n60) );
  NOR2X0 U579 ( .IN1(n1), .IN2(write_pointer[3]), .QN(n62) );
  NOR2X0 U580 ( .IN1(n3), .IN2(write_pointer[2]), .QN(n56) );
  MUX21X1 U581 ( .IN1(n47), .IN2(n74), .S(write_pointer[2]), .Q(n1329) );
  NAND3X0 U582 ( .IN1(n75), .IN2(n72), .IN3(n76), .QN(n74) );
  NAND2X0 U583 ( .IN1(n73), .IN2(n4), .QN(n76) );
  INVX0 U584 ( .INP(n77), .ZN(n72) );
  AND3X1 U585 ( .IN1(write_pointer[0]), .IN2(n73), .IN3(write_pointer[1]), .Q(
        n47) );
  NAND3X0 U586 ( .IN1(n70), .IN2(n68), .IN3(n78), .QN(n1328) );
  NAND2X0 U587 ( .IN1(n79), .IN2(write_pointer[1]), .QN(n78) );
  NAND2X0 U588 ( .IN1(n77), .IN2(write_pointer[1]), .QN(n68) );
  NAND3X0 U589 ( .IN1(n73), .IN2(n4), .IN3(write_pointer[0]), .QN(n70) );
  INVX0 U590 ( .INP(n80), .ZN(n73) );
  AO221X1 U591 ( .IN1(n79), .IN2(write_pointer[0]), .IN3(clear), .IN4(write), 
        .IN5(n77), .Q(n1327) );
  NOR2X0 U592 ( .IN1(n80), .IN2(write_pointer[0]), .QN(n77) );
  INVX0 U593 ( .INP(n75), .ZN(n79) );
  NAND2X0 U594 ( .IN1(n80), .IN2(n81), .QN(n75) );
  NAND3X0 U595 ( .IN1(n45), .IN2(n81), .IN3(write), .QN(n80) );
  NAND3X0 U596 ( .IN1(n82), .IN2(cnt[4]), .IN3(n1311), .QN(n45) );
  AO22X1 U597 ( .IN1(n83), .IN2(N17), .IN3(n84), .IN4(n85), .Q(n1326) );
  NAND2X0 U598 ( .IN1(n86), .IN2(n87), .QN(n85) );
  MUX21X1 U599 ( .IN1(n83), .IN2(n88), .S(n1845), .Q(n1325) );
  NOR2X0 U600 ( .IN1(n89), .IN2(n90), .QN(n88) );
  AO21X1 U601 ( .IN1(n84), .IN2(n89), .IN3(n91), .Q(n83) );
  INVX0 U602 ( .INP(n92), .ZN(n89) );
  AO22X1 U603 ( .IN1(n91), .IN2(N15), .IN3(n84), .IN4(n93), .Q(n1324) );
  OR2X1 U604 ( .IN1(n94), .IN2(n95), .Q(n93) );
  AO21X1 U605 ( .IN1(\U3/U1/Z_0 ), .IN2(clear), .IN3(n96), .Q(n1323) );
  MUX21X1 U606 ( .IN1(n91), .IN2(n84), .S(n426), .Q(n96) );
  NOR2X0 U607 ( .IN1(n84), .IN2(clear), .QN(n91) );
  INVX0 U608 ( .INP(n90), .ZN(n84) );
  NAND3X0 U609 ( .IN1(n97), .IN2(n81), .IN3(\U3/U1/Z_0 ), .QN(n90) );
  AO22X1 U610 ( .IN1(n98), .IN2(cnt[4]), .IN3(n99), .IN4(n100), .Q(n1322) );
  XOR3X1 U611 ( .IN1(n1848), .IN2(\U3/U1/Z_0 ), .IN3(n101), .Q(n100) );
  OA22X1 U612 ( .IN1(n1313), .IN2(n102), .IN3(n103), .IN4(n104), .Q(n101) );
  NOR2X0 U613 ( .IN1(\U3/U1/Z_0 ), .IN2(n105), .QN(n102) );
  AO22X1 U614 ( .IN1(n98), .IN2(cnt[3]), .IN3(n99), .IN4(n106), .Q(n1321) );
  XOR3X1 U615 ( .IN1(n1313), .IN2(\U3/U1/Z_0 ), .IN3(n103), .Q(n106) );
  INVX0 U616 ( .INP(n105), .ZN(n103) );
  AO22X1 U617 ( .IN1(\U3/U1/Z_0 ), .IN2(n107), .IN3(n108), .IN4(cnt[2]), .Q(
        n105) );
  OR2X1 U618 ( .IN1(n107), .IN2(\U3/U1/Z_0 ), .Q(n108) );
  AO22X1 U619 ( .IN1(n98), .IN2(cnt[2]), .IN3(n99), .IN4(n109), .Q(n1320) );
  XOR3X1 U620 ( .IN1(\U3/U1/Z_0 ), .IN2(cnt[2]), .IN3(n107), .Q(n109) );
  AO21X1 U621 ( .IN1(\U3/U1/Z_0 ), .IN2(n110), .IN3(n111), .Q(n107) );
  NAND2X0 U622 ( .IN1(n1311), .IN2(n1847), .QN(n110) );
  AO22X1 U623 ( .IN1(n98), .IN2(cnt[1]), .IN3(n99), .IN4(n112), .Q(n1319) );
  AO21X1 U624 ( .IN1(n111), .IN2(\U3/U1/Z_0 ), .IN3(n113), .Q(n112) );
  MUX21X1 U625 ( .IN1(n114), .IN2(n115), .S(n1847), .Q(n113) );
  XOR2X1 U626 ( .IN1(cnt[0]), .IN2(\U3/U1/Z_0 ), .Q(n115) );
  NOR2X0 U627 ( .IN1(\U3/U1/Z_0 ), .IN2(cnt[0]), .QN(n114) );
  AO21X1 U628 ( .IN1(clear), .IN2(n116), .IN3(n117), .Q(n1318) );
  MUX21X1 U629 ( .IN1(n98), .IN2(n99), .S(n1311), .Q(n117) );
  NOR2X0 U630 ( .IN1(n99), .IN2(clear), .QN(n98) );
  AND2X1 U631 ( .IN1(n116), .IN2(n81), .Q(n99) );
  INVX0 U632 ( .INP(clear), .ZN(n81) );
  XNOR2X1 U633 ( .IN1(write), .IN2(n104), .Q(n116) );
  INVX0 U634 ( .INP(\U3/U1/Z_0 ), .ZN(n104) );
  INVX0 U635 ( .INP(n97), .ZN(empty) );
  NAND3X0 U636 ( .IN1(n1311), .IN2(n82), .IN3(n1848), .QN(n97) );
  AND3X1 U637 ( .IN1(cnt[2]), .IN2(cnt[3]), .IN3(n111), .Q(almost_full) );
  NOR2X0 U638 ( .IN1(n1311), .IN2(n1847), .QN(n111) );
  AND3X1 U639 ( .IN1(n1848), .IN2(cnt[0]), .IN3(n82), .Q(almost_empty) );
  AND3X1 U640 ( .IN1(n1313), .IN2(n1312), .IN3(n1847), .Q(n82) );
  MUX21X1 U641 ( .IN1(n118), .IN2(\fifo[0][31] ), .S(clear), .Q(N155) );
  NAND4X0 U642 ( .IN1(n119), .IN2(n120), .IN3(n121), .IN4(n122), .QN(n118) );
  OA221X1 U643 ( .IN1(n1156), .IN2(n123), .IN3(n1935), .IN4(n124), .IN5(n125), 
        .Q(n122) );
  OA22X1 U644 ( .IN1(n1028), .IN2(n126), .IN3(n1913), .IN4(n127), .Q(n125) );
  OA221X1 U645 ( .IN1(n964), .IN2(n128), .IN3(n1092), .IN4(n129), .IN5(n130), 
        .Q(n121) );
  OA22X1 U646 ( .IN1(n1849), .IN2(n131), .IN3(n1220), .IN4(n132), .Q(n130) );
  OA221X1 U647 ( .IN1(n932), .IN2(n133), .IN3(n1060), .IN4(n134), .IN5(n135), 
        .Q(n120) );
  OA22X1 U648 ( .IN1(n1284), .IN2(n136), .IN3(n1188), .IN4(n137), .Q(n135) );
  OA221X1 U649 ( .IN1(n1252), .IN2(n138), .IN3(n1881), .IN4(n139), .IN5(n140), 
        .Q(n119) );
  OA22X1 U650 ( .IN1(n1124), .IN2(n141), .IN3(n996), .IN4(n86), .Q(n140) );
  MUX21X1 U651 ( .IN1(n142), .IN2(\fifo[0][30] ), .S(clear), .Q(N154) );
  NAND4X0 U652 ( .IN1(n143), .IN2(n144), .IN3(n145), .IN4(n146), .QN(n142) );
  OA221X1 U653 ( .IN1(n1157), .IN2(n123), .IN3(n1936), .IN4(n124), .IN5(n147), 
        .Q(n146) );
  OA22X1 U654 ( .IN1(n1029), .IN2(n126), .IN3(n1914), .IN4(n127), .Q(n147) );
  OA221X1 U655 ( .IN1(n965), .IN2(n128), .IN3(n1093), .IN4(n129), .IN5(n148), 
        .Q(n145) );
  OA22X1 U656 ( .IN1(n1850), .IN2(n131), .IN3(n1221), .IN4(n132), .Q(n148) );
  OA221X1 U657 ( .IN1(n933), .IN2(n133), .IN3(n1061), .IN4(n134), .IN5(n149), 
        .Q(n144) );
  OA22X1 U658 ( .IN1(n1285), .IN2(n136), .IN3(n1189), .IN4(n137), .Q(n149) );
  OA221X1 U659 ( .IN1(n1253), .IN2(n138), .IN3(n1882), .IN4(n139), .IN5(n150), 
        .Q(n143) );
  OA22X1 U660 ( .IN1(n1125), .IN2(n141), .IN3(n997), .IN4(n86), .Q(n150) );
  MUX21X1 U661 ( .IN1(n151), .IN2(\fifo[0][29] ), .S(clear), .Q(N153) );
  NAND4X0 U662 ( .IN1(n152), .IN2(n153), .IN3(n154), .IN4(n155), .QN(n151) );
  OA221X1 U663 ( .IN1(n1158), .IN2(n123), .IN3(n1937), .IN4(n124), .IN5(n156), 
        .Q(n155) );
  OA22X1 U664 ( .IN1(n1030), .IN2(n126), .IN3(n1915), .IN4(n127), .Q(n156) );
  OA221X1 U665 ( .IN1(n966), .IN2(n128), .IN3(n1094), .IN4(n129), .IN5(n157), 
        .Q(n154) );
  OA22X1 U666 ( .IN1(n1851), .IN2(n131), .IN3(n1222), .IN4(n132), .Q(n157) );
  OA221X1 U667 ( .IN1(n934), .IN2(n133), .IN3(n1062), .IN4(n134), .IN5(n158), 
        .Q(n153) );
  OA22X1 U668 ( .IN1(n1286), .IN2(n136), .IN3(n1190), .IN4(n137), .Q(n158) );
  OA221X1 U669 ( .IN1(n1254), .IN2(n138), .IN3(n1883), .IN4(n139), .IN5(n159), 
        .Q(n152) );
  OA22X1 U670 ( .IN1(n1126), .IN2(n141), .IN3(n998), .IN4(n86), .Q(n159) );
  MUX21X1 U671 ( .IN1(n160), .IN2(\fifo[0][28] ), .S(clear), .Q(N152) );
  NAND4X0 U672 ( .IN1(n161), .IN2(n162), .IN3(n163), .IN4(n164), .QN(n160) );
  OA221X1 U673 ( .IN1(n1159), .IN2(n123), .IN3(n1938), .IN4(n124), .IN5(n165), 
        .Q(n164) );
  OA22X1 U674 ( .IN1(n1031), .IN2(n126), .IN3(n1916), .IN4(n127), .Q(n165) );
  OA221X1 U675 ( .IN1(n967), .IN2(n128), .IN3(n1095), .IN4(n129), .IN5(n166), 
        .Q(n163) );
  OA22X1 U676 ( .IN1(n1852), .IN2(n131), .IN3(n1223), .IN4(n132), .Q(n166) );
  OA221X1 U677 ( .IN1(n935), .IN2(n133), .IN3(n1063), .IN4(n134), .IN5(n167), 
        .Q(n162) );
  OA22X1 U678 ( .IN1(n1287), .IN2(n136), .IN3(n1191), .IN4(n137), .Q(n167) );
  OA221X1 U679 ( .IN1(n1255), .IN2(n138), .IN3(n1884), .IN4(n139), .IN5(n168), 
        .Q(n161) );
  OA22X1 U680 ( .IN1(n1127), .IN2(n141), .IN3(n999), .IN4(n86), .Q(n168) );
  MUX21X1 U681 ( .IN1(n169), .IN2(\fifo[0][27] ), .S(clear), .Q(N151) );
  NAND4X0 U682 ( .IN1(n170), .IN2(n171), .IN3(n172), .IN4(n173), .QN(n169) );
  OA221X1 U683 ( .IN1(n1160), .IN2(n123), .IN3(n1939), .IN4(n124), .IN5(n174), 
        .Q(n173) );
  OA22X1 U684 ( .IN1(n1032), .IN2(n126), .IN3(n1917), .IN4(n127), .Q(n174) );
  OA221X1 U685 ( .IN1(n968), .IN2(n128), .IN3(n1096), .IN4(n129), .IN5(n175), 
        .Q(n172) );
  OA22X1 U686 ( .IN1(n1853), .IN2(n131), .IN3(n1224), .IN4(n132), .Q(n175) );
  OA221X1 U687 ( .IN1(n936), .IN2(n133), .IN3(n1064), .IN4(n134), .IN5(n176), 
        .Q(n171) );
  OA22X1 U688 ( .IN1(n1288), .IN2(n136), .IN3(n1192), .IN4(n137), .Q(n176) );
  OA221X1 U689 ( .IN1(n1256), .IN2(n138), .IN3(n1885), .IN4(n139), .IN5(n177), 
        .Q(n170) );
  OA22X1 U690 ( .IN1(n1128), .IN2(n141), .IN3(n1000), .IN4(n86), .Q(n177) );
  MUX21X1 U691 ( .IN1(n178), .IN2(\fifo[0][26] ), .S(clear), .Q(N150) );
  NAND4X0 U692 ( .IN1(n179), .IN2(n180), .IN3(n181), .IN4(n182), .QN(n178) );
  OA221X1 U693 ( .IN1(n1161), .IN2(n123), .IN3(n1940), .IN4(n124), .IN5(n183), 
        .Q(n182) );
  OA22X1 U694 ( .IN1(n1033), .IN2(n126), .IN3(n1918), .IN4(n127), .Q(n183) );
  OA221X1 U695 ( .IN1(n969), .IN2(n128), .IN3(n1097), .IN4(n129), .IN5(n184), 
        .Q(n181) );
  OA22X1 U696 ( .IN1(n1854), .IN2(n131), .IN3(n1225), .IN4(n132), .Q(n184) );
  OA221X1 U697 ( .IN1(n937), .IN2(n133), .IN3(n1065), .IN4(n134), .IN5(n185), 
        .Q(n180) );
  OA22X1 U698 ( .IN1(n1289), .IN2(n136), .IN3(n1193), .IN4(n137), .Q(n185) );
  OA221X1 U699 ( .IN1(n1257), .IN2(n138), .IN3(n1886), .IN4(n139), .IN5(n186), 
        .Q(n179) );
  OA22X1 U700 ( .IN1(n1129), .IN2(n141), .IN3(n1001), .IN4(n86), .Q(n186) );
  MUX21X1 U701 ( .IN1(n187), .IN2(\fifo[0][25] ), .S(clear), .Q(N149) );
  NAND4X0 U702 ( .IN1(n188), .IN2(n189), .IN3(n190), .IN4(n191), .QN(n187) );
  OA221X1 U703 ( .IN1(n1162), .IN2(n123), .IN3(n1941), .IN4(n124), .IN5(n192), 
        .Q(n191) );
  OA22X1 U704 ( .IN1(n1034), .IN2(n126), .IN3(n1919), .IN4(n127), .Q(n192) );
  OA221X1 U705 ( .IN1(n970), .IN2(n128), .IN3(n1098), .IN4(n129), .IN5(n193), 
        .Q(n190) );
  OA22X1 U706 ( .IN1(n1855), .IN2(n131), .IN3(n1226), .IN4(n132), .Q(n193) );
  OA221X1 U707 ( .IN1(n938), .IN2(n133), .IN3(n1066), .IN4(n134), .IN5(n194), 
        .Q(n189) );
  OA22X1 U708 ( .IN1(n1290), .IN2(n136), .IN3(n1194), .IN4(n137), .Q(n194) );
  OA221X1 U709 ( .IN1(n1258), .IN2(n138), .IN3(n1887), .IN4(n139), .IN5(n195), 
        .Q(n188) );
  OA22X1 U710 ( .IN1(n1130), .IN2(n141), .IN3(n1002), .IN4(n86), .Q(n195) );
  MUX21X1 U711 ( .IN1(n196), .IN2(\fifo[0][24] ), .S(clear), .Q(N148) );
  NAND4X0 U712 ( .IN1(n197), .IN2(n198), .IN3(n199), .IN4(n200), .QN(n196) );
  OA221X1 U713 ( .IN1(n1163), .IN2(n123), .IN3(n1942), .IN4(n124), .IN5(n201), 
        .Q(n200) );
  OA22X1 U714 ( .IN1(n1035), .IN2(n126), .IN3(n1920), .IN4(n127), .Q(n201) );
  OA221X1 U715 ( .IN1(n971), .IN2(n128), .IN3(n1099), .IN4(n129), .IN5(n202), 
        .Q(n199) );
  OA22X1 U716 ( .IN1(n1856), .IN2(n131), .IN3(n1227), .IN4(n132), .Q(n202) );
  OA221X1 U717 ( .IN1(n939), .IN2(n133), .IN3(n1067), .IN4(n134), .IN5(n203), 
        .Q(n198) );
  OA22X1 U718 ( .IN1(n1291), .IN2(n136), .IN3(n1195), .IN4(n137), .Q(n203) );
  OA221X1 U719 ( .IN1(n1259), .IN2(n138), .IN3(n1888), .IN4(n139), .IN5(n204), 
        .Q(n197) );
  OA22X1 U720 ( .IN1(n1131), .IN2(n141), .IN3(n1003), .IN4(n86), .Q(n204) );
  MUX21X1 U721 ( .IN1(n205), .IN2(\fifo[0][23] ), .S(clear), .Q(N147) );
  NAND4X0 U722 ( .IN1(n206), .IN2(n207), .IN3(n208), .IN4(n209), .QN(n205) );
  OA221X1 U723 ( .IN1(n1164), .IN2(n123), .IN3(n1943), .IN4(n124), .IN5(n210), 
        .Q(n209) );
  OA22X1 U724 ( .IN1(n1036), .IN2(n126), .IN3(n1921), .IN4(n127), .Q(n210) );
  OA221X1 U725 ( .IN1(n972), .IN2(n128), .IN3(n1100), .IN4(n129), .IN5(n211), 
        .Q(n208) );
  OA22X1 U726 ( .IN1(n1857), .IN2(n131), .IN3(n1228), .IN4(n132), .Q(n211) );
  OA221X1 U727 ( .IN1(n940), .IN2(n133), .IN3(n1068), .IN4(n134), .IN5(n212), 
        .Q(n207) );
  OA22X1 U728 ( .IN1(n1292), .IN2(n136), .IN3(n1196), .IN4(n137), .Q(n212) );
  OA221X1 U729 ( .IN1(n1260), .IN2(n138), .IN3(n1889), .IN4(n139), .IN5(n213), 
        .Q(n206) );
  OA22X1 U730 ( .IN1(n1132), .IN2(n141), .IN3(n1004), .IN4(n86), .Q(n213) );
  MUX21X1 U731 ( .IN1(n214), .IN2(\fifo[0][22] ), .S(clear), .Q(N146) );
  NAND4X0 U732 ( .IN1(n215), .IN2(n216), .IN3(n217), .IN4(n218), .QN(n214) );
  OA221X1 U733 ( .IN1(n1165), .IN2(n123), .IN3(n1944), .IN4(n124), .IN5(n219), 
        .Q(n218) );
  OA22X1 U734 ( .IN1(n1037), .IN2(n126), .IN3(n1922), .IN4(n127), .Q(n219) );
  OA221X1 U735 ( .IN1(n973), .IN2(n128), .IN3(n1101), .IN4(n129), .IN5(n220), 
        .Q(n217) );
  OA22X1 U736 ( .IN1(n1858), .IN2(n131), .IN3(n1229), .IN4(n132), .Q(n220) );
  OA221X1 U737 ( .IN1(n941), .IN2(n133), .IN3(n1069), .IN4(n134), .IN5(n221), 
        .Q(n216) );
  OA22X1 U738 ( .IN1(n1293), .IN2(n136), .IN3(n1197), .IN4(n137), .Q(n221) );
  OA221X1 U739 ( .IN1(n1261), .IN2(n138), .IN3(n1890), .IN4(n139), .IN5(n222), 
        .Q(n215) );
  OA22X1 U740 ( .IN1(n1133), .IN2(n141), .IN3(n1005), .IN4(n86), .Q(n222) );
  MUX21X1 U741 ( .IN1(n223), .IN2(\fifo[0][21] ), .S(clear), .Q(N145) );
  NAND4X0 U742 ( .IN1(n224), .IN2(n225), .IN3(n226), .IN4(n227), .QN(n223) );
  OA221X1 U743 ( .IN1(n1166), .IN2(n123), .IN3(n1945), .IN4(n124), .IN5(n228), 
        .Q(n227) );
  OA22X1 U744 ( .IN1(n1038), .IN2(n126), .IN3(n1923), .IN4(n127), .Q(n228) );
  OA221X1 U745 ( .IN1(n974), .IN2(n128), .IN3(n1102), .IN4(n129), .IN5(n229), 
        .Q(n226) );
  OA22X1 U746 ( .IN1(n1859), .IN2(n131), .IN3(n1230), .IN4(n132), .Q(n229) );
  OA221X1 U747 ( .IN1(n942), .IN2(n133), .IN3(n1070), .IN4(n134), .IN5(n230), 
        .Q(n225) );
  OA22X1 U748 ( .IN1(n1294), .IN2(n136), .IN3(n1198), .IN4(n137), .Q(n230) );
  OA221X1 U749 ( .IN1(n1262), .IN2(n138), .IN3(n1891), .IN4(n139), .IN5(n231), 
        .Q(n224) );
  OA22X1 U750 ( .IN1(n1134), .IN2(n141), .IN3(n1006), .IN4(n86), .Q(n231) );
  MUX21X1 U751 ( .IN1(n232), .IN2(\fifo[0][20] ), .S(clear), .Q(N144) );
  NAND4X0 U752 ( .IN1(n233), .IN2(n234), .IN3(n235), .IN4(n236), .QN(n232) );
  OA221X1 U753 ( .IN1(n1167), .IN2(n123), .IN3(n1946), .IN4(n124), .IN5(n237), 
        .Q(n236) );
  OA22X1 U754 ( .IN1(n1039), .IN2(n126), .IN3(n1924), .IN4(n127), .Q(n237) );
  OA221X1 U755 ( .IN1(n975), .IN2(n128), .IN3(n1103), .IN4(n129), .IN5(n238), 
        .Q(n235) );
  OA22X1 U756 ( .IN1(n1860), .IN2(n131), .IN3(n1231), .IN4(n132), .Q(n238) );
  OA221X1 U757 ( .IN1(n943), .IN2(n133), .IN3(n1071), .IN4(n134), .IN5(n239), 
        .Q(n234) );
  OA22X1 U758 ( .IN1(n1295), .IN2(n136), .IN3(n1199), .IN4(n137), .Q(n239) );
  OA221X1 U759 ( .IN1(n1263), .IN2(n138), .IN3(n1892), .IN4(n139), .IN5(n240), 
        .Q(n233) );
  OA22X1 U760 ( .IN1(n1135), .IN2(n141), .IN3(n1007), .IN4(n86), .Q(n240) );
  MUX21X1 U761 ( .IN1(n241), .IN2(\fifo[0][19] ), .S(clear), .Q(N143) );
  NAND4X0 U762 ( .IN1(n242), .IN2(n243), .IN3(n244), .IN4(n245), .QN(n241) );
  OA221X1 U763 ( .IN1(n1168), .IN2(n123), .IN3(n1947), .IN4(n124), .IN5(n246), 
        .Q(n245) );
  OA22X1 U764 ( .IN1(n1040), .IN2(n126), .IN3(n1925), .IN4(n127), .Q(n246) );
  OA221X1 U765 ( .IN1(n976), .IN2(n128), .IN3(n1104), .IN4(n129), .IN5(n247), 
        .Q(n244) );
  OA22X1 U766 ( .IN1(n1861), .IN2(n131), .IN3(n1232), .IN4(n132), .Q(n247) );
  OA221X1 U767 ( .IN1(n944), .IN2(n133), .IN3(n1072), .IN4(n134), .IN5(n248), 
        .Q(n243) );
  OA22X1 U768 ( .IN1(n1296), .IN2(n136), .IN3(n1200), .IN4(n137), .Q(n248) );
  OA221X1 U769 ( .IN1(n1264), .IN2(n138), .IN3(n1893), .IN4(n139), .IN5(n249), 
        .Q(n242) );
  OA22X1 U770 ( .IN1(n1136), .IN2(n141), .IN3(n1008), .IN4(n86), .Q(n249) );
  MUX21X1 U771 ( .IN1(n250), .IN2(\fifo[0][18] ), .S(clear), .Q(N142) );
  NAND4X0 U772 ( .IN1(n251), .IN2(n252), .IN3(n253), .IN4(n254), .QN(n250) );
  OA221X1 U773 ( .IN1(n1169), .IN2(n123), .IN3(n1948), .IN4(n124), .IN5(n255), 
        .Q(n254) );
  OA22X1 U774 ( .IN1(n1041), .IN2(n126), .IN3(n1926), .IN4(n127), .Q(n255) );
  OA221X1 U775 ( .IN1(n977), .IN2(n128), .IN3(n1105), .IN4(n129), .IN5(n256), 
        .Q(n253) );
  OA22X1 U776 ( .IN1(n1862), .IN2(n131), .IN3(n1233), .IN4(n132), .Q(n256) );
  OA221X1 U777 ( .IN1(n945), .IN2(n133), .IN3(n1073), .IN4(n134), .IN5(n257), 
        .Q(n252) );
  OA22X1 U778 ( .IN1(n1297), .IN2(n136), .IN3(n1201), .IN4(n137), .Q(n257) );
  OA221X1 U779 ( .IN1(n1265), .IN2(n138), .IN3(n1894), .IN4(n139), .IN5(n258), 
        .Q(n251) );
  OA22X1 U780 ( .IN1(n1137), .IN2(n141), .IN3(n1009), .IN4(n86), .Q(n258) );
  MUX21X1 U781 ( .IN1(n259), .IN2(\fifo[0][17] ), .S(clear), .Q(N141) );
  NAND4X0 U782 ( .IN1(n260), .IN2(n261), .IN3(n262), .IN4(n263), .QN(n259) );
  OA221X1 U783 ( .IN1(n1170), .IN2(n123), .IN3(n1949), .IN4(n124), .IN5(n264), 
        .Q(n263) );
  OA22X1 U784 ( .IN1(n1042), .IN2(n126), .IN3(n1927), .IN4(n127), .Q(n264) );
  OA221X1 U785 ( .IN1(n978), .IN2(n128), .IN3(n1106), .IN4(n129), .IN5(n265), 
        .Q(n262) );
  OA22X1 U786 ( .IN1(n1863), .IN2(n131), .IN3(n1234), .IN4(n132), .Q(n265) );
  OA221X1 U787 ( .IN1(n946), .IN2(n133), .IN3(n1074), .IN4(n134), .IN5(n266), 
        .Q(n261) );
  OA22X1 U788 ( .IN1(n1298), .IN2(n136), .IN3(n1202), .IN4(n137), .Q(n266) );
  OA221X1 U789 ( .IN1(n1266), .IN2(n138), .IN3(n1895), .IN4(n139), .IN5(n267), 
        .Q(n260) );
  OA22X1 U790 ( .IN1(n1138), .IN2(n141), .IN3(n1010), .IN4(n86), .Q(n267) );
  MUX21X1 U791 ( .IN1(n268), .IN2(\fifo[0][16] ), .S(clear), .Q(N140) );
  NAND4X0 U792 ( .IN1(n269), .IN2(n270), .IN3(n271), .IN4(n272), .QN(n268) );
  OA221X1 U793 ( .IN1(n1171), .IN2(n123), .IN3(n1950), .IN4(n124), .IN5(n273), 
        .Q(n272) );
  OA22X1 U794 ( .IN1(n1043), .IN2(n126), .IN3(n1928), .IN4(n127), .Q(n273) );
  OA221X1 U795 ( .IN1(n979), .IN2(n128), .IN3(n1107), .IN4(n129), .IN5(n274), 
        .Q(n271) );
  OA22X1 U796 ( .IN1(n1864), .IN2(n131), .IN3(n1235), .IN4(n132), .Q(n274) );
  OA221X1 U797 ( .IN1(n947), .IN2(n133), .IN3(n1075), .IN4(n134), .IN5(n275), 
        .Q(n270) );
  OA22X1 U798 ( .IN1(n1299), .IN2(n136), .IN3(n1203), .IN4(n137), .Q(n275) );
  OA221X1 U799 ( .IN1(n1267), .IN2(n138), .IN3(n1896), .IN4(n139), .IN5(n276), 
        .Q(n269) );
  OA22X1 U800 ( .IN1(n1139), .IN2(n141), .IN3(n1011), .IN4(n86), .Q(n276) );
  MUX21X1 U801 ( .IN1(n277), .IN2(\fifo[0][15] ), .S(clear), .Q(N139) );
  NAND4X0 U802 ( .IN1(n278), .IN2(n279), .IN3(n280), .IN4(n281), .QN(n277) );
  OA221X1 U803 ( .IN1(n1172), .IN2(n123), .IN3(n1951), .IN4(n124), .IN5(n282), 
        .Q(n281) );
  OA22X1 U804 ( .IN1(n1044), .IN2(n126), .IN3(n1929), .IN4(n127), .Q(n282) );
  OA221X1 U805 ( .IN1(n980), .IN2(n128), .IN3(n1108), .IN4(n129), .IN5(n283), 
        .Q(n280) );
  OA22X1 U806 ( .IN1(n1865), .IN2(n131), .IN3(n1236), .IN4(n132), .Q(n283) );
  OA221X1 U807 ( .IN1(n948), .IN2(n133), .IN3(n1076), .IN4(n134), .IN5(n284), 
        .Q(n279) );
  OA22X1 U808 ( .IN1(n1300), .IN2(n136), .IN3(n1204), .IN4(n137), .Q(n284) );
  OA221X1 U809 ( .IN1(n1268), .IN2(n138), .IN3(n1897), .IN4(n139), .IN5(n285), 
        .Q(n278) );
  OA22X1 U810 ( .IN1(n1140), .IN2(n141), .IN3(n1012), .IN4(n86), .Q(n285) );
  MUX21X1 U811 ( .IN1(n286), .IN2(\fifo[0][14] ), .S(clear), .Q(N138) );
  NAND4X0 U812 ( .IN1(n287), .IN2(n288), .IN3(n289), .IN4(n290), .QN(n286) );
  OA221X1 U813 ( .IN1(n1173), .IN2(n123), .IN3(n1952), .IN4(n124), .IN5(n291), 
        .Q(n290) );
  OA22X1 U814 ( .IN1(n1045), .IN2(n126), .IN3(n1930), .IN4(n127), .Q(n291) );
  OA221X1 U815 ( .IN1(n981), .IN2(n128), .IN3(n1109), .IN4(n129), .IN5(n292), 
        .Q(n289) );
  OA22X1 U816 ( .IN1(n1866), .IN2(n131), .IN3(n1237), .IN4(n132), .Q(n292) );
  OA221X1 U817 ( .IN1(n949), .IN2(n133), .IN3(n1077), .IN4(n134), .IN5(n293), 
        .Q(n288) );
  OA22X1 U818 ( .IN1(n1301), .IN2(n136), .IN3(n1205), .IN4(n137), .Q(n293) );
  OA221X1 U819 ( .IN1(n1269), .IN2(n138), .IN3(n1898), .IN4(n139), .IN5(n294), 
        .Q(n287) );
  OA22X1 U820 ( .IN1(n1141), .IN2(n141), .IN3(n1013), .IN4(n86), .Q(n294) );
  MUX21X1 U821 ( .IN1(n295), .IN2(\fifo[0][13] ), .S(clear), .Q(N137) );
  NAND4X0 U822 ( .IN1(n296), .IN2(n297), .IN3(n298), .IN4(n299), .QN(n295) );
  OA221X1 U823 ( .IN1(n1174), .IN2(n123), .IN3(n1953), .IN4(n124), .IN5(n300), 
        .Q(n299) );
  OA22X1 U824 ( .IN1(n1046), .IN2(n126), .IN3(n1931), .IN4(n127), .Q(n300) );
  OA221X1 U825 ( .IN1(n982), .IN2(n128), .IN3(n1110), .IN4(n129), .IN5(n301), 
        .Q(n298) );
  OA22X1 U826 ( .IN1(n1867), .IN2(n131), .IN3(n1238), .IN4(n132), .Q(n301) );
  OA221X1 U827 ( .IN1(n950), .IN2(n133), .IN3(n1078), .IN4(n134), .IN5(n302), 
        .Q(n297) );
  OA22X1 U828 ( .IN1(n1302), .IN2(n136), .IN3(n1206), .IN4(n137), .Q(n302) );
  OA221X1 U829 ( .IN1(n1270), .IN2(n138), .IN3(n1899), .IN4(n139), .IN5(n303), 
        .Q(n296) );
  OA22X1 U830 ( .IN1(n1142), .IN2(n141), .IN3(n1014), .IN4(n86), .Q(n303) );
  MUX21X1 U831 ( .IN1(n304), .IN2(\fifo[0][12] ), .S(clear), .Q(N136) );
  NAND4X0 U832 ( .IN1(n305), .IN2(n306), .IN3(n307), .IN4(n308), .QN(n304) );
  OA221X1 U833 ( .IN1(n1175), .IN2(n123), .IN3(n1954), .IN4(n124), .IN5(n309), 
        .Q(n308) );
  OA22X1 U834 ( .IN1(n1047), .IN2(n126), .IN3(n1932), .IN4(n127), .Q(n309) );
  OA221X1 U835 ( .IN1(n983), .IN2(n128), .IN3(n1111), .IN4(n129), .IN5(n310), 
        .Q(n307) );
  OA22X1 U836 ( .IN1(n1868), .IN2(n131), .IN3(n1239), .IN4(n132), .Q(n310) );
  OA221X1 U837 ( .IN1(n951), .IN2(n133), .IN3(n1079), .IN4(n134), .IN5(n311), 
        .Q(n306) );
  OA22X1 U838 ( .IN1(n1303), .IN2(n136), .IN3(n1207), .IN4(n137), .Q(n311) );
  OA221X1 U839 ( .IN1(n1271), .IN2(n138), .IN3(n1900), .IN4(n139), .IN5(n312), 
        .Q(n305) );
  OA22X1 U840 ( .IN1(n1143), .IN2(n141), .IN3(n1015), .IN4(n86), .Q(n312) );
  MUX21X1 U841 ( .IN1(n313), .IN2(\fifo[0][11] ), .S(clear), .Q(N135) );
  NAND4X0 U842 ( .IN1(n314), .IN2(n315), .IN3(n316), .IN4(n317), .QN(n313) );
  OA221X1 U843 ( .IN1(n1176), .IN2(n123), .IN3(n1955), .IN4(n124), .IN5(n318), 
        .Q(n317) );
  OA22X1 U844 ( .IN1(n1048), .IN2(n126), .IN3(n1933), .IN4(n127), .Q(n318) );
  OA221X1 U845 ( .IN1(n984), .IN2(n128), .IN3(n1112), .IN4(n129), .IN5(n319), 
        .Q(n316) );
  OA22X1 U846 ( .IN1(n1869), .IN2(n131), .IN3(n1240), .IN4(n132), .Q(n319) );
  OA221X1 U847 ( .IN1(n952), .IN2(n133), .IN3(n1080), .IN4(n134), .IN5(n320), 
        .Q(n315) );
  OA22X1 U848 ( .IN1(n1304), .IN2(n136), .IN3(n1208), .IN4(n137), .Q(n320) );
  OA221X1 U849 ( .IN1(n1272), .IN2(n138), .IN3(n1901), .IN4(n139), .IN5(n321), 
        .Q(n314) );
  OA22X1 U850 ( .IN1(n1144), .IN2(n141), .IN3(n1016), .IN4(n86), .Q(n321) );
  MUX21X1 U851 ( .IN1(n322), .IN2(\fifo[0][10] ), .S(clear), .Q(N134) );
  NAND4X0 U852 ( .IN1(n323), .IN2(n324), .IN3(n325), .IN4(n326), .QN(n322) );
  OA221X1 U853 ( .IN1(n1177), .IN2(n123), .IN3(n1956), .IN4(n124), .IN5(n327), 
        .Q(n326) );
  OA22X1 U854 ( .IN1(n1049), .IN2(n126), .IN3(n1934), .IN4(n127), .Q(n327) );
  OA221X1 U855 ( .IN1(n985), .IN2(n128), .IN3(n1113), .IN4(n129), .IN5(n328), 
        .Q(n325) );
  OA22X1 U856 ( .IN1(n1870), .IN2(n131), .IN3(n1241), .IN4(n132), .Q(n328) );
  OA221X1 U857 ( .IN1(n953), .IN2(n133), .IN3(n1081), .IN4(n134), .IN5(n329), 
        .Q(n324) );
  OA22X1 U858 ( .IN1(n1305), .IN2(n136), .IN3(n1209), .IN4(n137), .Q(n329) );
  OA221X1 U859 ( .IN1(n1273), .IN2(n138), .IN3(n1902), .IN4(n139), .IN5(n330), 
        .Q(n323) );
  OA22X1 U860 ( .IN1(n1145), .IN2(n141), .IN3(n1017), .IN4(n86), .Q(n330) );
  MUX21X1 U861 ( .IN1(n331), .IN2(\fifo[0][9] ), .S(clear), .Q(N133) );
  NAND4X0 U862 ( .IN1(n332), .IN2(n333), .IN3(n334), .IN4(n335), .QN(n331) );
  OA221X1 U863 ( .IN1(n1178), .IN2(n123), .IN3(n1957), .IN4(n124), .IN5(n336), 
        .Q(n335) );
  OA22X1 U864 ( .IN1(n1050), .IN2(n126), .IN3(n922), .IN4(n127), .Q(n336) );
  OA221X1 U865 ( .IN1(n986), .IN2(n128), .IN3(n1114), .IN4(n129), .IN5(n337), 
        .Q(n334) );
  OA22X1 U866 ( .IN1(n1871), .IN2(n131), .IN3(n1242), .IN4(n132), .Q(n337) );
  OA221X1 U867 ( .IN1(n954), .IN2(n133), .IN3(n1082), .IN4(n134), .IN5(n338), 
        .Q(n333) );
  OA22X1 U868 ( .IN1(n1306), .IN2(n136), .IN3(n1210), .IN4(n137), .Q(n338) );
  OA221X1 U869 ( .IN1(n1274), .IN2(n138), .IN3(n1903), .IN4(n139), .IN5(n339), 
        .Q(n332) );
  OA22X1 U870 ( .IN1(n1146), .IN2(n141), .IN3(n1018), .IN4(n86), .Q(n339) );
  MUX21X1 U871 ( .IN1(n340), .IN2(\fifo[0][8] ), .S(clear), .Q(N132) );
  NAND4X0 U872 ( .IN1(n341), .IN2(n342), .IN3(n343), .IN4(n344), .QN(n340) );
  OA221X1 U873 ( .IN1(n1179), .IN2(n123), .IN3(n1958), .IN4(n124), .IN5(n345), 
        .Q(n344) );
  OA22X1 U874 ( .IN1(n1051), .IN2(n126), .IN3(n923), .IN4(n127), .Q(n345) );
  OA221X1 U875 ( .IN1(n987), .IN2(n128), .IN3(n1115), .IN4(n129), .IN5(n346), 
        .Q(n343) );
  OA22X1 U876 ( .IN1(n1872), .IN2(n131), .IN3(n1243), .IN4(n132), .Q(n346) );
  OA221X1 U877 ( .IN1(n955), .IN2(n133), .IN3(n1083), .IN4(n134), .IN5(n347), 
        .Q(n342) );
  OA22X1 U878 ( .IN1(n1307), .IN2(n136), .IN3(n1211), .IN4(n137), .Q(n347) );
  OA221X1 U879 ( .IN1(n1275), .IN2(n138), .IN3(n1904), .IN4(n139), .IN5(n348), 
        .Q(n341) );
  OA22X1 U880 ( .IN1(n1147), .IN2(n141), .IN3(n1019), .IN4(n86), .Q(n348) );
  MUX21X1 U881 ( .IN1(n349), .IN2(\fifo[0][7] ), .S(clear), .Q(N131) );
  NAND4X0 U882 ( .IN1(n350), .IN2(n351), .IN3(n352), .IN4(n353), .QN(n349) );
  OA221X1 U883 ( .IN1(n1180), .IN2(n123), .IN3(n1959), .IN4(n124), .IN5(n354), 
        .Q(n353) );
  OA22X1 U884 ( .IN1(n1052), .IN2(n126), .IN3(n924), .IN4(n127), .Q(n354) );
  OA221X1 U885 ( .IN1(n988), .IN2(n128), .IN3(n1116), .IN4(n129), .IN5(n355), 
        .Q(n352) );
  OA22X1 U886 ( .IN1(n1873), .IN2(n131), .IN3(n1244), .IN4(n132), .Q(n355) );
  OA221X1 U887 ( .IN1(n956), .IN2(n133), .IN3(n1084), .IN4(n134), .IN5(n356), 
        .Q(n351) );
  OA22X1 U888 ( .IN1(n1308), .IN2(n136), .IN3(n1212), .IN4(n137), .Q(n356) );
  OA221X1 U889 ( .IN1(n1276), .IN2(n138), .IN3(n1905), .IN4(n139), .IN5(n357), 
        .Q(n350) );
  OA22X1 U890 ( .IN1(n1148), .IN2(n141), .IN3(n1020), .IN4(n86), .Q(n357) );
  MUX21X1 U891 ( .IN1(n358), .IN2(\fifo[0][6] ), .S(clear), .Q(N130) );
  NAND4X0 U892 ( .IN1(n359), .IN2(n360), .IN3(n361), .IN4(n362), .QN(n358) );
  OA221X1 U893 ( .IN1(n1181), .IN2(n123), .IN3(n1960), .IN4(n124), .IN5(n363), 
        .Q(n362) );
  OA22X1 U894 ( .IN1(n1053), .IN2(n126), .IN3(n925), .IN4(n127), .Q(n363) );
  OA221X1 U895 ( .IN1(n989), .IN2(n128), .IN3(n1117), .IN4(n129), .IN5(n364), 
        .Q(n361) );
  OA22X1 U896 ( .IN1(n1874), .IN2(n131), .IN3(n1245), .IN4(n132), .Q(n364) );
  OA221X1 U897 ( .IN1(n957), .IN2(n133), .IN3(n1085), .IN4(n134), .IN5(n365), 
        .Q(n360) );
  OA22X1 U898 ( .IN1(n1309), .IN2(n136), .IN3(n1213), .IN4(n137), .Q(n365) );
  OA221X1 U899 ( .IN1(n1277), .IN2(n138), .IN3(n1906), .IN4(n139), .IN5(n366), 
        .Q(n359) );
  OA22X1 U900 ( .IN1(n1149), .IN2(n141), .IN3(n1021), .IN4(n86), .Q(n366) );
  MUX21X1 U901 ( .IN1(n367), .IN2(\fifo[0][5] ), .S(clear), .Q(N129) );
  NAND4X0 U902 ( .IN1(n368), .IN2(n369), .IN3(n370), .IN4(n371), .QN(n367) );
  OA221X1 U903 ( .IN1(n1182), .IN2(n123), .IN3(n1961), .IN4(n124), .IN5(n372), 
        .Q(n371) );
  OA22X1 U904 ( .IN1(n1054), .IN2(n126), .IN3(n926), .IN4(n127), .Q(n372) );
  OA221X1 U905 ( .IN1(n990), .IN2(n128), .IN3(n1118), .IN4(n129), .IN5(n373), 
        .Q(n370) );
  OA22X1 U906 ( .IN1(n1875), .IN2(n131), .IN3(n1246), .IN4(n132), .Q(n373) );
  OA221X1 U907 ( .IN1(n958), .IN2(n133), .IN3(n1086), .IN4(n134), .IN5(n374), 
        .Q(n369) );
  OA22X1 U908 ( .IN1(n1310), .IN2(n136), .IN3(n1214), .IN4(n137), .Q(n374) );
  OA221X1 U909 ( .IN1(n1278), .IN2(n138), .IN3(n1907), .IN4(n139), .IN5(n375), 
        .Q(n368) );
  OA22X1 U910 ( .IN1(n1150), .IN2(n141), .IN3(n1022), .IN4(n86), .Q(n375) );
  MUX21X1 U911 ( .IN1(n376), .IN2(\fifo[0][4] ), .S(clear), .Q(N128) );
  NAND4X0 U912 ( .IN1(n377), .IN2(n378), .IN3(n379), .IN4(n380), .QN(n376) );
  OA221X1 U913 ( .IN1(n1183), .IN2(n123), .IN3(n1962), .IN4(n124), .IN5(n381), 
        .Q(n380) );
  OA22X1 U914 ( .IN1(n1055), .IN2(n126), .IN3(n927), .IN4(n127), .Q(n381) );
  OA221X1 U915 ( .IN1(n991), .IN2(n128), .IN3(n1119), .IN4(n129), .IN5(n382), 
        .Q(n379) );
  OA22X1 U916 ( .IN1(n1876), .IN2(n131), .IN3(n1247), .IN4(n132), .Q(n382) );
  OA221X1 U917 ( .IN1(n959), .IN2(n133), .IN3(n1087), .IN4(n134), .IN5(n383), 
        .Q(n378) );
  OA22X1 U918 ( .IN1(n1314), .IN2(n136), .IN3(n1215), .IN4(n137), .Q(n383) );
  OA221X1 U919 ( .IN1(n1279), .IN2(n138), .IN3(n1908), .IN4(n139), .IN5(n384), 
        .Q(n377) );
  OA22X1 U920 ( .IN1(n1151), .IN2(n141), .IN3(n1023), .IN4(n86), .Q(n384) );
  MUX21X1 U921 ( .IN1(n385), .IN2(\fifo[0][3] ), .S(clear), .Q(N127) );
  NAND4X0 U922 ( .IN1(n386), .IN2(n387), .IN3(n388), .IN4(n389), .QN(n385) );
  OA221X1 U923 ( .IN1(n1184), .IN2(n123), .IN3(n1963), .IN4(n124), .IN5(n390), 
        .Q(n389) );
  OA22X1 U924 ( .IN1(n1056), .IN2(n126), .IN3(n928), .IN4(n127), .Q(n390) );
  OA221X1 U925 ( .IN1(n992), .IN2(n128), .IN3(n1120), .IN4(n129), .IN5(n391), 
        .Q(n388) );
  OA22X1 U926 ( .IN1(n1877), .IN2(n131), .IN3(n1248), .IN4(n132), .Q(n391) );
  OA221X1 U927 ( .IN1(n960), .IN2(n133), .IN3(n1088), .IN4(n134), .IN5(n392), 
        .Q(n387) );
  OA22X1 U928 ( .IN1(n1315), .IN2(n136), .IN3(n1216), .IN4(n137), .Q(n392) );
  OA221X1 U929 ( .IN1(n1280), .IN2(n138), .IN3(n1909), .IN4(n139), .IN5(n393), 
        .Q(n386) );
  OA22X1 U930 ( .IN1(n1152), .IN2(n141), .IN3(n1024), .IN4(n86), .Q(n393) );
  MUX21X1 U931 ( .IN1(n394), .IN2(\fifo[0][2] ), .S(clear), .Q(N126) );
  NAND4X0 U932 ( .IN1(n395), .IN2(n396), .IN3(n397), .IN4(n398), .QN(n394) );
  OA221X1 U933 ( .IN1(n1185), .IN2(n123), .IN3(n1964), .IN4(n124), .IN5(n399), 
        .Q(n398) );
  OA22X1 U934 ( .IN1(n1057), .IN2(n126), .IN3(n929), .IN4(n127), .Q(n399) );
  OA221X1 U935 ( .IN1(n993), .IN2(n128), .IN3(n1121), .IN4(n129), .IN5(n400), 
        .Q(n397) );
  OA22X1 U936 ( .IN1(n1878), .IN2(n131), .IN3(n1249), .IN4(n132), .Q(n400) );
  OA221X1 U937 ( .IN1(n961), .IN2(n133), .IN3(n1089), .IN4(n134), .IN5(n401), 
        .Q(n396) );
  OA22X1 U938 ( .IN1(n1316), .IN2(n136), .IN3(n1217), .IN4(n137), .Q(n401) );
  OA221X1 U939 ( .IN1(n1281), .IN2(n138), .IN3(n1910), .IN4(n139), .IN5(n402), 
        .Q(n395) );
  OA22X1 U940 ( .IN1(n1153), .IN2(n141), .IN3(n1025), .IN4(n86), .Q(n402) );
  MUX21X1 U941 ( .IN1(n403), .IN2(\fifo[0][1] ), .S(clear), .Q(N125) );
  NAND4X0 U942 ( .IN1(n404), .IN2(n405), .IN3(n406), .IN4(n407), .QN(n403) );
  OA221X1 U943 ( .IN1(n1186), .IN2(n123), .IN3(n1965), .IN4(n124), .IN5(n408), 
        .Q(n407) );
  OA22X1 U944 ( .IN1(n1058), .IN2(n126), .IN3(n930), .IN4(n127), .Q(n408) );
  OA221X1 U945 ( .IN1(n994), .IN2(n128), .IN3(n1122), .IN4(n129), .IN5(n409), 
        .Q(n406) );
  OA22X1 U946 ( .IN1(n1879), .IN2(n131), .IN3(n1250), .IN4(n132), .Q(n409) );
  OA221X1 U947 ( .IN1(n962), .IN2(n133), .IN3(n1090), .IN4(n134), .IN5(n410), 
        .Q(n405) );
  OA22X1 U948 ( .IN1(n1317), .IN2(n136), .IN3(n1218), .IN4(n137), .Q(n410) );
  OA221X1 U949 ( .IN1(n1282), .IN2(n138), .IN3(n1911), .IN4(n139), .IN5(n411), 
        .Q(n404) );
  OA22X1 U950 ( .IN1(n1154), .IN2(n141), .IN3(n1026), .IN4(n86), .Q(n411) );
  MUX21X1 U951 ( .IN1(n412), .IN2(\fifo[0][0] ), .S(clear), .Q(N124) );
  NAND4X0 U952 ( .IN1(n413), .IN2(n414), .IN3(n415), .IN4(n416), .QN(n412) );
  OA221X1 U953 ( .IN1(n1187), .IN2(n123), .IN3(n1966), .IN4(n124), .IN5(n417), 
        .Q(n416) );
  OA22X1 U954 ( .IN1(n1059), .IN2(n126), .IN3(n931), .IN4(n127), .Q(n417) );
  NAND2X0 U955 ( .IN1(n418), .IN2(n419), .QN(n127) );
  NAND2X0 U956 ( .IN1(n420), .IN2(n418), .QN(n126) );
  NAND2X0 U957 ( .IN1(n421), .IN2(n418), .QN(n124) );
  NAND2X0 U958 ( .IN1(n422), .IN2(n418), .QN(n123) );
  AND2X1 U959 ( .IN1(n1844), .IN2(n426), .Q(n418) );
  OA221X1 U960 ( .IN1(n995), .IN2(n128), .IN3(n1123), .IN4(n129), .IN5(n423), 
        .Q(n415) );
  OA22X1 U961 ( .IN1(n1880), .IN2(n131), .IN3(n1251), .IN4(n132), .Q(n423) );
  NAND2X0 U962 ( .IN1(n95), .IN2(n422), .QN(n132) );
  NAND2X0 U963 ( .IN1(n95), .IN2(n421), .QN(n131) );
  NAND2X0 U964 ( .IN1(n95), .IN2(n420), .QN(n129) );
  NAND2X0 U965 ( .IN1(n95), .IN2(n419), .QN(n128) );
  AND2X1 U966 ( .IN1(n426), .IN2(N15), .Q(n95) );
  OA221X1 U967 ( .IN1(n963), .IN2(n133), .IN3(n1091), .IN4(n134), .IN5(n424), 
        .Q(n414) );
  OA22X1 U968 ( .IN1(n1843), .IN2(n136), .IN3(n1219), .IN4(n137), .Q(n424) );
  NAND2X0 U969 ( .IN1(n94), .IN2(n422), .QN(n137) );
  NAND2X0 U970 ( .IN1(n94), .IN2(n421), .QN(n136) );
  NAND2X0 U971 ( .IN1(n94), .IN2(n420), .QN(n134) );
  NAND2X0 U972 ( .IN1(n94), .IN2(n419), .QN(n133) );
  NOR2X0 U973 ( .IN1(N15), .IN2(n426), .QN(n94) );
  OA221X1 U974 ( .IN1(n1283), .IN2(n138), .IN3(n1912), .IN4(n139), .IN5(n425), 
        .Q(n413) );
  OA22X1 U975 ( .IN1(n1155), .IN2(n141), .IN3(n1027), .IN4(n86), .Q(n425) );
  NAND2X0 U976 ( .IN1(n92), .IN2(n419), .QN(n86) );
  NOR2X0 U977 ( .IN1(N17), .IN2(n1845), .QN(n419) );
  NAND2X0 U978 ( .IN1(n420), .IN2(n92), .QN(n141) );
  INVX0 U979 ( .INP(n87), .ZN(n420) );
  NAND2X0 U980 ( .IN1(n1845), .IN2(N17), .QN(n87) );
  NAND2X0 U981 ( .IN1(n421), .IN2(n92), .QN(n139) );
  AND2X1 U982 ( .IN1(n1846), .IN2(n1845), .Q(n421) );
  NAND2X0 U983 ( .IN1(n422), .IN2(n92), .QN(n138) );
  NOR2X0 U984 ( .IN1(n1844), .IN2(n426), .QN(n92) );
  NOR2X0 U985 ( .IN1(n1846), .IN2(n1845), .QN(n422) );
endmodule


module eth_wishbone_DW01_inc_0 ( A, SUM );
  input [29:0] A;
  output [29:0] SUM;

  wire   [29:2] carry;

  HADDX1 U1_1_28 ( .A0(A[28]), .B0(carry[28]), .C1(carry[29]), .SO(SUM[28]) );
  HADDX1 U1_1_27 ( .A0(A[27]), .B0(carry[27]), .C1(carry[28]), .SO(SUM[27]) );
  HADDX1 U1_1_26 ( .A0(A[26]), .B0(carry[26]), .C1(carry[27]), .SO(SUM[26]) );
  HADDX1 U1_1_25 ( .A0(A[25]), .B0(carry[25]), .C1(carry[26]), .SO(SUM[25]) );
  HADDX1 U1_1_24 ( .A0(A[24]), .B0(carry[24]), .C1(carry[25]), .SO(SUM[24]) );
  HADDX1 U1_1_23 ( .A0(A[23]), .B0(carry[23]), .C1(carry[24]), .SO(SUM[23]) );
  HADDX1 U1_1_22 ( .A0(A[22]), .B0(carry[22]), .C1(carry[23]), .SO(SUM[22]) );
  HADDX1 U1_1_21 ( .A0(A[21]), .B0(carry[21]), .C1(carry[22]), .SO(SUM[21]) );
  HADDX1 U1_1_20 ( .A0(A[20]), .B0(carry[20]), .C1(carry[21]), .SO(SUM[20]) );
  HADDX1 U1_1_19 ( .A0(A[19]), .B0(carry[19]), .C1(carry[20]), .SO(SUM[19]) );
  HADDX1 U1_1_18 ( .A0(A[18]), .B0(carry[18]), .C1(carry[19]), .SO(SUM[18]) );
  HADDX1 U1_1_17 ( .A0(A[17]), .B0(carry[17]), .C1(carry[18]), .SO(SUM[17]) );
  HADDX1 U1_1_16 ( .A0(A[16]), .B0(carry[16]), .C1(carry[17]), .SO(SUM[16]) );
  HADDX1 U1_1_15 ( .A0(A[15]), .B0(carry[15]), .C1(carry[16]), .SO(SUM[15]) );
  HADDX1 U1_1_14 ( .A0(A[14]), .B0(carry[14]), .C1(carry[15]), .SO(SUM[14]) );
  HADDX1 U1_1_13 ( .A0(A[13]), .B0(carry[13]), .C1(carry[14]), .SO(SUM[13]) );
  HADDX1 U1_1_12 ( .A0(A[12]), .B0(carry[12]), .C1(carry[13]), .SO(SUM[12]) );
  HADDX1 U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1 U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1 U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1 U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  XOR2X1 U2 ( .IN1(carry[29]), .IN2(A[29]), .Q(SUM[29]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module eth_wishbone_DW01_inc_1 ( A, SUM );
  input [29:0] A;
  output [29:0] SUM;

  wire   [29:2] carry;

  HADDX1 U1_1_28 ( .A0(A[28]), .B0(carry[28]), .C1(carry[29]), .SO(SUM[28]) );
  HADDX1 U1_1_27 ( .A0(A[27]), .B0(carry[27]), .C1(carry[28]), .SO(SUM[27]) );
  HADDX1 U1_1_26 ( .A0(A[26]), .B0(carry[26]), .C1(carry[27]), .SO(SUM[26]) );
  HADDX1 U1_1_25 ( .A0(A[25]), .B0(carry[25]), .C1(carry[26]), .SO(SUM[25]) );
  HADDX1 U1_1_24 ( .A0(A[24]), .B0(carry[24]), .C1(carry[25]), .SO(SUM[24]) );
  HADDX1 U1_1_23 ( .A0(A[23]), .B0(carry[23]), .C1(carry[24]), .SO(SUM[23]) );
  HADDX1 U1_1_22 ( .A0(A[22]), .B0(carry[22]), .C1(carry[23]), .SO(SUM[22]) );
  HADDX1 U1_1_21 ( .A0(A[21]), .B0(carry[21]), .C1(carry[22]), .SO(SUM[21]) );
  HADDX1 U1_1_20 ( .A0(A[20]), .B0(carry[20]), .C1(carry[21]), .SO(SUM[20]) );
  HADDX1 U1_1_19 ( .A0(A[19]), .B0(carry[19]), .C1(carry[20]), .SO(SUM[19]) );
  HADDX1 U1_1_18 ( .A0(A[18]), .B0(carry[18]), .C1(carry[19]), .SO(SUM[18]) );
  HADDX1 U1_1_17 ( .A0(A[17]), .B0(carry[17]), .C1(carry[18]), .SO(SUM[17]) );
  HADDX1 U1_1_16 ( .A0(A[16]), .B0(carry[16]), .C1(carry[17]), .SO(SUM[16]) );
  HADDX1 U1_1_15 ( .A0(A[15]), .B0(carry[15]), .C1(carry[16]), .SO(SUM[15]) );
  HADDX1 U1_1_14 ( .A0(A[14]), .B0(carry[14]), .C1(carry[15]), .SO(SUM[14]) );
  HADDX1 U1_1_13 ( .A0(A[13]), .B0(carry[13]), .C1(carry[14]), .SO(SUM[13]) );
  HADDX1 U1_1_12 ( .A0(A[12]), .B0(carry[12]), .C1(carry[13]), .SO(SUM[12]) );
  HADDX1 U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1 U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1 U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1 U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  XOR2X1 U2 ( .IN1(carry[29]), .IN2(A[29]), .Q(SUM[29]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module eth_wishbone_DW01_inc_2 ( A, SUM );
  input [29:0] A;
  output [29:0] SUM;

  wire   [29:2] carry;

  HADDX1 U1_1_28 ( .A0(A[28]), .B0(carry[28]), .C1(carry[29]), .SO(SUM[28]) );
  HADDX1 U1_1_27 ( .A0(A[27]), .B0(carry[27]), .C1(carry[28]), .SO(SUM[27]) );
  HADDX1 U1_1_26 ( .A0(A[26]), .B0(carry[26]), .C1(carry[27]), .SO(SUM[26]) );
  HADDX1 U1_1_25 ( .A0(A[25]), .B0(carry[25]), .C1(carry[26]), .SO(SUM[25]) );
  HADDX1 U1_1_24 ( .A0(A[24]), .B0(carry[24]), .C1(carry[25]), .SO(SUM[24]) );
  HADDX1 U1_1_23 ( .A0(A[23]), .B0(carry[23]), .C1(carry[24]), .SO(SUM[23]) );
  HADDX1 U1_1_22 ( .A0(A[22]), .B0(carry[22]), .C1(carry[23]), .SO(SUM[22]) );
  HADDX1 U1_1_21 ( .A0(A[21]), .B0(carry[21]), .C1(carry[22]), .SO(SUM[21]) );
  HADDX1 U1_1_20 ( .A0(A[20]), .B0(carry[20]), .C1(carry[21]), .SO(SUM[20]) );
  HADDX1 U1_1_19 ( .A0(A[19]), .B0(carry[19]), .C1(carry[20]), .SO(SUM[19]) );
  HADDX1 U1_1_18 ( .A0(A[18]), .B0(carry[18]), .C1(carry[19]), .SO(SUM[18]) );
  HADDX1 U1_1_17 ( .A0(A[17]), .B0(carry[17]), .C1(carry[18]), .SO(SUM[17]) );
  HADDX1 U1_1_16 ( .A0(A[16]), .B0(carry[16]), .C1(carry[17]), .SO(SUM[16]) );
  HADDX1 U1_1_15 ( .A0(A[15]), .B0(carry[15]), .C1(carry[16]), .SO(SUM[15]) );
  HADDX1 U1_1_14 ( .A0(A[14]), .B0(carry[14]), .C1(carry[15]), .SO(SUM[14]) );
  HADDX1 U1_1_13 ( .A0(A[13]), .B0(carry[13]), .C1(carry[14]), .SO(SUM[13]) );
  HADDX1 U1_1_12 ( .A0(A[12]), .B0(carry[12]), .C1(carry[13]), .SO(SUM[12]) );
  HADDX1 U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1 U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1 U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1 U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  XOR2X1 U2 ( .IN1(carry[29]), .IN2(A[29]), .Q(SUM[29]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module eth_wishbone_DW01_inc_3 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  XOR2X1 U2 ( .IN1(carry[6]), .IN2(A[6]), .Q(SUM[6]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module eth_wishbone_DW01_inc_4 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  XOR2X1 U2 ( .IN1(carry[6]), .IN2(A[6]), .Q(SUM[6]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module eth_wishbone_test_1 ( WB_CLK_I, WB_DAT_I, WB_DAT_O, WB_ADR_I, WB_WE_I, 
        WB_ACK_O, BDCs, Reset, m_wb_adr_o, m_wb_sel_o, m_wb_we_o, m_wb_dat_o, 
        m_wb_dat_i, m_wb_cyc_o, m_wb_stb_o, m_wb_ack_i, m_wb_err_i, MTxClk, 
        TxStartFrm, TxEndFrm, TxUsedData, TxData, TxRetry, TxAbort, TxUnderRun, 
        TxDone, PerPacketCrcEn, PerPacketPad, MRxClk, RxData, RxValid, 
        RxStartFrm, RxEndFrm, RxAbort, RxStatusWriteLatched_sync2, r_TxEn, 
        r_RxEn, r_TxBDNum, r_RxFlow, r_PassAll, TxB_IRQ, TxE_IRQ, RxB_IRQ, 
        RxE_IRQ, Busy_IRQ, InvalidSymbol, LatchedCrcError, RxLateCollision, 
        ShortFrame, DribbleNibble, ReceivedPacketTooBig, RxLength, 
        LoadRxStatus, ReceivedPacketGood, AddressMiss, ReceivedPauseFrm, 
        RetryCntLatched, RetryLimit, LateCollLatched, DeferLatched, 
        RstDeferLatched, CarrierSenseLost, eth_top_test_point_11887_in, 
        test_si8, test_si7, test_si6, test_si5, test_si4, test_si3, test_si2, 
        test_si1, test_so7, test_so6, test_so5, test_so4, test_so3, test_so2, 
        test_so1, test_se );
  input [31:0] WB_DAT_I;
  output [31:0] WB_DAT_O;
  input [9:2] WB_ADR_I;
  input [3:0] BDCs;
  output [29:0] m_wb_adr_o;
  output [3:0] m_wb_sel_o;
  output [31:0] m_wb_dat_o;
  input [31:0] m_wb_dat_i;
  output [7:0] TxData;
  input [7:0] RxData;
  input [7:0] r_TxBDNum;
  input [15:0] RxLength;
  input [3:0] RetryCntLatched;
  input WB_CLK_I, WB_WE_I, Reset, m_wb_ack_i, m_wb_err_i, MTxClk, TxUsedData,
         TxRetry, TxAbort, TxDone, MRxClk, RxValid, RxStartFrm, RxEndFrm,
         RxAbort, r_TxEn, r_RxEn, r_RxFlow, r_PassAll, InvalidSymbol,
         LatchedCrcError, RxLateCollision, ShortFrame, DribbleNibble,
         ReceivedPacketTooBig, LoadRxStatus, ReceivedPacketGood, AddressMiss,
         ReceivedPauseFrm, RetryLimit, LateCollLatched, DeferLatched,
         CarrierSenseLost, eth_top_test_point_11887_in, test_si8, test_si7,
         test_si6, test_si5, test_si4, test_si3, test_si2, test_si1, test_se;
  output WB_ACK_O, m_wb_we_o, m_wb_cyc_o, m_wb_stb_o, TxStartFrm, TxEndFrm,
         TxUnderRun, PerPacketCrcEn, PerPacketPad, RxStatusWriteLatched_sync2,
         TxB_IRQ, TxE_IRQ, RxB_IRQ, RxE_IRQ, Busy_IRQ, RstDeferLatched,
         test_so7, test_so6, test_so5, test_so4, test_so3, test_so2, test_so1;
  wire   m_wb_cyc_o, WbEn, N76, ram_oe, TxEn, RxEn, BlockingTxStatusWrite,
         TxDone_wb, TxAbort_wb, BlockingTxStatusWrite_sync1,
         BlockingTxStatusWrite_sync2, BlockingTxStatusWrite_sync3, N350, N351,
         N352, N353, N354, N355, N356, N357, N358, N359, N360, N361, N362,
         N363, N364, N365, N366, N367, N368, N369, N370, N371, N372, N373,
         N374, N375, N376, N377, N378, N379, tx_burst_en, TxBufferAlmostFull,
         rx_burst_en, N651, N652, N653, N654, N655, N656, N657, N658, N659,
         N660, N661, N662, N663, N664, N665, N666, N667, N668, N669, N670,
         N671, N672, N673, N674, N675, N676, N677, N678, N679, N680, _1_net_,
         TxBufferFull, TxBufferAlmostEmpty, TxBufferEmpty, TxStartFrm_wb,
         TxStartFrm_sync1, TxStartFrm_sync2, TxStartFrm_syncb1,
         LatchValidBytes, N792, N800, N801, N802, N803, N804, N805, N806, N807,
         N808, N809, N810, N811, N812, N813, TxRetry_wb, N837, N848, N857,
         ReadTxDataFromFifo_tck, ReadTxDataFromFifo_syncb2,
         ReadTxDataFromFifo_sync1, ReadTxDataFromFifo_sync2,
         ReadTxDataFromFifo_syncb1, TxRetrySync1, TxDoneSync1, TxAbortSync1,
         RxAbortSync3, RxAbortSync2, N998, N999, N1000, N1001, N1002, N1003,
         N1004, N1005, N1006, N1007, N1008, N1009, N1010, N1011, N1012, N1013,
         N1014, N1015, N1016, N1017, N1018, N1019, N1020, N1021, N1022, N1023,
         N1024, N1025, N1026, N1027, ShiftEnded_rck, WriteRxDataToFifo,
         WriteRxDataToFifoSync2, WriteRxDataToFifoSync1, SyncRxStartFrm_q,
         LatchedRxStartFrm, SyncRxStartFrm, SyncRxStartFrm_q2, RxFifoReset,
         _2_net_, RxBufferFull, RxBufferAlmostEmpty, RxBufferEmpty,
         ShiftEndedSync_c1, ShiftEndedSync1, ShiftEndedSync2, RxAbortSync1,
         RxAbortLatched, RxAbortSyncb1, RxStatusWriteLatched,
         RxStatusWriteLatched_sync1, RxStatusWriteLatched_syncb1, N1258, N1261,
         N1265, N1268, Busy_IRQ_rck, Busy_IRQ_sync1, Busy_IRQ_sync3,
         Busy_IRQ_sync2, Busy_IRQ_syncb1, n676, n679, n705, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n723, n724, n838, n840, n842, n847, n848, n849, n860, n883,
         n1088, n1091, n1094, n1097, n1100, n1103, n1106, n1109, n1112, n1115,
         n1118, n1121, n1124, n1127, n1130, n1133, n1157, n1159, n1264, n1266,
         n1288, n1297, n1299, n1301, n1335, n1338, n1340, n1342, n1344, n1346,
         n1348, n1350, n1352, n1354, n1356, n1358, n1360, n1362, n1364, n1366,
         n1368, n1370, n1372, n1374, n1376, n1378, n1380, n1382, n1384, n1419,
         n1420, n1429, n1433, n1435, n1445, n1448, n1449, n1450, n1451, n1452,
         n1463, n1464, n1465, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n3, n4, n8, n9, n11, n12, n19, n28, n29, n30, n32, n33,
         n35, n36, n37, n38, n43, n50, n54, n59, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n675, n677, n678, n680, n681, n682,
         n683, n684, n685, n686, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n706,
         n722, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n738, n739, n740, n741, n742, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n985, n987, n989, n990, n991, n993, n994, n995, n996, n1188, n1, n2,
         n5, n6, n7, n10, n13, n14, n15, n16, n17, n18, n20, n21, n22, n23,
         n24, n25, n26, n27, n31, n34, n39, n40, n41, n42, n44, n45, n46, n47,
         n48, n49, n51, n52, n53, n55, n56, n57, n58, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n652, n674, n687, n737,
         n743, n744, n745, n746, n747, n748, n749, n765, n766, n767;
  wire   [3:0] ram_we;
  wire   [7:0] ram_addr;
  wire   [31:0] ram_di;
  wire   [7:1] TxBDAddress;
  wire   [7:1] RxBDAddress;
  wire   [31:2] TxPointerMSB;
  wire   [2:0] tx_burst_cnt;
  wire   [2:0] rx_burst_cnt;
  wire   [31:2] RxPointerMSB;
  wire   [4:0] txfifo_cnt;
  wire   [31:0] TxData_wb;
  wire   [31:0] RxDataLatched2;
  wire   [4:0] rxfifo_cnt;
  tri   [31:0] WB_DAT_O;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;
  assign m_wb_stb_o = m_wb_cyc_o;

  SDFFARX1 r_TxEn_q_reg ( .D(r_TxEn), .SI(n741), .SE(test_se), .CLK(n75), 
        .RSTB(n26), .Q(n740), .QN(n766) );
  SDFFARX1 r_RxEn_q_reg ( .D(r_RxEn), .SI(m_wb_we_o), .SE(test_se), .CLK(n72), 
        .RSTB(n46), .Q(n741), .QN(n765) );
  SDFFARX1 TxRetry_q_reg ( .D(TxRetry), .SI(TxRetrySync1), .SE(test_se), .CLK(
        n78), .RSTB(n26), .Q(n691), .QN(n536) );
  SDFFARX1 Flop_reg ( .D(n1806), .SI(n764), .SE(test_se), .CLK(n78), .RSTB(n26), .Q(n686), .QN(n749) );
  SDFFARX1 TxUsedData_q_reg ( .D(TxUsedData), .SI(n654), .SE(test_se), .CLK(
        n80), .RSTB(n39), .Q(n750), .QN(n724) );
  SDFFARX1 TxAbort_q_reg ( .D(TxAbort), .SI(TxAbortSync1), .SE(test_se), .CLK(
        n78), .RSTB(n22), .Q(n690), .QN(n537) );
  SDFFARX1 TxRetrySync1_reg ( .D(TxRetry), .SI(n729), .SE(test_se), .CLK(n71), 
        .RSTB(n23), .Q(TxRetrySync1) );
  SDFFARX1 TxRetry_wb_reg ( .D(TxRetrySync1), .SI(n554), .SE(test_se), .CLK(
        n71), .RSTB(n23), .Q(TxRetry_wb), .QN(n1450) );
  SDFFARX1 TxRetry_wb_q_reg ( .D(TxRetry_wb), .SI(n691), .SE(test_se), .CLK(
        n75), .RSTB(n26), .Q(n554), .QN(n996) );
  SDFFARX1 TxDoneSync1_reg ( .D(TxDone), .SI(n753), .SE(test_se), .CLK(n72), 
        .RSTB(n41), .Q(TxDoneSync1) );
  SDFFARX1 TxDone_wb_reg ( .D(TxDoneSync1), .SI(n698), .SE(test_se), .CLK(n72), 
        .RSTB(n41), .Q(TxDone_wb), .QN(n1451) );
  SDFFARX1 TxDone_wb_q_reg ( .D(TxDone_wb), .SI(TxDoneSync1), .SE(test_se), 
        .CLK(n72), .RSTB(n42), .Q(n698), .QN(n995) );
  SDFFARX1 TxAbortSync1_reg ( .D(TxAbort), .SI(n730), .SE(test_se), .CLK(n74), 
        .RSTB(n60), .Q(TxAbortSync1) );
  SDFFARX1 TxAbort_wb_reg ( .D(TxAbortSync1), .SI(n696), .SE(test_se), .CLK(
        n71), .RSTB(n22), .Q(TxAbort_wb), .QN(n1452) );
  SDFFARX1 TxAbort_wb_q_reg ( .D(TxAbort_wb), .SI(n690), .SE(test_se), .CLK(
        n71), .RSTB(n22), .Q(n696) );
  SDFFARX1 SyncRxStartFrm_q_reg ( .D(SyncRxStartFrm), .SI(SyncRxStartFrm_q2), 
        .SE(test_se), .CLK(n74), .RSTB(n31), .Q(SyncRxStartFrm_q), .QN(n1464)
         );
  SDFFARX1 LatchedRxStartFrm_reg ( .D(n1805), .SI(n684), .SE(test_se), .CLK(
        n83), .RSTB(n31), .Q(LatchedRxStartFrm) );
  SDFFARX1 SyncRxStartFrm_reg ( .D(LatchedRxStartFrm), .SI(SyncRxStartFrm_q), 
        .SE(test_se), .CLK(n74), .RSTB(n31), .Q(SyncRxStartFrm) );
  SDFFARX1 SyncRxStartFrm_q2_reg ( .D(SyncRxStartFrm_q), .SI(n590), .SE(
        test_se), .CLK(n74), .RSTB(n31), .Q(SyncRxStartFrm_q2) );
  SDFFARX1 RxEnableWindow_reg ( .D(n1804), .SI(RxEn), .SE(test_se), .CLK(n83), 
        .RSTB(n60), .Q(n685) );
  SDFFARX1 RxAbortLatched_reg ( .D(n1803), .SI(n760), .SE(test_se), .CLK(n81), 
        .RSTB(n22), .Q(RxAbortLatched) );
  SDFFARX1 RxAbortSync1_reg ( .D(RxAbortLatched), .SI(RxAbortLatched), .SE(
        test_se), .CLK(n71), .RSTB(n23), .Q(RxAbortSync1) );
  SDFFARX1 RxAbortSync2_reg ( .D(RxAbortSync1), .SI(RxAbortSync1), .SE(test_se), .CLK(n71), .RSTB(n23), .Q(RxAbortSync2), .QN(n676) );
  SDFFARX1 RxAbortSync3_reg ( .D(RxAbortSync2), .SI(RxAbortSync2), .SE(test_se), .CLK(n71), .RSTB(n23), .Q(RxAbortSync3) );
  SDFFARX1 RxAbortSync4_reg ( .D(RxAbortSync3), .SI(RxAbortSync3), .SE(test_se), .CLK(n71), .RSTB(n23), .Q(n759), .QN(n532) );
  SDFFARX1 RxAbortSyncb1_reg ( .D(RxAbortSync2), .SI(n759), .SE(test_se), 
        .CLK(n81), .RSTB(n23), .Q(RxAbortSyncb1) );
  SDFFARX1 RxAbortSyncb2_reg ( .D(RxAbortSyncb1), .SI(RxAbortSyncb1), .SE(
        test_se), .CLK(n81), .RSTB(n23), .Q(n758), .QN(n842) );
  SDFFARX1 \LatchedRxLength_reg[15]  ( .D(n1384), .SI(n683), .SE(test_se), 
        .CLK(n83), .RSTB(n31), .Q(n684) );
  SDFFARX1 \LatchedRxLength_reg[14]  ( .D(n1382), .SI(n682), .SE(test_se), 
        .CLK(n83), .RSTB(n31), .Q(n683) );
  SDFFARX1 \LatchedRxLength_reg[13]  ( .D(n1380), .SI(n681), .SE(test_se), 
        .CLK(n82), .RSTB(n31), .Q(n682) );
  SDFFARX1 \LatchedRxLength_reg[12]  ( .D(n1378), .SI(n680), .SE(test_se), 
        .CLK(n82), .RSTB(n27), .Q(n681) );
  SDFFARX1 \LatchedRxLength_reg[11]  ( .D(n1376), .SI(n678), .SE(test_se), 
        .CLK(n82), .RSTB(n27), .Q(n680) );
  SDFFARX1 \LatchedRxLength_reg[10]  ( .D(n1374), .SI(n677), .SE(test_se), 
        .CLK(n82), .RSTB(n27), .Q(n678) );
  SDFFARX1 \LatchedRxLength_reg[9]  ( .D(n1372), .SI(n675), .SE(test_se), 
        .CLK(n82), .RSTB(n27), .Q(n677) );
  SDFFARX1 \LatchedRxLength_reg[8]  ( .D(n1370), .SI(n673), .SE(test_se), 
        .CLK(n82), .RSTB(n27), .Q(n675) );
  SDFFARX1 \LatchedRxLength_reg[7]  ( .D(n1368), .SI(n672), .SE(test_se), 
        .CLK(n82), .RSTB(n27), .Q(n673) );
  SDFFARX1 \LatchedRxLength_reg[6]  ( .D(n1366), .SI(n671), .SE(test_se), 
        .CLK(n82), .RSTB(n27), .Q(n672) );
  SDFFARX1 \LatchedRxLength_reg[5]  ( .D(n1364), .SI(n670), .SE(test_se), 
        .CLK(n82), .RSTB(n27), .Q(n671) );
  SDFFARX1 \LatchedRxLength_reg[4]  ( .D(n1362), .SI(n669), .SE(test_se), 
        .CLK(n82), .RSTB(n27), .Q(n670) );
  SDFFARX1 \LatchedRxLength_reg[3]  ( .D(n1360), .SI(n668), .SE(test_se), 
        .CLK(n82), .RSTB(n27), .Q(n669) );
  SDFFARX1 \LatchedRxLength_reg[2]  ( .D(n1358), .SI(n667), .SE(test_se), 
        .CLK(n82), .RSTB(n27), .Q(n668) );
  SDFFARX1 \LatchedRxLength_reg[1]  ( .D(n1356), .SI(n666), .SE(test_se), 
        .CLK(n81), .RSTB(n27), .Q(n667) );
  SDFFARX1 \LatchedRxLength_reg[0]  ( .D(n1354), .SI(LatchValidBytes), .SE(
        test_se), .CLK(n81), .RSTB(n26), .Q(n666) );
  SDFFARX1 \RxStatusInLatched_reg[8]  ( .D(n1352), .SI(n664), .SE(test_se), 
        .CLK(n83), .RSTB(n63), .Q(n665) );
  SDFFARX1 \RxStatusInLatched_reg[7]  ( .D(n1350), .SI(n656), .SE(test_se), 
        .CLK(n83), .RSTB(n63), .Q(n664) );
  SDFFARX1 \RxStatusInLatched_reg[5]  ( .D(n1348), .SI(n662), .SE(test_se), 
        .CLK(n83), .RSTB(n31), .Q(n663) );
  SDFFARX1 \RxStatusInLatched_reg[4]  ( .D(n1346), .SI(n661), .SE(test_se), 
        .CLK(n83), .RSTB(n31), .Q(n662) );
  SDFFARX1 \RxStatusInLatched_reg[3]  ( .D(n1344), .SI(n660), .SE(test_se), 
        .CLK(n82), .RSTB(n31), .Q(n661) );
  SDFFARX1 \RxStatusInLatched_reg[2]  ( .D(n1342), .SI(n659), .SE(test_se), 
        .CLK(n81), .RSTB(n22), .Q(n660) );
  SDFFARX1 \RxStatusInLatched_reg[1]  ( .D(n1340), .SI(n658), .SE(test_se), 
        .CLK(n81), .RSTB(n22), .Q(n659) );
  SDFFARX1 \RxStatusInLatched_reg[0]  ( .D(n1338), .SI(n640), .SE(test_se), 
        .CLK(n84), .RSTB(n22), .Q(n658) );
  SDFFARX1 RxOverrun_reg ( .D(n1802), .SI(n685), .SE(test_se), .CLK(n74), 
        .RSTB(n63), .Q(n657) );
  SDFFARX1 \RxStatusInLatched_reg[6]  ( .D(n1335), .SI(n663), .SE(test_se), 
        .CLK(n83), .RSTB(n63), .Q(n656) );
  SDFFARX1 \ram_di_reg[6]  ( .D(n1677), .SI(ram_di[5]), .SE(test_se), .CLK(n72), .RSTB(n48), .Q(ram_di[6]) );
  SDFFARX1 \TxLength_reg[15]  ( .D(n1800), .SI(n32), .SE(test_se), .CLK(n73), 
        .RSTB(n51), .Q(n54) );
  SDFFARX1 LatchValidBytes_reg ( .D(N792), .SI(n763), .SE(test_se), .CLK(n72), 
        .RSTB(n39), .Q(LatchValidBytes) );
  SDFFARX1 LatchValidBytes_q_reg ( .D(LatchValidBytes), .SI(n692), .SE(test_se), .CLK(n72), .RSTB(n39), .Q(n763), .QN(n1435) );
  SDFFARX1 \TxValidBytesLatched_reg[0]  ( .D(n1632), .SI(n750), .SE(test_se), 
        .CLK(n72), .RSTB(n39), .Q(n655), .QN(n990) );
  SDFFARX1 TxEndFrm_reg ( .D(n1630), .SI(TxEn), .SE(test_se), .CLK(n80), 
        .RSTB(n39), .Q(TxEndFrm), .QN(n1445) );
  SDFFARX1 LastWord_reg ( .D(n1629), .SI(n706), .SE(test_se), .CLK(n80), 
        .RSTB(n39), .Q(n692), .QN(n748) );
  SDFFARX1 ReadTxDataFromFifo_tck_reg ( .D(n1628), .SI(n761), .SE(test_se), 
        .CLK(n80), .RSTB(n39), .Q(ReadTxDataFromFifo_tck) );
  SDFFARX1 ReadTxDataFromFifo_sync1_reg ( .D(ReadTxDataFromFifo_tck), .SI(n727), .SE(test_se), .CLK(n72), .RSTB(n39), .Q(ReadTxDataFromFifo_sync1) );
  SDFFARX1 ReadTxDataFromFifo_sync2_reg ( .D(ReadTxDataFromFifo_sync1), .SI(
        ReadTxDataFromFifo_sync1), .SE(test_se), .CLK(n72), .RSTB(n39), .Q(
        ReadTxDataFromFifo_sync2) );
  SDFFARX1 ReadTxDataFromFifo_syncb1_reg ( .D(ReadTxDataFromFifo_sync2), .SI(
        n762), .SE(test_se), .CLK(n76), .RSTB(n60), .Q(
        ReadTxDataFromFifo_syncb1) );
  SDFFARX1 ReadTxDataFromFifo_syncb2_reg ( .D(ReadTxDataFromFifo_syncb1), .SI(
        ReadTxDataFromFifo_syncb1), .SE(test_se), .CLK(n76), .RSTB(n60), .Q(
        ReadTxDataFromFifo_syncb2) );
  SDFFARX1 ReadTxDataFromFifo_syncb3_reg ( .D(ReadTxDataFromFifo_syncb2), .SI(
        ReadTxDataFromFifo_syncb2), .SE(test_se), .CLK(n76), .RSTB(n20), .Q(
        n761), .QN(n1448) );
  SDFFARX1 ReadTxDataFromFifo_sync3_reg ( .D(ReadTxDataFromFifo_sync2), .SI(
        ReadTxDataFromFifo_sync2), .SE(test_se), .CLK(n72), .RSTB(n39), .Q(
        n762), .QN(n1449) );
  SDFFARX1 TxUnderRun_wb_reg ( .D(n1581), .SI(n648), .SE(test_se), .CLK(n72), 
        .RSTB(n39), .Q(n654) );
  SDFFARX1 BlockReadTxDataFromMemory_reg ( .D(n1799), .SI(n641), .SE(test_se), 
        .CLK(n73), .RSTB(n34), .Q(n653) );
  SDFFARX1 \tx_burst_cnt_reg[2]  ( .D(n1798), .SI(tx_burst_cnt[1]), .SE(
        test_se), .CLK(n74), .RSTB(n49), .Q(tx_burst_cnt[2]) );
  SDFFASX1 tx_burst_en_reg ( .D(n1797), .SI(tx_burst_cnt[2]), .SE(test_se), 
        .CLK(n70), .SETB(n69), .Q(tx_burst_en), .QN(n6) );
  SDFFARX1 TxDonePacket_reg ( .D(N857), .SI(n735), .SE(test_se), .CLK(n72), 
        .RSTB(n41), .Q(n753), .QN(n534) );
  SDFFARX1 TxDonePacketBlocked_reg ( .D(n1709), .SI(TxData[7]), .SE(test_se), 
        .CLK(n72), .RSTB(n41), .Q(n651) );
  SDFFARX1 TxRetryPacket_reg ( .D(N848), .SI(n726), .SE(test_se), .CLK(n71), 
        .RSTB(n23), .Q(n729), .QN(n14) );
  SDFFARX1 TxRetryPacketBlocked_reg ( .D(n1708), .SI(n725), .SE(test_se), 
        .CLK(n73), .RSTB(n57), .Q(n650) );
  SDFFARX1 TxAbortPacket_reg ( .D(N837), .SI(n736), .SE(test_se), .CLK(n71), 
        .RSTB(n22), .Q(n730) );
  SDFFARX1 TxAbortPacketBlocked_reg ( .D(n1796), .SI(SyncRxStartFrm), .SE(
        test_se), .CLK(n74), .RSTB(n31), .Q(n649) );
  SDFFARX1 TxAbortPacket_NotCleared_reg ( .D(n1795), .SI(n649), .SE(test_se), 
        .CLK(n74), .RSTB(n61), .Q(n736), .QN(n747) );
  SDFFARX1 BlockingTxStatusWrite_reg ( .D(n1564), .SI(n555), .SE(test_se), 
        .CLK(n72), .RSTB(n42), .Q(BlockingTxStatusWrite), .QN(n1419) );
  SDFFARX1 BlockingTxStatusWrite_sync1_reg ( .D(BlockingTxStatusWrite), .SI(
        BlockingTxStatusWrite), .SE(test_se), .CLK(n78), .RSTB(n42), .Q(
        BlockingTxStatusWrite_sync1) );
  SDFFARX1 BlockingTxStatusWrite_sync2_reg ( .D(BlockingTxStatusWrite_sync1), 
        .SI(BlockingTxStatusWrite_sync1), .SE(test_se), .CLK(n78), .RSTB(n42), 
        .Q(BlockingTxStatusWrite_sync2), .QN(n1420) );
  SDFFARX1 BlockingTxStatusWrite_sync3_reg ( .D(BlockingTxStatusWrite_sync2), 
        .SI(BlockingTxStatusWrite_sync2), .SE(test_se), .CLK(n78), .RSTB(n42), 
        .Q(BlockingTxStatusWrite_sync3) );
  SDFFARX1 TxUnderRun_sync1_reg ( .D(n1563), .SI(TxUnderRun), .SE(test_se), 
        .CLK(n78), .RSTB(n31), .Q(n648) );
  SDFFARX1 TxUnderRun_reg ( .D(n1562), .SI(n646), .SE(test_se), .CLK(n78), 
        .RSTB(n25), .Q(TxUnderRun) );
  SDFFASX1 TxBDRead_reg ( .D(n1794), .SI(TxBDAddress[7]), .SE(test_se), .CLK(
        n70), .SETB(n69), .Q(n731) );
  SDFFARX1 \TxStatus_reg[11]  ( .D(n1301), .SI(TxStartFrm_wb), .SE(test_se), 
        .CLK(n72), .RSTB(n25), .Q(PerPacketCrcEn) );
  SDFFARX1 \TxStatus_reg[12]  ( .D(n1299), .SI(PerPacketCrcEn), .SE(test_se), 
        .CLK(n74), .RSTB(n25), .Q(PerPacketPad) );
  SDFFARX1 \TxStatus_reg[13]  ( .D(n1297), .SI(PerPacketPad), .SE(test_se), 
        .CLK(n75), .RSTB(n25), .Q(n647) );
  SDFFARX1 \TxBDAddress_reg[1]  ( .D(n1579), .SI(TxAbort_wb), .SE(test_se), 
        .CLK(n75), .RSTB(n26), .Q(TxBDAddress[1]) );
  SDFFARX1 \TxBDAddress_reg[2]  ( .D(n1578), .SI(TxBDAddress[1]), .SE(test_se), 
        .CLK(n74), .RSTB(n26), .Q(TxBDAddress[2]) );
  SDFFARX1 \TxBDAddress_reg[3]  ( .D(n1577), .SI(TxBDAddress[2]), .SE(test_se), 
        .CLK(n75), .RSTB(n26), .Q(TxBDAddress[3]) );
  SDFFARX1 \TxBDAddress_reg[4]  ( .D(n1576), .SI(TxBDAddress[3]), .SE(test_se), 
        .CLK(n74), .RSTB(n26), .Q(TxBDAddress[4]) );
  SDFFARX1 \TxBDAddress_reg[5]  ( .D(n1575), .SI(TxBDAddress[4]), .SE(test_se), 
        .CLK(n74), .RSTB(n26), .Q(TxBDAddress[5]) );
  SDFFARX1 \TxBDAddress_reg[6]  ( .D(n1574), .SI(TxBDAddress[5]), .SE(test_se), 
        .CLK(n74), .RSTB(n26), .Q(TxBDAddress[6]) );
  SDFFARX1 \TxBDAddress_reg[7]  ( .D(n1573), .SI(TxBDAddress[6]), .SE(test_se), 
        .CLK(n74), .RSTB(n26), .Q(TxBDAddress[7]) );
  SDFFARX1 \TxStatus_reg[14]  ( .D(n1288), .SI(n647), .SE(test_se), .CLK(n75), 
        .RSTB(n25), .Q(n646), .QN(n10) );
  SDFFARX1 TxBDReady_reg ( .D(n1652), .SI(n731), .SE(test_se), .CLK(n73), 
        .RSTB(n39), .Q(n733), .QN(n746) );
  SDFFARX1 TxEn_needed_reg ( .D(n1792), .SI(TxE_IRQ), .SE(test_se), .CLK(n74), 
        .RSTB(n34), .Q(n645), .QN(n538) );
  SDFFARX1 TxEn_reg ( .D(n1791), .SI(n752), .SE(test_se), .CLK(n74), .RSTB(n65), .Q(TxEn), .QN(n883) );
  SDFFARX1 TxEn_q_reg ( .D(TxEn), .SI(n645), .SE(test_se), .CLK(n74), .RSTB(
        n60), .Q(n752), .QN(n745) );
  SDFFARX1 TxPointerRead_reg ( .D(n1793), .SI(TxPointerMSB[31]), .SE(test_se), 
        .CLK(n71), .RSTB(n24), .Q(n725) );
  SDFFARX1 \BDWrite_reg[0]  ( .D(n1691), .SI(n608), .SE(test_se), .CLK(n74), 
        .RSTB(n61), .Q(n644) );
  SDFFARX1 \BDWrite_reg[1]  ( .D(n1690), .SI(n644), .SE(test_se), .CLK(n74), 
        .RSTB(n61), .Q(n643) );
  SDFFARX1 \BDWrite_reg[2]  ( .D(n1689), .SI(n643), .SE(test_se), .CLK(n74), 
        .RSTB(n61), .Q(n642) );
  SDFFARX1 \BDWrite_reg[3]  ( .D(n1688), .SI(n642), .SE(test_se), .CLK(n74), 
        .RSTB(n61), .Q(n641) );
  SDFFASX1 WbEn_reg ( .D(n1686), .SI(n734), .SE(test_se), .CLK(n70), .SETB(n69), .Q(WbEn), .QN(n838) );
  SDFFARX1 WbEn_q_reg ( .D(WbEn), .SI(WB_ACK_O), .SE(test_se), .CLK(n71), 
        .RSTB(n23), .Q(n734), .QN(n744) );
  SDFFARX1 RxEn_needed_reg ( .D(n1692), .SI(RxE_IRQ), .SE(test_se), .CLK(n73), 
        .RSTB(n42), .Q(n732), .QN(n743) );
  SDFFARX1 \ram_di_reg[15]  ( .D(n1668), .SI(ram_di[14]), .SE(test_se), .CLK(
        n71), .RSTB(n20), .Q(ram_di[15]) );
  SDFFARX1 \ram_di_reg[10]  ( .D(n1673), .SI(ram_di[9]), .SE(test_se), .CLK(
        n72), .RSTB(n48), .Q(ram_di[10]) );
  SDFFARX1 \ram_di_reg[9]  ( .D(n1674), .SI(ram_di[8]), .SE(test_se), .CLK(n72), .RSTB(n48), .Q(ram_di[9]) );
  SDFFARX1 RxEn_reg ( .D(n1790), .SI(n757), .SE(test_se), .CLK(n74), .RSTB(n60), .Q(RxEn) );
  SDFFARX1 RxEn_q_reg ( .D(RxEn), .SI(n732), .SE(test_se), .CLK(n74), .RSTB(
        n61), .Q(n757), .QN(n737) );
  SDFFARX1 ShiftEnded_reg ( .D(n1789), .SI(ShiftEnded_rck), .SE(test_se), 
        .CLK(n74), .RSTB(n64), .Q(n754), .QN(n687) );
  SDFFARX1 RxReady_reg ( .D(n1788), .SI(n722), .SE(test_se), .CLK(n71), .RSTB(
        n21), .Q(n640), .QN(n8) );
  SDFFARX1 RxBDRead_reg ( .D(n1787), .SI(RxBDAddress[7]), .SE(test_se), .CLK(
        n71), .RSTB(n24), .Q(n697) );
  SDFFARX1 \RxStatus_reg[14]  ( .D(n1266), .SI(n638), .SE(test_se), .CLK(n71), 
        .RSTB(n25), .Q(n639), .QN(n674) );
  SDFFARX1 \RxStatus_reg[13]  ( .D(n1264), .SI(n756), .SE(test_se), .CLK(n74), 
        .RSTB(n65), .Q(n638) );
  SDFFARX1 RxBDReady_reg ( .D(n1685), .SI(n697), .SE(test_se), .CLK(n71), 
        .RSTB(n24), .Q(n637), .QN(n535) );
  SDFFARX1 RxPointerRead_reg ( .D(n1779), .SI(RxPointerMSB[31]), .SE(test_se), 
        .CLK(n71), .RSTB(n21), .Q(n722) );
  SDFFARX1 \RxByteCnt_reg[1]  ( .D(n1766), .SI(n702), .SE(test_se), .CLK(n84), 
        .RSTB(n65), .Q(n701), .QN(n985) );
  SDFFARX1 ShiftEnded_rck_reg ( .D(n1764), .SI(n755), .SE(test_se), .CLK(n81), 
        .RSTB(n25), .Q(ShiftEnded_rck), .QN(n847) );
  SDFFARX1 ShiftEndedSync1_reg ( .D(ShiftEnded_rck), .SI(n699), .SE(test_se), 
        .CLK(n74), .RSTB(n64), .Q(ShiftEndedSync1) );
  SDFFARX1 ShiftEndedSync2_reg ( .D(ShiftEndedSync1), .SI(ShiftEndedSync1), 
        .SE(test_se), .CLK(n74), .RSTB(n64), .Q(ShiftEndedSync2), .QN(n1465)
         );
  SDFFARX1 ShiftEndedSync_c1_reg ( .D(ShiftEndedSync2), .SI(n609), .SE(test_se), .CLK(n83), .RSTB(n64), .Q(ShiftEndedSync_c1), .QN(n848) );
  SDFFARX1 ShiftEndedSync_c2_reg ( .D(ShiftEndedSync_c1), .SI(
        ShiftEndedSync_c1), .SE(test_se), .CLK(n84), .RSTB(n64), .Q(n755), 
        .QN(n849) );
  SDFFARX1 ShiftWillEnd_reg ( .D(n1762), .SI(n754), .SE(test_se), .CLK(n81), 
        .RSTB(n25), .Q(n636), .QN(n652) );
  SDFFARX1 LastByteIn_reg ( .D(n1761), .SI(n634), .SE(test_se), .CLK(n83), 
        .RSTB(n63), .Q(n706), .QN(n552) );
  SDFFARX1 WriteRxDataToFifo_reg ( .D(n1765), .SI(n556), .SE(test_se), .CLK(
        n83), .RSTB(n62), .Q(WriteRxDataToFifo), .QN(n679) );
  SDFFARX1 WriteRxDataToFifoSync1_reg ( .D(WriteRxDataToFifo), .SI(WbEn), .SE(
        test_se), .CLK(n74), .RSTB(n63), .Q(WriteRxDataToFifoSync1) );
  SDFFARX1 WriteRxDataToFifoSync2_reg ( .D(WriteRxDataToFifoSync1), .SI(
        WriteRxDataToFifoSync1), .SE(test_se), .CLK(n74), .RSTB(n63), .Q(
        WriteRxDataToFifoSync2), .QN(n1463) );
  SDFFARX1 WriteRxDataToFifoSync3_reg ( .D(WriteRxDataToFifoSync2), .SI(
        WriteRxDataToFifoSync2), .SE(test_se), .CLK(n74), .RSTB(n63), .Q(n556), 
        .QN(n59) );
  SDFFARX1 cyc_cleared_reg ( .D(n1706), .SI(n742), .SE(test_se), .CLK(n73), 
        .RSTB(n34), .Q(n728), .QN(n540) );
  SDFFARX1 \tx_burst_cnt_reg[0]  ( .D(n1705), .SI(n739), .SE(test_se), .CLK(
        n74), .RSTB(n49), .Q(tx_burst_cnt[0]) );
  SDFFARX1 \rx_burst_cnt_reg[0]  ( .D(n1703), .SI(ram_di[31]), .SE(test_se), 
        .CLK(n73), .RSTB(n34), .Q(rx_burst_cnt[0]), .QN(n7) );
  SDFFARX1 \rx_burst_cnt_reg[1]  ( .D(n1702), .SI(rx_burst_cnt[0]), .SE(
        test_se), .CLK(n73), .RSTB(n34), .Q(rx_burst_cnt[1]), .QN(n2) );
  SDFFARX1 \tx_burst_cnt_reg[1]  ( .D(n1704), .SI(tx_burst_cnt[0]), .SE(
        test_se), .CLK(n74), .RSTB(n49), .Q(tx_burst_cnt[1]), .QN(n5) );
  SDFFARX1 \rx_burst_cnt_reg[2]  ( .D(n1701), .SI(rx_burst_cnt[1]), .SE(
        test_se), .CLK(n73), .RSTB(n34), .Q(rx_burst_cnt[2]), .QN(n1) );
  SDFFARX1 MasterWbRX_reg ( .D(n1768), .SI(n607), .SE(test_se), .CLK(n72), 
        .RSTB(n42), .Q(n635), .QN(n551) );
  SDFFARX1 rx_burst_en_reg ( .D(n1711), .SI(rx_burst_cnt[2]), .SE(test_se), 
        .CLK(n73), .RSTB(n34), .Q(rx_burst_en) );
  SDFFARX1 MasterWbTX_reg ( .D(n1710), .SI(n635), .SE(test_se), .CLK(n74), 
        .RSTB(n63), .Q(n727), .QN(n550) );
  SDFFARX1 \m_wb_sel_o_reg[0]  ( .D(n1698), .SI(m_wb_cyc_o), .SE(test_se), 
        .CLK(n72), .RSTB(n46), .Q(m_wb_sel_o[0]), .QN(n705) );
  SDFFARX1 m_wb_cyc_o_reg ( .D(n1699), .SI(m_wb_adr_o[29]), .SE(test_se), 
        .CLK(n72), .RSTB(n46), .Q(m_wb_cyc_o) );
  SDFFARX1 m_wb_we_o_reg ( .D(n1700), .SI(m_wb_sel_o[3]), .SE(test_se), .CLK(
        n72), .RSTB(n46), .Q(m_wb_we_o) );
  SDFFARX1 IncrTxPointer_reg ( .D(n1694), .SI(n686), .SE(test_se), .CLK(n74), 
        .RSTB(n63), .Q(n634), .QN(n539) );
  SDFFARX1 BlockingIncrementTxPointer_reg ( .D(n1693), .SI(n653), .SE(test_se), 
        .CLK(n73), .RSTB(n34), .Q(n553) );
  SDFFARX1 \RxPointerLSB_rst_reg[0]  ( .D(n1767), .SI(n657), .SE(test_se), 
        .CLK(n74), .RSTB(n64), .Q(n703), .QN(n549) );
  SDFFARX1 \RxByteCnt_reg[0]  ( .D(n1763), .SI(RxB_IRQ), .SE(test_se), .CLK(
        n81), .RSTB(n25), .Q(n702), .QN(n548) );
  SDFFASX1 \RxValidBytes_reg[0]  ( .D(n1737), .SI(n639), .SE(test_se), .CLK(
        n81), .SETB(n69), .Q(n700), .QN(n9) );
  SDFFARX1 \RxPointerLSB_rst_reg[1]  ( .D(n1778), .SI(n703), .SE(test_se), 
        .CLK(n74), .RSTB(n64), .Q(n704), .QN(n987) );
  SDFFARX1 \RxValidBytes_reg[1]  ( .D(n1736), .SI(n700), .SE(test_se), .CLK(
        n83), .RSTB(n64), .Q(n699), .QN(n547) );
  SDFFARX1 \RxDataLatched2_reg[7]  ( .D(n1728), .SI(RxDataLatched2[6]), .SE(
        test_se), .CLK(n86), .RSTB(n68), .Q(RxDataLatched2[7]) );
  SDFFARX1 \RxDataLatched2_reg[6]  ( .D(n1729), .SI(RxDataLatched2[5]), .SE(
        test_se), .CLK(n86), .RSTB(n68), .Q(RxDataLatched2[6]) );
  SDFFARX1 \RxDataLatched2_reg[5]  ( .D(n1730), .SI(RxDataLatched2[4]), .SE(
        test_se), .CLK(n86), .RSTB(n68), .Q(RxDataLatched2[5]) );
  SDFFARX1 \RxDataLatched2_reg[4]  ( .D(n1731), .SI(RxDataLatched2[3]), .SE(
        test_se), .CLK(n86), .RSTB(n68), .Q(RxDataLatched2[4]) );
  SDFFARX1 \RxDataLatched2_reg[3]  ( .D(n1732), .SI(RxDataLatched2[2]), .SE(
        test_se), .CLK(n86), .RSTB(n67), .Q(RxDataLatched2[3]) );
  SDFFARX1 \RxDataLatched2_reg[2]  ( .D(n1733), .SI(RxDataLatched2[1]), .SE(
        test_se), .CLK(n86), .RSTB(n68), .Q(RxDataLatched2[2]) );
  SDFFARX1 \RxDataLatched2_reg[1]  ( .D(n1734), .SI(RxDataLatched2[0]), .SE(
        test_se), .CLK(n86), .RSTB(n67), .Q(RxDataLatched2[1]) );
  SDFFARX1 \RxDataLatched2_reg[0]  ( .D(n1735), .SI(n624), .SE(test_se), .CLK(
        n86), .RSTB(n68), .Q(RxDataLatched2[0]) );
  SDFFARX1 \RxDataLatched1_reg[16]  ( .D(n1745), .SI(n610), .SE(test_se), 
        .CLK(n85), .RSTB(n66), .Q(n633) );
  SDFFARX1 \RxDataLatched2_reg[16]  ( .D(n1719), .SI(RxDataLatched2[15]), .SE(
        test_se), .CLK(n87), .RSTB(n69), .Q(RxDataLatched2[16]) );
  SDFFARX1 \RxDataLatched1_reg[23]  ( .D(n1744), .SI(n631), .SE(test_se), 
        .CLK(n85), .RSTB(n67), .Q(n632) );
  SDFFARX1 \RxDataLatched2_reg[23]  ( .D(n1712), .SI(RxDataLatched2[22]), .SE(
        test_se), .CLK(n88), .RSTB(n48), .Q(RxDataLatched2[23]) );
  SDFFARX1 \RxDataLatched1_reg[22]  ( .D(n1743), .SI(n630), .SE(test_se), 
        .CLK(n85), .RSTB(n66), .Q(n631) );
  SDFFARX1 \RxDataLatched2_reg[22]  ( .D(n1713), .SI(RxDataLatched2[21]), .SE(
        test_se), .CLK(n87), .RSTB(n55), .Q(RxDataLatched2[22]) );
  SDFFARX1 \RxDataLatched1_reg[21]  ( .D(n1742), .SI(n629), .SE(test_se), 
        .CLK(n85), .RSTB(n67), .Q(n630) );
  SDFFARX1 \RxDataLatched2_reg[21]  ( .D(n1714), .SI(RxDataLatched2[20]), .SE(
        test_se), .CLK(n87), .RSTB(n68), .Q(RxDataLatched2[21]) );
  SDFFARX1 \RxDataLatched1_reg[20]  ( .D(n1741), .SI(n628), .SE(test_se), 
        .CLK(n85), .RSTB(n66), .Q(n629) );
  SDFFARX1 \RxDataLatched2_reg[20]  ( .D(n1715), .SI(RxDataLatched2[19]), .SE(
        test_se), .CLK(n87), .RSTB(n69), .Q(RxDataLatched2[20]) );
  SDFFARX1 \RxDataLatched1_reg[19]  ( .D(n1740), .SI(n627), .SE(test_se), 
        .CLK(n85), .RSTB(n67), .Q(n628) );
  SDFFARX1 \RxDataLatched2_reg[19]  ( .D(n1716), .SI(RxDataLatched2[18]), .SE(
        test_se), .CLK(n87), .RSTB(n69), .Q(RxDataLatched2[19]) );
  SDFFARX1 \RxDataLatched1_reg[18]  ( .D(n1739), .SI(n626), .SE(test_se), 
        .CLK(n85), .RSTB(n66), .Q(n627) );
  SDFFARX1 \RxDataLatched2_reg[18]  ( .D(n1717), .SI(RxDataLatched2[17]), .SE(
        test_se), .CLK(n87), .RSTB(n69), .Q(RxDataLatched2[18]) );
  SDFFARX1 \RxDataLatched1_reg[17]  ( .D(n1738), .SI(n633), .SE(test_se), 
        .CLK(n85), .RSTB(n66), .Q(n626) );
  SDFFARX1 \RxDataLatched2_reg[17]  ( .D(n1718), .SI(RxDataLatched2[16]), .SE(
        test_se), .CLK(n87), .RSTB(n69), .Q(RxDataLatched2[17]) );
  SDFFARX1 \RxDataLatched1_reg[24]  ( .D(n1777), .SI(n632), .SE(test_se), 
        .CLK(n85), .RSTB(n67), .Q(n625) );
  SDFFARX1 \RxDataLatched2_reg[24]  ( .D(n1760), .SI(RxDataLatched2[23]), .SE(
        test_se), .CLK(n88), .RSTB(n48), .Q(RxDataLatched2[24]) );
  SDFFARX1 \RxDataLatched1_reg[31]  ( .D(n1776), .SI(n623), .SE(test_se), 
        .CLK(n86), .RSTB(n68), .Q(n624) );
  SDFFARX1 \RxDataLatched2_reg[31]  ( .D(n1754), .SI(RxDataLatched2[30]), .SE(
        test_se), .CLK(n81), .RSTB(n49), .Q(RxDataLatched2[31]) );
  SDFFARX1 \RxDataLatched1_reg[30]  ( .D(n1775), .SI(n622), .SE(test_se), 
        .CLK(n86), .RSTB(n67), .Q(n623) );
  SDFFARX1 \RxDataLatched2_reg[30]  ( .D(n1755), .SI(RxDataLatched2[29]), .SE(
        test_se), .CLK(n88), .RSTB(n49), .Q(RxDataLatched2[30]) );
  SDFFARX1 \RxDataLatched1_reg[29]  ( .D(n1774), .SI(n621), .SE(test_se), 
        .CLK(n86), .RSTB(n67), .Q(n622) );
  SDFFARX1 \RxDataLatched2_reg[29]  ( .D(n1756), .SI(RxDataLatched2[28]), .SE(
        test_se), .CLK(n88), .RSTB(n49), .Q(RxDataLatched2[29]) );
  SDFFARX1 \RxDataLatched1_reg[28]  ( .D(n1773), .SI(n620), .SE(test_se), 
        .CLK(n85), .RSTB(n67), .Q(n621) );
  SDFFARX1 \RxDataLatched2_reg[28]  ( .D(n1757), .SI(RxDataLatched2[27]), .SE(
        test_se), .CLK(n88), .RSTB(n48), .Q(RxDataLatched2[28]) );
  SDFFARX1 \RxDataLatched1_reg[27]  ( .D(n1772), .SI(n619), .SE(test_se), 
        .CLK(n85), .RSTB(n67), .Q(n620) );
  SDFFARX1 \RxDataLatched2_reg[27]  ( .D(n1758), .SI(RxDataLatched2[26]), .SE(
        test_se), .CLK(n88), .RSTB(n48), .Q(RxDataLatched2[27]) );
  SDFFARX1 \RxDataLatched1_reg[26]  ( .D(n1771), .SI(n618), .SE(test_se), 
        .CLK(n85), .RSTB(n67), .Q(n619) );
  SDFFARX1 \RxDataLatched2_reg[26]  ( .D(n1759), .SI(RxDataLatched2[25]), .SE(
        test_se), .CLK(n88), .RSTB(n48), .Q(RxDataLatched2[26]) );
  SDFFARX1 \RxDataLatched1_reg[25]  ( .D(n1770), .SI(n625), .SE(test_se), 
        .CLK(n85), .RSTB(n67), .Q(n618) );
  SDFFARX1 \RxDataLatched2_reg[25]  ( .D(n1769), .SI(RxDataLatched2[24]), .SE(
        test_se), .CLK(n88), .RSTB(n48), .Q(RxDataLatched2[25]) );
  SDFFARX1 \RxDataLatched1_reg[8]  ( .D(n1753), .SI(n701), .SE(test_se), .CLK(
        n84), .RSTB(n65), .Q(n617) );
  SDFFARX1 \RxDataLatched2_reg[8]  ( .D(n1727), .SI(RxDataLatched2[7]), .SE(
        test_se), .CLK(n86), .RSTB(n68), .Q(RxDataLatched2[8]) );
  SDFFARX1 \RxDataLatched1_reg[9]  ( .D(n1752), .SI(n617), .SE(test_se), .CLK(
        n84), .RSTB(n66), .Q(n616) );
  SDFFARX1 \RxDataLatched2_reg[9]  ( .D(n1726), .SI(RxDataLatched2[8]), .SE(
        test_se), .CLK(n86), .RSTB(n68), .Q(RxDataLatched2[9]) );
  SDFFARX1 \RxDataLatched1_reg[10]  ( .D(n1751), .SI(n616), .SE(test_se), 
        .CLK(n84), .RSTB(n66), .Q(n615) );
  SDFFARX1 \RxDataLatched2_reg[10]  ( .D(n1725), .SI(RxDataLatched2[9]), .SE(
        test_se), .CLK(n87), .RSTB(n68), .Q(RxDataLatched2[10]) );
  SDFFARX1 \RxDataLatched1_reg[11]  ( .D(n1750), .SI(n615), .SE(test_se), 
        .CLK(n84), .RSTB(n66), .Q(n614) );
  SDFFARX1 \RxDataLatched2_reg[11]  ( .D(n1724), .SI(RxDataLatched2[10]), .SE(
        test_se), .CLK(n87), .RSTB(n68), .Q(RxDataLatched2[11]) );
  SDFFARX1 \RxDataLatched1_reg[12]  ( .D(n1749), .SI(n614), .SE(test_se), 
        .CLK(n84), .RSTB(n66), .Q(n613) );
  SDFFARX1 \RxDataLatched2_reg[12]  ( .D(n1723), .SI(RxDataLatched2[11]), .SE(
        test_se), .CLK(n87), .RSTB(n69), .Q(RxDataLatched2[12]) );
  SDFFARX1 \RxDataLatched1_reg[13]  ( .D(n1748), .SI(n613), .SE(test_se), 
        .CLK(n84), .RSTB(n66), .Q(n612) );
  SDFFARX1 \RxDataLatched2_reg[13]  ( .D(n1722), .SI(RxDataLatched2[12]), .SE(
        test_se), .CLK(n87), .RSTB(n69), .Q(RxDataLatched2[13]) );
  SDFFARX1 \RxDataLatched1_reg[14]  ( .D(n1747), .SI(n612), .SE(test_se), 
        .CLK(n84), .RSTB(n66), .Q(n611) );
  SDFFARX1 \RxDataLatched2_reg[14]  ( .D(n1721), .SI(RxDataLatched2[13]), .SE(
        test_se), .CLK(n87), .RSTB(n69), .Q(RxDataLatched2[14]) );
  SDFFARX1 \RxDataLatched1_reg[15]  ( .D(n1746), .SI(n611), .SE(test_se), 
        .CLK(n84), .RSTB(n66), .Q(n610) );
  SDFFARX1 \RxDataLatched2_reg[15]  ( .D(n1720), .SI(RxDataLatched2[14]), .SE(
        test_se), .CLK(n87), .RSTB(n69), .Q(RxDataLatched2[15]) );
  SDFFARX1 \m_wb_sel_o_reg[2]  ( .D(n1696), .SI(m_wb_sel_o[1]), .SE(test_se), 
        .CLK(n72), .RSTB(n46), .Q(m_wb_sel_o[2]) );
  SDFFARX1 \m_wb_sel_o_reg[1]  ( .D(n1697), .SI(m_wb_sel_o[0]), .SE(test_se), 
        .CLK(n72), .RSTB(n46), .Q(m_wb_sel_o[1]) );
  SDFFARX1 \m_wb_sel_o_reg[3]  ( .D(n1695), .SI(m_wb_sel_o[2]), .SE(test_se), 
        .CLK(n72), .RSTB(n46), .Q(m_wb_sel_o[3]) );
  SDFFARX1 ShiftEndedSync3_reg ( .D(n1684), .SI(ShiftEndedSync2), .SE(test_se), 
        .CLK(n74), .RSTB(n64), .Q(n609) );
  SDFFARX1 \RxBDAddress_reg[1]  ( .D(n1786), .SI(n758), .SE(test_se), .CLK(n72), .RSTB(n46), .Q(RxBDAddress[1]) );
  SDFFARX1 \RxBDAddress_reg[2]  ( .D(n1785), .SI(RxBDAddress[1]), .SE(test_se), 
        .CLK(n74), .RSTB(n65), .Q(RxBDAddress[2]) );
  SDFFARX1 \RxBDAddress_reg[3]  ( .D(n1784), .SI(RxBDAddress[2]), .SE(test_se), 
        .CLK(n74), .RSTB(n65), .Q(RxBDAddress[3]) );
  SDFFARX1 \RxBDAddress_reg[4]  ( .D(n1783), .SI(RxBDAddress[3]), .SE(test_se), 
        .CLK(n74), .RSTB(n65), .Q(RxBDAddress[4]) );
  SDFFARX1 \RxBDAddress_reg[5]  ( .D(n1782), .SI(RxBDAddress[4]), .SE(test_se), 
        .CLK(n74), .RSTB(n65), .Q(RxBDAddress[5]) );
  SDFFARX1 \RxBDAddress_reg[6]  ( .D(n1781), .SI(RxBDAddress[5]), .SE(test_se), 
        .CLK(n74), .RSTB(n65), .Q(RxBDAddress[6]) );
  SDFFARX1 \RxBDAddress_reg[7]  ( .D(n1780), .SI(RxBDAddress[6]), .SE(test_se), 
        .CLK(n74), .RSTB(n65), .Q(RxBDAddress[7]) );
  SDFFARX1 BDRead_reg ( .D(n1687), .SI(test_si1), .SE(test_se), .CLK(n74), 
        .RSTB(n61), .Q(n608) );
  SDFFX1 WB_ACK_O_reg ( .D(N76), .SI(n591), .SE(test_se), .CLK(n75), .Q(
        WB_ACK_O) );
  SDFFARX1 TxDonePacket_NotCleared_reg ( .D(n1651), .SI(n651), .SE(test_se), 
        .CLK(n74), .RSTB(n61), .Q(n735), .QN(n13) );
  SDFFARX1 \TxPointerLSB_reg[1]  ( .D(n1159), .SI(n689), .SE(test_se), .CLK(
        n73), .RSTB(n52), .Q(n688), .QN(n546) );
  SDFFARX1 \TxPointerLSB_reg[0]  ( .D(n1157), .SI(n54), .SE(test_se), .CLK(n73), .RSTB(n51), .Q(n689), .QN(n545) );
  SDFFARX1 \TxPointerLSB_rst_reg[1]  ( .D(n1649), .SI(n28), .SE(test_se), 
        .CLK(n73), .RSTB(n52), .Q(n695), .QN(n989) );
  SDFFARX1 \TxPointerLSB_rst_reg[0]  ( .D(n1650), .SI(n688), .SE(test_se), 
        .CLK(n73), .RSTB(n52), .Q(n28), .QN(n840) );
  SDFFARX1 \ram_di_reg[0]  ( .D(n1683), .SI(ram_addr[7]), .SE(test_se), .CLK(
        n72), .RSTB(n47), .Q(ram_di[0]) );
  SDFFARX1 \ram_di_reg[1]  ( .D(n1682), .SI(ram_di[0]), .SE(test_se), .CLK(n72), .RSTB(n47), .Q(ram_di[1]) );
  SDFFARX1 \ram_di_reg[2]  ( .D(n1681), .SI(ram_di[1]), .SE(test_se), .CLK(n72), .RSTB(n47), .Q(ram_di[2]) );
  SDFFARX1 \ram_di_reg[3]  ( .D(n1680), .SI(ram_di[2]), .SE(test_se), .CLK(n72), .RSTB(n47), .Q(ram_di[3]) );
  SDFFARX1 \ram_di_reg[4]  ( .D(n1679), .SI(ram_di[3]), .SE(test_se), .CLK(n72), .RSTB(n47), .Q(ram_di[4]) );
  SDFFARX1 \ram_di_reg[5]  ( .D(n1678), .SI(ram_di[4]), .SE(test_se), .CLK(n72), .RSTB(n47), .Q(ram_di[5]) );
  SDFFARX1 \ram_di_reg[7]  ( .D(n1676), .SI(ram_di[6]), .SE(test_se), .CLK(n72), .RSTB(n48), .Q(ram_di[7]) );
  SDFFARX1 \ram_di_reg[8]  ( .D(n1675), .SI(ram_di[7]), .SE(test_se), .CLK(n72), .RSTB(n48), .Q(ram_di[8]) );
  SDFFARX1 \ram_di_reg[11]  ( .D(n1672), .SI(ram_di[10]), .SE(test_se), .CLK(
        n72), .RSTB(n24), .Q(ram_di[11]) );
  SDFFARX1 \ram_di_reg[12]  ( .D(n1671), .SI(ram_di[11]), .SE(test_se), .CLK(
        n71), .RSTB(n20), .Q(ram_di[12]) );
  SDFFARX1 \ram_di_reg[13]  ( .D(n1670), .SI(ram_di[12]), .SE(test_se), .CLK(
        n71), .RSTB(n20), .Q(ram_di[13]) );
  SDFFARX1 \ram_di_reg[14]  ( .D(n1669), .SI(ram_di[13]), .SE(test_se), .CLK(
        n71), .RSTB(n20), .Q(ram_di[14]) );
  SDFFARX1 \ram_addr_reg[0]  ( .D(n1572), .SI(n740), .SE(test_se), .CLK(n74), 
        .RSTB(n61), .Q(ram_addr[0]) );
  SDFFARX1 \ram_addr_reg[1]  ( .D(n1571), .SI(ram_addr[0]), .SE(test_se), 
        .CLK(n72), .RSTB(n46), .Q(ram_addr[1]) );
  SDFFARX1 \ram_addr_reg[2]  ( .D(n1570), .SI(ram_addr[1]), .SE(test_se), 
        .CLK(n72), .RSTB(n47), .Q(ram_addr[2]) );
  SDFFARX1 \ram_addr_reg[3]  ( .D(n1569), .SI(ram_addr[2]), .SE(test_se), 
        .CLK(n72), .RSTB(n47), .Q(ram_addr[3]) );
  SDFFARX1 \ram_addr_reg[4]  ( .D(n1568), .SI(ram_addr[3]), .SE(test_se), 
        .CLK(n72), .RSTB(n47), .Q(ram_addr[4]) );
  SDFFARX1 \ram_addr_reg[5]  ( .D(n1567), .SI(ram_addr[4]), .SE(test_se), 
        .CLK(n72), .RSTB(n47), .Q(ram_addr[5]) );
  SDFFARX1 \ram_addr_reg[6]  ( .D(n1566), .SI(ram_addr[5]), .SE(test_se), 
        .CLK(n72), .RSTB(n47), .Q(ram_addr[6]) );
  SDFFARX1 \ram_addr_reg[7]  ( .D(n1565), .SI(ram_addr[6]), .SE(test_se), 
        .CLK(n72), .RSTB(n47), .Q(ram_addr[7]) );
  SDFFARX1 \LatchedTxLength_reg[15]  ( .D(n1133), .SI(n606), .SE(test_se), 
        .CLK(n72), .RSTB(n42), .Q(n607) );
  SDFFARX1 \ram_di_reg[31]  ( .D(n1801), .SI(ram_di[30]), .SE(test_se), .CLK(
        n73), .RSTB(n34), .Q(ram_di[31]) );
  SDFFARX1 \LatchedTxLength_reg[14]  ( .D(n1130), .SI(n605), .SE(test_se), 
        .CLK(n71), .RSTB(n60), .Q(n606) );
  SDFFARX1 \ram_di_reg[30]  ( .D(n1653), .SI(ram_di[29]), .SE(test_se), .CLK(
        n71), .RSTB(n21), .Q(ram_di[30]) );
  SDFFARX1 \LatchedTxLength_reg[13]  ( .D(n1127), .SI(n604), .SE(test_se), 
        .CLK(n73), .RSTB(n57), .Q(n605) );
  SDFFARX1 \ram_di_reg[29]  ( .D(n1654), .SI(ram_di[28]), .SE(test_se), .CLK(
        n71), .RSTB(n21), .Q(ram_di[29]) );
  SDFFARX1 \LatchedTxLength_reg[12]  ( .D(n1124), .SI(n603), .SE(test_se), 
        .CLK(n73), .RSTB(n57), .Q(n604) );
  SDFFARX1 \ram_di_reg[28]  ( .D(n1655), .SI(ram_di[27]), .SE(test_se), .CLK(
        n71), .RSTB(n21), .Q(ram_di[28]) );
  SDFFARX1 \LatchedTxLength_reg[11]  ( .D(n1121), .SI(n602), .SE(test_se), 
        .CLK(n73), .RSTB(n57), .Q(n603) );
  SDFFARX1 \ram_di_reg[27]  ( .D(n1656), .SI(ram_di[26]), .SE(test_se), .CLK(
        n71), .RSTB(n21), .Q(ram_di[27]) );
  SDFFARX1 \LatchedTxLength_reg[10]  ( .D(n1118), .SI(n601), .SE(test_se), 
        .CLK(n73), .RSTB(n57), .Q(n602) );
  SDFFARX1 \ram_di_reg[26]  ( .D(n1657), .SI(ram_di[25]), .SE(test_se), .CLK(
        n71), .RSTB(n21), .Q(ram_di[26]) );
  SDFFARX1 \LatchedTxLength_reg[9]  ( .D(n1115), .SI(n600), .SE(test_se), 
        .CLK(n73), .RSTB(n56), .Q(n601) );
  SDFFARX1 \ram_di_reg[25]  ( .D(n1658), .SI(ram_di[24]), .SE(test_se), .CLK(
        n71), .RSTB(n21), .Q(ram_di[25]) );
  SDFFARX1 \LatchedTxLength_reg[8]  ( .D(n1112), .SI(n599), .SE(test_se), 
        .CLK(n73), .RSTB(n56), .Q(n600) );
  SDFFARX1 \ram_di_reg[24]  ( .D(n1659), .SI(ram_di[23]), .SE(test_se), .CLK(
        n71), .RSTB(n21), .Q(ram_di[24]) );
  SDFFARX1 \LatchedTxLength_reg[7]  ( .D(n1109), .SI(n598), .SE(test_se), 
        .CLK(n73), .RSTB(n56), .Q(n599) );
  SDFFARX1 \ram_di_reg[23]  ( .D(n1660), .SI(ram_di[22]), .SE(test_se), .CLK(
        n71), .RSTB(n21), .Q(ram_di[23]) );
  SDFFARX1 \LatchedTxLength_reg[6]  ( .D(n1106), .SI(n597), .SE(test_se), 
        .CLK(n73), .RSTB(n51), .Q(n598) );
  SDFFARX1 \ram_di_reg[22]  ( .D(n1661), .SI(ram_di[21]), .SE(test_se), .CLK(
        n71), .RSTB(n20), .Q(ram_di[22]) );
  SDFFARX1 \LatchedTxLength_reg[5]  ( .D(n1103), .SI(n596), .SE(test_se), 
        .CLK(n73), .RSTB(n51), .Q(n597) );
  SDFFARX1 \ram_di_reg[21]  ( .D(n1662), .SI(ram_di[20]), .SE(test_se), .CLK(
        n71), .RSTB(n20), .Q(ram_di[21]) );
  SDFFARX1 \LatchedTxLength_reg[4]  ( .D(n1100), .SI(n595), .SE(test_se), 
        .CLK(n73), .RSTB(n51), .Q(n596) );
  SDFFARX1 \ram_di_reg[20]  ( .D(n1663), .SI(ram_di[19]), .SE(test_se), .CLK(
        n71), .RSTB(n20), .Q(ram_di[20]) );
  SDFFARX1 \LatchedTxLength_reg[3]  ( .D(n1097), .SI(n594), .SE(test_se), 
        .CLK(n74), .RSTB(n51), .Q(n595) );
  SDFFARX1 \ram_di_reg[19]  ( .D(n1664), .SI(ram_di[18]), .SE(test_se), .CLK(
        n71), .RSTB(n20), .Q(ram_di[19]) );
  SDFFARX1 \LatchedTxLength_reg[2]  ( .D(n1094), .SI(n593), .SE(test_se), 
        .CLK(n74), .RSTB(n51), .Q(n594) );
  SDFFARX1 \ram_di_reg[18]  ( .D(n1665), .SI(ram_di[17]), .SE(test_se), .CLK(
        n71), .RSTB(n20), .Q(ram_di[18]) );
  SDFFARX1 \LatchedTxLength_reg[1]  ( .D(n1091), .SI(n592), .SE(test_se), 
        .CLK(n74), .RSTB(n49), .Q(n593) );
  SDFFARX1 \ram_di_reg[17]  ( .D(n1666), .SI(ram_di[16]), .SE(test_se), .CLK(
        n71), .RSTB(n20), .Q(ram_di[17]) );
  SDFFARX1 \LatchedTxLength_reg[0]  ( .D(n1088), .SI(LatchedRxStartFrm), .SE(
        test_se), .CLK(n74), .RSTB(n49), .Q(n592) );
  SDFFARX1 \ram_di_reg[16]  ( .D(n1667), .SI(ram_di[15]), .SE(test_se), .CLK(
        n71), .RSTB(n20), .Q(ram_di[16]) );
  SDFFARX1 \TxLength_reg[0]  ( .D(n1648), .SI(n589), .SE(test_se), .CLK(n71), 
        .RSTB(n22), .Q(n35), .QN(n720) );
  SDFFARX1 \TxLength_reg[1]  ( .D(n1647), .SI(n35), .SE(test_se), .CLK(n73), 
        .RSTB(n55), .Q(n38), .QN(n721) );
  SDFFARX1 \TxValidBytesLatched_reg[1]  ( .D(n1631), .SI(n655), .SE(test_se), 
        .CLK(n71), .RSTB(n23), .Q(n591), .QN(n991) );
  SDFFARX1 \TxLength_reg[2]  ( .D(n1646), .SI(n38), .SE(test_se), .CLK(n73), 
        .RSTB(n55), .Q(n33), .QN(n707) );
  SDFFARX1 \TxLength_reg[3]  ( .D(n1645), .SI(n33), .SE(test_se), .CLK(n73), 
        .RSTB(n55), .Q(n11), .QN(n708) );
  SDFFARX1 \TxLength_reg[4]  ( .D(n1644), .SI(n11), .SE(test_se), .CLK(n73), 
        .RSTB(n55), .Q(n30), .QN(n709) );
  SDFFARX1 \TxLength_reg[5]  ( .D(n1643), .SI(n30), .SE(test_se), .CLK(n73), 
        .RSTB(n55), .Q(n29), .QN(n710) );
  SDFFARX1 \TxLength_reg[6]  ( .D(n1642), .SI(n29), .SE(test_se), .CLK(n73), 
        .RSTB(n55), .Q(n50), .QN(n711) );
  SDFFARX1 \TxLength_reg[7]  ( .D(n1641), .SI(n50), .SE(test_se), .CLK(n73), 
        .RSTB(n55), .Q(n12), .QN(n712) );
  SDFFARX1 \TxLength_reg[8]  ( .D(n1640), .SI(n12), .SE(test_se), .CLK(n73), 
        .RSTB(n55), .Q(n37), .QN(n713) );
  SDFFARX1 \TxLength_reg[9]  ( .D(n1639), .SI(n37), .SE(test_se), .CLK(n73), 
        .RSTB(n55), .Q(n3), .QN(n714) );
  SDFFARX1 \TxLength_reg[10]  ( .D(n1638), .SI(n3), .SE(test_se), .CLK(n73), 
        .RSTB(n55), .Q(n36), .QN(n715) );
  SDFFARX1 \TxLength_reg[11]  ( .D(n1637), .SI(n36), .SE(test_se), .CLK(n73), 
        .RSTB(n55), .Q(n4), .QN(n716) );
  SDFFARX1 \TxLength_reg[12]  ( .D(n1636), .SI(n4), .SE(test_se), .CLK(n73), 
        .RSTB(n56), .Q(n19), .QN(n717) );
  SDFFARX1 \TxLength_reg[13]  ( .D(n1635), .SI(n19), .SE(test_se), .CLK(n73), 
        .RSTB(n51), .Q(n43), .QN(n718) );
  SDFFARX1 \TxLength_reg[14]  ( .D(n1634), .SI(n43), .SE(test_se), .CLK(n73), 
        .RSTB(n56), .Q(n32), .QN(n719) );
  SDFFARX1 TxStartFrm_wb_reg ( .D(n1626), .SI(n751), .SE(test_se), .CLK(n71), 
        .RSTB(n25), .Q(TxStartFrm_wb), .QN(n993) );
  SDFFARX1 TxStartFrm_sync1_reg ( .D(TxStartFrm_wb), .SI(TxStartFrm), .SE(
        test_se), .CLK(n78), .RSTB(n61), .Q(TxStartFrm_sync1) );
  SDFFARX1 TxStartFrm_sync2_reg ( .D(TxStartFrm_sync1), .SI(TxStartFrm_sync1), 
        .SE(test_se), .CLK(n78), .RSTB(n61), .Q(TxStartFrm_sync2), .QN(n1433)
         );
  SDFFARX1 TxStartFrm_syncb1_reg ( .D(TxStartFrm_sync2), .SI(TxStartFrm_sync2), 
        .SE(test_se), .CLK(n74), .RSTB(n61), .Q(TxStartFrm_syncb1) );
  SDFFARX1 TxStartFrm_syncb2_reg ( .D(TxStartFrm_syncb1), .SI(
        TxStartFrm_syncb1), .SE(test_se), .CLK(n74), .RSTB(n62), .Q(n751), 
        .QN(n723) );
  SDFFARX1 TxStartFrm_reg ( .D(n1625), .SI(TxRetry_wb), .SE(test_se), .CLK(n80), .RSTB(n40), .Q(TxStartFrm) );
  SDFFARX1 \TxByteCnt_reg[0]  ( .D(n1624), .SI(TxB_IRQ), .SE(test_se), .CLK(
        n80), .RSTB(n40), .Q(n693), .QN(n544) );
  SDFFARX1 \TxByteCnt_reg[1]  ( .D(n1623), .SI(n693), .SE(test_se), .CLK(n80), 
        .RSTB(n40), .Q(n694), .QN(n543) );
  SDFFARX1 StartOccured_reg ( .D(n1622), .SI(n636), .SE(test_se), .CLK(n71), 
        .RSTB(n25), .Q(n590), .QN(n994) );
  SDFFARX1 ReadTxDataFromMemory_reg ( .D(n1633), .SI(ReadTxDataFromFifo_tck), 
        .SE(test_se), .CLK(n71), .RSTB(n22), .Q(n760), .QN(n533) );
  SDFFARX1 TxEndFrm_wb_reg ( .D(n1627), .SI(TxEndFrm), .SE(test_se), .CLK(n71), 
        .RSTB(n22), .Q(n589) );
  SDFFARX1 BlockingTxBDRead_reg ( .D(n1580), .SI(n553), .SE(test_se), .CLK(n73), .RSTB(n34), .Q(n555), .QN(n542) );
  SDFFARX1 TxRetryPacket_NotCleared_reg ( .D(n1707), .SI(n650), .SE(test_se), 
        .CLK(n73), .RSTB(n57), .Q(n726), .QN(n541) );
  SDFFARX1 \TxDataLatched_reg[0]  ( .D(n1621), .SI(n694), .SE(test_se), .CLK(
        n80), .RSTB(n40), .Q(n588) );
  SDFFARX1 \TxDataLatched_reg[1]  ( .D(n1620), .SI(n588), .SE(test_se), .CLK(
        n80), .RSTB(n40), .Q(n587) );
  SDFFARX1 \TxDataLatched_reg[2]  ( .D(n1619), .SI(n587), .SE(test_se), .CLK(
        n80), .RSTB(n40), .Q(n586) );
  SDFFARX1 \TxDataLatched_reg[3]  ( .D(n1618), .SI(n586), .SE(test_se), .CLK(
        n80), .RSTB(n40), .Q(n585) );
  SDFFARX1 \TxDataLatched_reg[4]  ( .D(n1617), .SI(n585), .SE(test_se), .CLK(
        n80), .RSTB(n40), .Q(n584) );
  SDFFARX1 \TxDataLatched_reg[5]  ( .D(n1616), .SI(n584), .SE(test_se), .CLK(
        n79), .RSTB(n40), .Q(n583) );
  SDFFARX1 \TxDataLatched_reg[6]  ( .D(n1615), .SI(n583), .SE(test_se), .CLK(
        n79), .RSTB(n40), .Q(n582) );
  SDFFARX1 \TxDataLatched_reg[7]  ( .D(n1614), .SI(n582), .SE(test_se), .CLK(
        n79), .RSTB(n40), .Q(n581) );
  SDFFARX1 \TxDataLatched_reg[8]  ( .D(n1613), .SI(n581), .SE(test_se), .CLK(
        n79), .RSTB(n40), .Q(n580) );
  SDFFARX1 \TxDataLatched_reg[9]  ( .D(n1612), .SI(n580), .SE(test_se), .CLK(
        n78), .RSTB(n57), .Q(n579) );
  SDFFARX1 \TxDataLatched_reg[10]  ( .D(n1611), .SI(n579), .SE(test_se), .CLK(
        n78), .RSTB(n57), .Q(n578) );
  SDFFARX1 \TxDataLatched_reg[11]  ( .D(n1610), .SI(n578), .SE(test_se), .CLK(
        n77), .RSTB(n57), .Q(n577) );
  SDFFARX1 \TxDataLatched_reg[12]  ( .D(n1609), .SI(n577), .SE(test_se), .CLK(
        n77), .RSTB(n57), .Q(n576) );
  SDFFARX1 \TxDataLatched_reg[13]  ( .D(n1608), .SI(n576), .SE(test_se), .CLK(
        n77), .RSTB(n57), .Q(n575) );
  SDFFARX1 \TxDataLatched_reg[14]  ( .D(n1607), .SI(n575), .SE(test_se), .CLK(
        n77), .RSTB(n57), .Q(n574) );
  SDFFARX1 \TxDataLatched_reg[15]  ( .D(n1606), .SI(n574), .SE(test_se), .CLK(
        n77), .RSTB(n58), .Q(n573) );
  SDFFARX1 \TxDataLatched_reg[16]  ( .D(n1605), .SI(n573), .SE(test_se), .CLK(
        n77), .RSTB(n58), .Q(n572) );
  SDFFARX1 \TxDataLatched_reg[17]  ( .D(n1604), .SI(n572), .SE(test_se), .CLK(
        n77), .RSTB(n58), .Q(n571) );
  SDFFARX1 \TxDataLatched_reg[18]  ( .D(n1603), .SI(n571), .SE(test_se), .CLK(
        n77), .RSTB(n58), .Q(n570) );
  SDFFARX1 \TxDataLatched_reg[19]  ( .D(n1602), .SI(n570), .SE(test_se), .CLK(
        n77), .RSTB(n58), .Q(n569) );
  SDFFARX1 \TxDataLatched_reg[20]  ( .D(n1601), .SI(n569), .SE(test_se), .CLK(
        n77), .RSTB(n58), .Q(n568) );
  SDFFARX1 \TxDataLatched_reg[21]  ( .D(n1600), .SI(n568), .SE(test_se), .CLK(
        n77), .RSTB(n58), .Q(n567) );
  SDFFARX1 \TxDataLatched_reg[22]  ( .D(n1599), .SI(n567), .SE(test_se), .CLK(
        n77), .RSTB(n58), .Q(n566) );
  SDFFARX1 \TxDataLatched_reg[23]  ( .D(n1598), .SI(n566), .SE(test_se), .CLK(
        n76), .RSTB(n58), .Q(n565) );
  SDFFARX1 \TxDataLatched_reg[24]  ( .D(n1597), .SI(n565), .SE(test_se), .CLK(
        n76), .RSTB(n58), .Q(n564) );
  SDFFARX1 \TxData_reg[0]  ( .D(n1589), .SI(n557), .SE(test_se), .CLK(n79), 
        .RSTB(n41), .Q(TxData[0]) );
  SDFFARX1 \TxDataLatched_reg[25]  ( .D(n1596), .SI(n564), .SE(test_se), .CLK(
        n76), .RSTB(n58), .Q(n563) );
  SDFFARX1 \TxData_reg[1]  ( .D(n1588), .SI(TxData[0]), .SE(test_se), .CLK(n79), .RSTB(n41), .Q(TxData[1]) );
  SDFFARX1 \TxDataLatched_reg[26]  ( .D(n1595), .SI(n563), .SE(test_se), .CLK(
        n76), .RSTB(n58), .Q(n562) );
  SDFFARX1 \TxData_reg[2]  ( .D(n1587), .SI(TxData[1]), .SE(test_se), .CLK(n79), .RSTB(n41), .Q(TxData[2]) );
  SDFFARX1 \TxDataLatched_reg[27]  ( .D(n1594), .SI(n562), .SE(test_se), .CLK(
        n76), .RSTB(n60), .Q(n561) );
  SDFFARX1 \TxData_reg[3]  ( .D(n1586), .SI(TxData[2]), .SE(test_se), .CLK(n79), .RSTB(n41), .Q(TxData[3]) );
  SDFFARX1 \TxDataLatched_reg[28]  ( .D(n1593), .SI(n561), .SE(test_se), .CLK(
        n76), .RSTB(n60), .Q(n560) );
  SDFFARX1 \TxData_reg[4]  ( .D(n1585), .SI(TxData[3]), .SE(test_se), .CLK(n79), .RSTB(n41), .Q(TxData[4]) );
  SDFFARX1 \TxDataLatched_reg[29]  ( .D(n1592), .SI(n560), .SE(test_se), .CLK(
        n76), .RSTB(n60), .Q(n559) );
  SDFFARX1 \TxData_reg[5]  ( .D(n1584), .SI(TxData[4]), .SE(test_se), .CLK(n79), .RSTB(n41), .Q(TxData[5]) );
  SDFFARX1 \TxDataLatched_reg[30]  ( .D(n1591), .SI(n559), .SE(test_se), .CLK(
        n76), .RSTB(n60), .Q(n558) );
  SDFFARX1 \TxData_reg[6]  ( .D(n1583), .SI(TxData[5]), .SE(test_se), .CLK(n79), .RSTB(n41), .Q(TxData[6]) );
  SDFFARX1 \TxDataLatched_reg[31]  ( .D(n1590), .SI(n558), .SE(test_se), .CLK(
        n76), .RSTB(n60), .Q(n557) );
  SDFFARX1 \TxData_reg[7]  ( .D(n1582), .SI(TxData[6]), .SE(test_se), .CLK(n79), .RSTB(n41), .Q(TxData[7]) );
  SDFFARX1 \TxPointerMSB_reg[31]  ( .D(n1532), .SI(TxPointerMSB[30]), .SE(
        test_se), .CLK(n71), .RSTB(n24), .Q(TxPointerMSB[31]) );
  SDFFARX1 \TxPointerMSB_reg[2]  ( .D(n1561), .SI(n695), .SE(test_se), .CLK(
        n73), .RSTB(n52), .Q(TxPointerMSB[2]) );
  SDFFARX1 \TxPointerMSB_reg[3]  ( .D(n1560), .SI(TxPointerMSB[2]), .SE(
        test_se), .CLK(n73), .RSTB(n52), .Q(TxPointerMSB[3]) );
  SDFFARX1 \TxPointerMSB_reg[4]  ( .D(n1559), .SI(TxPointerMSB[3]), .SE(
        test_se), .CLK(n73), .RSTB(n52), .Q(TxPointerMSB[4]) );
  SDFFARX1 \TxPointerMSB_reg[5]  ( .D(n1558), .SI(TxPointerMSB[4]), .SE(
        test_se), .CLK(n73), .RSTB(n52), .Q(TxPointerMSB[5]) );
  SDFFARX1 \TxPointerMSB_reg[6]  ( .D(n1557), .SI(TxPointerMSB[5]), .SE(
        test_se), .CLK(n73), .RSTB(n52), .Q(TxPointerMSB[6]) );
  SDFFARX1 \TxPointerMSB_reg[7]  ( .D(n1556), .SI(TxPointerMSB[6]), .SE(
        test_se), .CLK(n73), .RSTB(n52), .Q(TxPointerMSB[7]) );
  SDFFARX1 \TxPointerMSB_reg[8]  ( .D(n1555), .SI(TxPointerMSB[7]), .SE(
        test_se), .CLK(n73), .RSTB(n52), .Q(TxPointerMSB[8]) );
  SDFFARX1 \TxPointerMSB_reg[9]  ( .D(n1554), .SI(TxPointerMSB[8]), .SE(
        test_se), .CLK(n73), .RSTB(n52), .Q(TxPointerMSB[9]) );
  SDFFARX1 \TxPointerMSB_reg[10]  ( .D(n1553), .SI(TxPointerMSB[9]), .SE(
        test_se), .CLK(n73), .RSTB(n52), .Q(TxPointerMSB[10]) );
  SDFFARX1 \TxPointerMSB_reg[11]  ( .D(n1552), .SI(TxPointerMSB[10]), .SE(
        test_se), .CLK(n73), .RSTB(n53), .Q(TxPointerMSB[11]) );
  SDFFARX1 \TxPointerMSB_reg[12]  ( .D(n1551), .SI(TxPointerMSB[11]), .SE(
        test_se), .CLK(n73), .RSTB(n53), .Q(TxPointerMSB[12]) );
  SDFFARX1 \TxPointerMSB_reg[13]  ( .D(n1550), .SI(TxPointerMSB[12]), .SE(
        test_se), .CLK(n73), .RSTB(n53), .Q(TxPointerMSB[13]) );
  SDFFARX1 \TxPointerMSB_reg[14]  ( .D(n1549), .SI(TxPointerMSB[13]), .SE(
        test_se), .CLK(n73), .RSTB(n53), .Q(TxPointerMSB[14]) );
  SDFFARX1 \TxPointerMSB_reg[15]  ( .D(n1548), .SI(TxPointerMSB[14]), .SE(
        test_se), .CLK(n73), .RSTB(n53), .Q(TxPointerMSB[15]) );
  SDFFARX1 \TxPointerMSB_reg[16]  ( .D(n1547), .SI(TxPointerMSB[15]), .SE(
        test_se), .CLK(n73), .RSTB(n53), .Q(TxPointerMSB[16]) );
  SDFFARX1 \TxPointerMSB_reg[17]  ( .D(n1546), .SI(TxPointerMSB[16]), .SE(
        test_se), .CLK(n73), .RSTB(n53), .Q(TxPointerMSB[17]) );
  SDFFARX1 \TxPointerMSB_reg[18]  ( .D(n1545), .SI(TxPointerMSB[17]), .SE(
        test_se), .CLK(n73), .RSTB(n53), .Q(TxPointerMSB[18]) );
  SDFFARX1 \TxPointerMSB_reg[19]  ( .D(n1544), .SI(TxPointerMSB[18]), .SE(
        test_se), .CLK(n73), .RSTB(n53), .Q(TxPointerMSB[19]) );
  SDFFARX1 \TxPointerMSB_reg[20]  ( .D(n1543), .SI(TxPointerMSB[19]), .SE(
        test_se), .CLK(n73), .RSTB(n53), .Q(TxPointerMSB[20]) );
  SDFFARX1 \TxPointerMSB_reg[21]  ( .D(n1542), .SI(TxPointerMSB[20]), .SE(
        test_se), .CLK(n73), .RSTB(n53), .Q(TxPointerMSB[21]) );
  SDFFARX1 \TxPointerMSB_reg[22]  ( .D(n1541), .SI(TxPointerMSB[21]), .SE(
        test_se), .CLK(n73), .RSTB(n53), .Q(TxPointerMSB[22]) );
  SDFFARX1 \TxPointerMSB_reg[23]  ( .D(n1540), .SI(TxPointerMSB[22]), .SE(
        test_se), .CLK(n71), .RSTB(n23), .Q(TxPointerMSB[23]) );
  SDFFARX1 \TxPointerMSB_reg[24]  ( .D(n1539), .SI(TxPointerMSB[23]), .SE(
        test_se), .CLK(n71), .RSTB(n24), .Q(TxPointerMSB[24]) );
  SDFFARX1 \TxPointerMSB_reg[25]  ( .D(n1538), .SI(TxPointerMSB[24]), .SE(
        test_se), .CLK(n71), .RSTB(n24), .Q(TxPointerMSB[25]) );
  SDFFARX1 \TxPointerMSB_reg[26]  ( .D(n1537), .SI(TxPointerMSB[25]), .SE(
        test_se), .CLK(n71), .RSTB(n24), .Q(TxPointerMSB[26]) );
  SDFFARX1 \TxPointerMSB_reg[27]  ( .D(n1536), .SI(TxPointerMSB[26]), .SE(
        test_se), .CLK(n71), .RSTB(n24), .Q(TxPointerMSB[27]) );
  SDFFARX1 \TxPointerMSB_reg[28]  ( .D(n1535), .SI(TxPointerMSB[27]), .SE(
        test_se), .CLK(n71), .RSTB(n24), .Q(TxPointerMSB[28]) );
  SDFFARX1 \TxPointerMSB_reg[29]  ( .D(n1534), .SI(TxPointerMSB[28]), .SE(
        test_se), .CLK(n71), .RSTB(n24), .Q(TxPointerMSB[29]) );
  SDFFARX1 \TxPointerMSB_reg[30]  ( .D(n1533), .SI(TxPointerMSB[29]), .SE(
        test_se), .CLK(n71), .RSTB(n24), .Q(TxPointerMSB[30]) );
  SDFFARX1 \RxPointerMSB_reg[31]  ( .D(n1502), .SI(RxPointerMSB[30]), .SE(
        test_se), .CLK(n71), .RSTB(n21), .Q(RxPointerMSB[31]) );
  SDFFARX1 \RxPointerMSB_reg[2]  ( .D(n1531), .SI(n704), .SE(test_se), .CLK(
        n72), .RSTB(n42), .Q(RxPointerMSB[2]) );
  SDFFARX1 \RxPointerMSB_reg[3]  ( .D(n1530), .SI(RxPointerMSB[2]), .SE(
        test_se), .CLK(n74), .RSTB(n62), .Q(RxPointerMSB[3]) );
  SDFFARX1 \RxPointerMSB_reg[4]  ( .D(n1529), .SI(RxPointerMSB[3]), .SE(
        test_se), .CLK(n74), .RSTB(n62), .Q(RxPointerMSB[4]) );
  SDFFARX1 \RxPointerMSB_reg[5]  ( .D(n1528), .SI(RxPointerMSB[4]), .SE(
        test_se), .CLK(n74), .RSTB(n62), .Q(RxPointerMSB[5]) );
  SDFFARX1 \RxPointerMSB_reg[6]  ( .D(n1527), .SI(RxPointerMSB[5]), .SE(
        test_se), .CLK(n74), .RSTB(n62), .Q(RxPointerMSB[6]) );
  SDFFARX1 \RxPointerMSB_reg[7]  ( .D(n1526), .SI(RxPointerMSB[6]), .SE(
        test_se), .CLK(n74), .RSTB(n62), .Q(RxPointerMSB[7]) );
  SDFFARX1 \RxPointerMSB_reg[8]  ( .D(n1525), .SI(RxPointerMSB[7]), .SE(
        test_se), .CLK(n74), .RSTB(n62), .Q(RxPointerMSB[8]) );
  SDFFARX1 \RxPointerMSB_reg[9]  ( .D(n1524), .SI(RxPointerMSB[8]), .SE(
        test_se), .CLK(n74), .RSTB(n62), .Q(RxPointerMSB[9]) );
  SDFFARX1 \RxPointerMSB_reg[10]  ( .D(n1523), .SI(RxPointerMSB[9]), .SE(
        test_se), .CLK(n74), .RSTB(n62), .Q(RxPointerMSB[10]) );
  SDFFARX1 \RxPointerMSB_reg[11]  ( .D(n1522), .SI(RxPointerMSB[10]), .SE(
        test_se), .CLK(n74), .RSTB(n62), .Q(RxPointerMSB[11]) );
  SDFFARX1 \RxPointerMSB_reg[12]  ( .D(n1521), .SI(RxPointerMSB[11]), .SE(
        test_se), .CLK(n74), .RSTB(n62), .Q(RxPointerMSB[12]) );
  SDFFARX1 \RxPointerMSB_reg[13]  ( .D(n1520), .SI(RxPointerMSB[12]), .SE(
        test_se), .CLK(n74), .RSTB(n63), .Q(RxPointerMSB[13]) );
  SDFFARX1 \RxPointerMSB_reg[14]  ( .D(n1519), .SI(RxPointerMSB[13]), .SE(
        test_se), .CLK(n74), .RSTB(n63), .Q(RxPointerMSB[14]) );
  SDFFARX1 \RxPointerMSB_reg[15]  ( .D(n1518), .SI(RxPointerMSB[14]), .SE(
        test_se), .CLK(n74), .RSTB(n49), .Q(RxPointerMSB[15]) );
  SDFFARX1 \RxPointerMSB_reg[16]  ( .D(n1517), .SI(RxPointerMSB[15]), .SE(
        test_se), .CLK(n74), .RSTB(n49), .Q(RxPointerMSB[16]) );
  SDFFARX1 \RxPointerMSB_reg[17]  ( .D(n1516), .SI(RxPointerMSB[16]), .SE(
        test_se), .CLK(n74), .RSTB(n49), .Q(RxPointerMSB[17]) );
  SDFFARX1 \RxPointerMSB_reg[18]  ( .D(n1515), .SI(RxPointerMSB[17]), .SE(
        test_se), .CLK(n74), .RSTB(n49), .Q(RxPointerMSB[18]) );
  SDFFARX1 \RxPointerMSB_reg[19]  ( .D(n1514), .SI(RxPointerMSB[18]), .SE(
        test_se), .CLK(n74), .RSTB(n51), .Q(RxPointerMSB[19]) );
  SDFFARX1 \RxPointerMSB_reg[20]  ( .D(n1513), .SI(RxPointerMSB[19]), .SE(
        test_se), .CLK(n73), .RSTB(n51), .Q(RxPointerMSB[20]) );
  SDFFARX1 \RxPointerMSB_reg[21]  ( .D(n1512), .SI(RxPointerMSB[20]), .SE(
        test_se), .CLK(n73), .RSTB(n51), .Q(RxPointerMSB[21]) );
  SDFFARX1 \RxPointerMSB_reg[22]  ( .D(n1511), .SI(RxPointerMSB[21]), .SE(
        test_se), .CLK(n73), .RSTB(n51), .Q(RxPointerMSB[22]) );
  SDFFARX1 \RxPointerMSB_reg[23]  ( .D(n1510), .SI(RxPointerMSB[22]), .SE(
        test_se), .CLK(n73), .RSTB(n56), .Q(RxPointerMSB[23]) );
  SDFFARX1 \RxPointerMSB_reg[24]  ( .D(n1509), .SI(RxPointerMSB[23]), .SE(
        test_se), .CLK(n73), .RSTB(n56), .Q(RxPointerMSB[24]) );
  SDFFARX1 \RxPointerMSB_reg[25]  ( .D(n1508), .SI(RxPointerMSB[24]), .SE(
        test_se), .CLK(n73), .RSTB(n56), .Q(RxPointerMSB[25]) );
  SDFFARX1 \RxPointerMSB_reg[26]  ( .D(n1507), .SI(RxPointerMSB[25]), .SE(
        test_se), .CLK(n73), .RSTB(n56), .Q(RxPointerMSB[26]) );
  SDFFARX1 \RxPointerMSB_reg[27]  ( .D(n1506), .SI(RxPointerMSB[26]), .SE(
        test_se), .CLK(n73), .RSTB(n56), .Q(RxPointerMSB[27]) );
  SDFFARX1 \RxPointerMSB_reg[28]  ( .D(n1505), .SI(RxPointerMSB[27]), .SE(
        test_se), .CLK(n73), .RSTB(n56), .Q(RxPointerMSB[28]) );
  SDFFARX1 \RxPointerMSB_reg[29]  ( .D(n1504), .SI(RxPointerMSB[28]), .SE(
        test_se), .CLK(n73), .RSTB(n56), .Q(RxPointerMSB[29]) );
  SDFFARX1 \RxPointerMSB_reg[30]  ( .D(n1503), .SI(RxPointerMSB[29]), .SE(
        test_se), .CLK(n71), .RSTB(n21), .Q(RxPointerMSB[30]) );
  SDFFARX1 \m_wb_adr_o_reg[29]  ( .D(n1472), .SI(m_wb_adr_o[28]), .SE(test_se), 
        .CLK(n72), .RSTB(n46), .Q(m_wb_adr_o[29]) );
  SDFFARX1 \m_wb_adr_o_reg[0]  ( .D(n1501), .SI(n728), .SE(test_se), .CLK(n72), 
        .RSTB(n42), .Q(m_wb_adr_o[0]) );
  SDFFARX1 \m_wb_adr_o_reg[1]  ( .D(n1500), .SI(m_wb_adr_o[0]), .SE(test_se), 
        .CLK(n72), .RSTB(n42), .Q(m_wb_adr_o[1]) );
  SDFFARX1 \m_wb_adr_o_reg[2]  ( .D(n1499), .SI(m_wb_adr_o[1]), .SE(test_se), 
        .CLK(n72), .RSTB(n42), .Q(m_wb_adr_o[2]) );
  SDFFARX1 \m_wb_adr_o_reg[3]  ( .D(n1498), .SI(m_wb_adr_o[2]), .SE(test_se), 
        .CLK(n72), .RSTB(n44), .Q(m_wb_adr_o[3]) );
  SDFFARX1 \m_wb_adr_o_reg[4]  ( .D(n1497), .SI(m_wb_adr_o[3]), .SE(test_se), 
        .CLK(n72), .RSTB(n44), .Q(m_wb_adr_o[4]) );
  SDFFARX1 \m_wb_adr_o_reg[5]  ( .D(n1496), .SI(m_wb_adr_o[4]), .SE(test_se), 
        .CLK(n72), .RSTB(n44), .Q(m_wb_adr_o[5]) );
  SDFFARX1 \m_wb_adr_o_reg[6]  ( .D(n1495), .SI(m_wb_adr_o[5]), .SE(test_se), 
        .CLK(n72), .RSTB(n44), .Q(m_wb_adr_o[6]) );
  SDFFARX1 \m_wb_adr_o_reg[7]  ( .D(n1494), .SI(m_wb_adr_o[6]), .SE(test_se), 
        .CLK(n72), .RSTB(n44), .Q(m_wb_adr_o[7]) );
  SDFFARX1 \m_wb_adr_o_reg[8]  ( .D(n1493), .SI(m_wb_adr_o[7]), .SE(test_se), 
        .CLK(n72), .RSTB(n44), .Q(m_wb_adr_o[8]) );
  SDFFARX1 \m_wb_adr_o_reg[9]  ( .D(n1492), .SI(m_wb_adr_o[8]), .SE(test_se), 
        .CLK(n72), .RSTB(n44), .Q(m_wb_adr_o[9]) );
  SDFFARX1 \m_wb_adr_o_reg[10]  ( .D(n1491), .SI(m_wb_adr_o[9]), .SE(test_se), 
        .CLK(n72), .RSTB(n44), .Q(m_wb_adr_o[10]) );
  SDFFARX1 \m_wb_adr_o_reg[11]  ( .D(n1490), .SI(m_wb_adr_o[10]), .SE(test_se), 
        .CLK(n72), .RSTB(n44), .Q(m_wb_adr_o[11]) );
  SDFFARX1 \m_wb_adr_o_reg[12]  ( .D(n1489), .SI(m_wb_adr_o[11]), .SE(test_se), 
        .CLK(n72), .RSTB(n44), .Q(m_wb_adr_o[12]) );
  SDFFARX1 \m_wb_adr_o_reg[13]  ( .D(n1488), .SI(m_wb_adr_o[12]), .SE(test_se), 
        .CLK(n72), .RSTB(n44), .Q(m_wb_adr_o[13]) );
  SDFFARX1 \m_wb_adr_o_reg[14]  ( .D(n1487), .SI(m_wb_adr_o[13]), .SE(test_se), 
        .CLK(n72), .RSTB(n44), .Q(m_wb_adr_o[14]) );
  SDFFARX1 \m_wb_adr_o_reg[15]  ( .D(n1486), .SI(m_wb_adr_o[14]), .SE(test_se), 
        .CLK(n72), .RSTB(n45), .Q(m_wb_adr_o[15]) );
  SDFFARX1 \m_wb_adr_o_reg[16]  ( .D(n1485), .SI(m_wb_adr_o[15]), .SE(test_se), 
        .CLK(n72), .RSTB(n45), .Q(m_wb_adr_o[16]) );
  SDFFARX1 \m_wb_adr_o_reg[17]  ( .D(n1484), .SI(m_wb_adr_o[16]), .SE(test_se), 
        .CLK(n72), .RSTB(n45), .Q(m_wb_adr_o[17]) );
  SDFFARX1 \m_wb_adr_o_reg[18]  ( .D(n1483), .SI(m_wb_adr_o[17]), .SE(test_se), 
        .CLK(n72), .RSTB(n45), .Q(m_wb_adr_o[18]) );
  SDFFARX1 \m_wb_adr_o_reg[19]  ( .D(n1482), .SI(m_wb_adr_o[18]), .SE(test_se), 
        .CLK(n72), .RSTB(n45), .Q(m_wb_adr_o[19]) );
  SDFFARX1 \m_wb_adr_o_reg[20]  ( .D(n1481), .SI(m_wb_adr_o[19]), .SE(test_se), 
        .CLK(n72), .RSTB(n45), .Q(m_wb_adr_o[20]) );
  SDFFARX1 \m_wb_adr_o_reg[21]  ( .D(n1480), .SI(m_wb_adr_o[20]), .SE(test_se), 
        .CLK(n72), .RSTB(n45), .Q(m_wb_adr_o[21]) );
  SDFFARX1 \m_wb_adr_o_reg[22]  ( .D(n1479), .SI(m_wb_adr_o[21]), .SE(test_se), 
        .CLK(n72), .RSTB(n45), .Q(m_wb_adr_o[22]) );
  SDFFARX1 \m_wb_adr_o_reg[23]  ( .D(n1478), .SI(m_wb_adr_o[22]), .SE(test_se), 
        .CLK(n72), .RSTB(n45), .Q(m_wb_adr_o[23]) );
  SDFFARX1 \m_wb_adr_o_reg[24]  ( .D(n1477), .SI(m_wb_adr_o[23]), .SE(test_se), 
        .CLK(n72), .RSTB(n45), .Q(m_wb_adr_o[24]) );
  SDFFARX1 \m_wb_adr_o_reg[25]  ( .D(n1476), .SI(m_wb_adr_o[24]), .SE(test_se), 
        .CLK(n72), .RSTB(n45), .Q(m_wb_adr_o[25]) );
  SDFFARX1 \m_wb_adr_o_reg[26]  ( .D(n1475), .SI(m_wb_adr_o[25]), .SE(test_se), 
        .CLK(n72), .RSTB(n45), .Q(m_wb_adr_o[26]) );
  SDFFARX1 \m_wb_adr_o_reg[27]  ( .D(n1474), .SI(m_wb_adr_o[26]), .SE(test_se), 
        .CLK(n72), .RSTB(n46), .Q(m_wb_adr_o[27]) );
  SDFFARX1 \m_wb_adr_o_reg[28]  ( .D(n1473), .SI(m_wb_adr_o[27]), .SE(test_se), 
        .CLK(n72), .RSTB(n46), .Q(m_wb_adr_o[28]) );
  SDFFARX1 RxStatusWriteLatched_syncb2_reg ( .D(RxStatusWriteLatched_syncb1), 
        .SI(RxStatusWriteLatched_syncb1), .SE(test_se), .CLK(n74), .RSTB(n65), 
        .Q(n756), .QN(n860) );
  SDFFARX1 RxStatusWriteLatched_reg ( .D(n1471), .SI(n665), .SE(test_se), 
        .CLK(n74), .RSTB(n64), .Q(RxStatusWriteLatched) );
  SDFFARX1 RxStatusWriteLatched_sync1_reg ( .D(RxStatusWriteLatched), .SI(
        RxStatusWriteLatched), .SE(test_se), .CLK(n84), .RSTB(n64), .Q(
        RxStatusWriteLatched_sync1) );
  SDFFARX1 RxStatusWriteLatched_sync2_reg ( .D(RxStatusWriteLatched_sync1), 
        .SI(RxStatusWriteLatched_sync1), .SE(test_se), .CLK(n84), .RSTB(n64), 
        .Q(RxStatusWriteLatched_sync2) );
  SDFFARX1 RxStatusWriteLatched_syncb1_reg ( .D(RxStatusWriteLatched_sync2), 
        .SI(RxStatusWriteLatched_sync2), .SE(test_se), .CLK(n74), .RSTB(n65), 
        .Q(RxStatusWriteLatched_syncb1) );
  SDFFARX1 TxB_IRQ_reg ( .D(N1258), .SI(n733), .SE(test_se), .CLK(n74), .RSTB(
        n34), .Q(TxB_IRQ) );
  SDFFARX1 TxE_IRQ_reg ( .D(N1261), .SI(TxDone_wb), .SE(test_se), .CLK(n74), 
        .RSTB(n34), .Q(TxE_IRQ) );
  SDFFARX1 RxB_IRQ_reg ( .D(N1265), .SI(n637), .SE(test_se), .CLK(n71), .RSTB(
        n25), .Q(RxB_IRQ) );
  SDFFARX1 RxE_IRQ_reg ( .D(N1268), .SI(RxDataLatched2[31]), .SE(test_se), 
        .CLK(n73), .RSTB(n48), .Q(RxE_IRQ) );
  SDFFX1 Busy_IRQ_syncb2_reg ( .D(Busy_IRQ_syncb1), .SI(Busy_IRQ_syncb1), .SE(
        test_se), .CLK(n88), .Q(n764), .QN(n1469) );
  SDFFARX1 Busy_IRQ_rck_reg ( .D(n1470), .SI(BlockingTxStatusWrite_sync3), 
        .SE(test_se), .CLK(n81), .RSTB(n22), .Q(Busy_IRQ_rck) );
  SDFFX1 Busy_IRQ_sync1_reg ( .D(Busy_IRQ_rck), .SI(Busy_IRQ_rck), .SE(test_se), .CLK(n75), .Q(Busy_IRQ_sync1) );
  SDFFX1 Busy_IRQ_sync2_reg ( .D(Busy_IRQ_sync1), .SI(Busy_IRQ_sync1), .SE(
        test_se), .CLK(n75), .Q(Busy_IRQ_sync2), .QN(n1468) );
  SDFFX1 Busy_IRQ_sync3_reg ( .D(Busy_IRQ_sync2), .SI(Busy_IRQ_sync2), .SE(
        test_se), .CLK(n75), .Q(Busy_IRQ_sync3) );
  SDFFX1 Busy_IRQ_syncb1_reg ( .D(Busy_IRQ_sync2), .SI(Busy_IRQ_sync3), .SE(
        test_se), .CLK(n88), .Q(Busy_IRQ_syncb1) );
  eth_spram_256x32_test_1 bd_ram ( .clk(n71), .rst(Reset), .ce(1'b1), .we(
        ram_we), .oe(ram_oe), .addr(ram_addr), .di(ram_di), .do(WB_DAT_O), 
        .test_si8(test_si8), .test_si7(test_si7), .test_si6(test_si6), 
        .test_si5(test_si5), .test_si4(test_si4), .test_si3(test_si3), 
        .test_si2(test_si2), .test_si1(WriteRxDataToFifo), .test_so8(n742), 
        .test_so7(test_so7), .test_so6(test_so6), .test_so5(test_so5), 
        .test_so4(test_so4), .test_so3(test_so3), .test_so2(test_so2), 
        .test_so1(test_so1), .test_se(test_se) );
  eth_fifo_DATA_WIDTH32_DEPTH16_CNT_WIDTH5_test_0 tx_fifo ( .data_in(
        m_wb_dat_i), .data_out(TxData_wb), .clk(n70), .reset(Reset), .write(
        n767), .read(_1_net_), .clear(n1188), .almost_full(TxBufferAlmostFull), 
        .full(TxBufferFull), .almost_empty(TxBufferAlmostEmpty), .empty(
        TxBufferEmpty), .cnt({txfifo_cnt[4:2], SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1}), .eth_top_test_point_11887_in(
        eth_top_test_point_11887_in), .test_si(tx_burst_en), .test_so(n738), 
        .test_se(test_se) );
  eth_fifo_DATA_WIDTH32_DEPTH16_CNT_WIDTH5_test_1 rx_fifo ( .data_in(
        RxDataLatched2), .data_out(m_wb_dat_o), .clk(n70), .reset(Reset), 
        .write(_2_net_), .read(n1429), .clear(RxFifoReset), .full(RxBufferFull), .almost_empty(RxBufferAlmostEmpty), .empty(RxBufferEmpty), .cnt(rxfifo_cnt), 
        .eth_top_test_point_11887_in(eth_top_test_point_11887_in), .test_si2(
        n738), .test_si1(rx_burst_en), .test_so1(n739), .test_se(test_se) );
  eth_wishbone_DW01_inc_0 add_1924 ( .A(RxPointerMSB), .SUM({N1027, N1026, 
        N1025, N1024, N1023, N1022, N1021, N1020, N1019, N1018, N1017, N1016, 
        N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, 
        N1005, N1004, N1003, N1002, N1001, N1000, N999, N998}) );
  eth_wishbone_DW01_inc_1 r272 ( .A(m_wb_adr_o), .SUM({N680, N679, N678, N677, 
        N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, 
        N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, 
        N652, N651}) );
  eth_wishbone_DW01_inc_2 add_915 ( .A(TxPointerMSB), .SUM({N379, N378, N377, 
        N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, 
        N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, 
        N352, N351, N350}) );
  eth_wishbone_DW01_inc_3 add_1363 ( .A(TxBDAddress), .SUM({N806, N805, N804, 
        N803, N802, N801, N800}) );
  eth_wishbone_DW01_inc_4 add_1364 ( .A(RxBDAddress), .SUM({N813, N812, N811, 
        N810, N809, N808, N807}) );
  NBUFFX2 U3 ( .INP(n17), .Z(n45) );
  NBUFFX2 U4 ( .INP(n18), .Z(n44) );
  NBUFFX2 U5 ( .INP(n18), .Z(n53) );
  NBUFFX2 U6 ( .INP(n16), .Z(n58) );
  NBUFFX2 U7 ( .INP(n15), .Z(n40) );
  NBUFFX2 U8 ( .INP(n17), .Z(n56) );
  NBUFFX2 U9 ( .INP(n16), .Z(n47) );
  NBUFFX2 U10 ( .INP(n15), .Z(n52) );
  NBUFFX2 U11 ( .INP(n17), .Z(n55) );
  NBUFFX2 U12 ( .INP(n18), .Z(n66) );
  NBUFFX2 U13 ( .INP(n15), .Z(n67) );
  INVX0 U14 ( .INP(eth_top_test_point_11887_in), .ZN(n15) );
  INVX0 U15 ( .INP(eth_top_test_point_11887_in), .ZN(n16) );
  INVX0 U16 ( .INP(eth_top_test_point_11887_in), .ZN(n17) );
  INVX0 U17 ( .INP(eth_top_test_point_11887_in), .ZN(n18) );
  INVX2 U18 ( .INP(n94), .ZN(n111) );
  NOR2X1 U19 ( .IN1(n378), .IN2(n377), .QN(n400) );
  INVX2 U20 ( .INP(n124), .ZN(n1188) );
  NOR2X1 U21 ( .IN1(n1464), .IN2(SyncRxStartFrm_q2), .QN(RxFifoReset) );
  NBUFFX2 U22 ( .INP(n15), .Z(n68) );
  NBUFFX2 U23 ( .INP(n16), .Z(n62) );
  NBUFFX2 U24 ( .INP(n17), .Z(n21) );
  NBUFFX2 U25 ( .INP(n18), .Z(n64) );
  NBUFFX2 U26 ( .INP(n15), .Z(n24) );
  NBUFFX2 U27 ( .INP(n16), .Z(n65) );
  NBUFFX2 U28 ( .INP(n17), .Z(n25) );
  NBUFFX2 U29 ( .INP(n18), .Z(n61) );
  NBUFFX2 U30 ( .INP(n15), .Z(n57) );
  NBUFFX2 U31 ( .INP(n16), .Z(n49) );
  NBUFFX2 U32 ( .INP(n17), .Z(n34) );
  NBUFFX2 U33 ( .INP(n18), .Z(n20) );
  NBUFFX2 U34 ( .INP(n15), .Z(n51) );
  NBUFFX2 U35 ( .INP(n16), .Z(n48) );
  NBUFFX2 U36 ( .INP(n17), .Z(n63) );
  NBUFFX2 U37 ( .INP(n18), .Z(n27) );
  NBUFFX2 U38 ( .INP(n15), .Z(n31) );
  NBUFFX2 U39 ( .INP(n16), .Z(n60) );
  NBUFFX2 U40 ( .INP(n17), .Z(n42) );
  NBUFFX2 U41 ( .INP(n18), .Z(n41) );
  NBUFFX2 U42 ( .INP(n15), .Z(n23) );
  NBUFFX2 U43 ( .INP(n16), .Z(n22) );
  NBUFFX2 U44 ( .INP(n17), .Z(n39) );
  NBUFFX2 U45 ( .INP(n18), .Z(n46) );
  NBUFFX2 U46 ( .INP(n15), .Z(n26) );
  NBUFFX2 U47 ( .INP(n16), .Z(n69) );
  DELLN1X2 U48 ( .INP(MRxClk), .Z(n86) );
  DELLN1X2 U49 ( .INP(MRxClk), .Z(n84) );
  DELLN1X2 U50 ( .INP(MRxClk), .Z(n82) );
  DELLN1X2 U51 ( .INP(MRxClk), .Z(n83) );
  NBUFFX4 U52 ( .INP(MRxClk), .Z(n88) );
  NBUFFX2 U53 ( .INP(MTxClk), .Z(n77) );
  NBUFFX2 U54 ( .INP(MTxClk), .Z(n79) );
  NBUFFX2 U55 ( .INP(MTxClk), .Z(n76) );
  NBUFFX2 U56 ( .INP(MTxClk), .Z(n80) );
  NBUFFX2 U57 ( .INP(MTxClk), .Z(n78) );
  NBUFFX2 U58 ( .INP(WB_CLK_I), .Z(n75) );
  DELLN1X2 U59 ( .INP(WB_CLK_I), .Z(n70) );
  DELLN1X2 U60 ( .INP(WB_CLK_I), .Z(n71) );
  DELLN1X2 U61 ( .INP(WB_CLK_I), .Z(n72) );
  DELLN1X2 U62 ( .INP(WB_CLK_I), .Z(n73) );
  DELLN1X2 U63 ( .INP(WB_CLK_I), .Z(n74) );
  DELLN2X2 U64 ( .INP(MRxClk), .Z(n81) );
  DELLN2X2 U65 ( .INP(MRxClk), .Z(n85) );
  DELLN2X2 U66 ( .INP(MRxClk), .Z(n87) );
  AO21X1 U67 ( .IN1(n641), .IN2(n89), .IN3(n90), .Q(ram_we[3]) );
  AO21X1 U68 ( .IN1(n642), .IN2(n89), .IN3(n90), .Q(ram_we[2]) );
  AO21X1 U69 ( .IN1(n643), .IN2(n89), .IN3(n90), .Q(ram_we[1]) );
  AO21X1 U70 ( .IN1(n644), .IN2(n89), .IN3(n90), .Q(ram_we[0]) );
  NAND2X0 U71 ( .IN1(n91), .IN2(n92), .QN(n90) );
  NAND4X0 U72 ( .IN1(n93), .IN2(n94), .IN3(n95), .IN4(n96), .QN(ram_oe) );
  AOI21X1 U73 ( .IN1(n89), .IN2(n608), .IN3(n97), .QN(n96) );
  NOR4X0 U74 ( .IN1(TxDone), .IN2(n98), .IN3(n99), .IN4(n100), .QN(n1806) );
  NOR2X0 U75 ( .IN1(TxUsedData), .IN2(n686), .QN(n99) );
  OA21X1 U76 ( .IN1(RxStartFrm), .IN2(LatchedRxStartFrm), .IN3(n1464), .Q(
        n1805) );
  NAND2X0 U77 ( .IN1(n101), .IN2(n102), .QN(n1804) );
  NAND3X0 U78 ( .IN1(n103), .IN2(n685), .IN3(n104), .QN(n102) );
  OA21X1 U79 ( .IN1(RxAbort), .IN2(RxAbortLatched), .IN3(n842), .Q(n1803) );
  OA21X1 U80 ( .IN1(n105), .IN2(n657), .IN3(n92), .Q(n1802) );
  AND3X1 U81 ( .IN1(n59), .IN2(WriteRxDataToFifoSync2), .IN3(RxBufferFull), 
        .Q(n105) );
  AO221X1 U82 ( .IN1(ram_di[31]), .IN2(n106), .IN3(WB_DAT_I[31]), .IN4(n107), 
        .IN5(n108), .Q(n1801) );
  AO22X1 U83 ( .IN1(n607), .IN2(n109), .IN3(n684), .IN4(n110), .Q(n108) );
  AO22X1 U84 ( .IN1(WB_DAT_O[31]), .IN2(n111), .IN3(n112), .IN4(n54), .Q(n1800) );
  AO21X1 U85 ( .IN1(n113), .IN2(n32), .IN3(n114), .Q(n112) );
  NAND2X0 U86 ( .IN1(n115), .IN2(n116), .QN(n1799) );
  NAND4X0 U87 ( .IN1(n541), .IN2(n117), .IN3(n747), .IN4(n118), .QN(n116) );
  OR3X1 U88 ( .IN1(TxBufferAlmostFull), .IN2(n119), .IN3(n120), .Q(n118) );
  NOR4X0 U89 ( .IN1(n121), .IN2(n30), .IN3(n122), .IN4(n11), .QN(n120) );
  NAND2X0 U90 ( .IN1(n721), .IN2(n720), .QN(n121) );
  NAND4X0 U91 ( .IN1(n534), .IN2(n653), .IN3(n123), .IN4(n124), .QN(n115) );
  AO22X1 U92 ( .IN1(n125), .IN2(n126), .IN3(tx_burst_cnt[2]), .IN4(n127), .Q(
        n1798) );
  MUX21X1 U93 ( .IN1(n128), .IN2(n129), .S(n130), .Q(n1797) );
  NOR2X0 U94 ( .IN1(n131), .IN2(n6), .QN(n129) );
  NOR3X0 U95 ( .IN1(n132), .IN2(tx_burst_cnt[2]), .IN3(n5), .QN(n131) );
  AOI221X1 U96 ( .IN1(txfifo_cnt[3]), .IN2(txfifo_cnt[2]), .IN3(n133), .IN4(
        n134), .IN5(txfifo_cnt[4]), .QN(n128) );
  AO21X1 U97 ( .IN1(n708), .IN2(n135), .IN3(n709), .Q(n134) );
  AO21X1 U98 ( .IN1(n721), .IN2(n720), .IN3(n707), .Q(n135) );
  MUX21X1 U99 ( .IN1(n136), .IN2(n649), .S(n137), .Q(n1796) );
  AOI21X1 U100 ( .IN1(n1452), .IN2(n696), .IN3(n730), .QN(n137) );
  NAND2X0 U101 ( .IN1(n696), .IN2(n1452), .QN(n136) );
  MUX21X1 U102 ( .IN1(n138), .IN2(N837), .S(n747), .Q(n1795) );
  AO21X1 U103 ( .IN1(n746), .IN2(n731), .IN3(n139), .Q(n1794) );
  INVX0 U104 ( .INP(n140), .ZN(n139) );
  AO22X1 U105 ( .IN1(n731), .IN2(n733), .IN3(n745), .IN4(n725), .Q(n1793) );
  AO22X1 U106 ( .IN1(n93), .IN2(n645), .IN3(n141), .IN4(r_TxEn), .Q(n1792) );
  NOR2X0 U107 ( .IN1(n733), .IN2(n142), .QN(n141) );
  AO21X1 U108 ( .IN1(n106), .IN2(TxEn), .IN3(n109), .Q(n1791) );
  AO21X1 U109 ( .IN1(n106), .IN2(RxEn), .IN3(n110), .Q(n1790) );
  MUX21X1 U110 ( .IN1(n92), .IN2(n143), .S(n687), .Q(n1789) );
  AND3X1 U111 ( .IN1(n1429), .IN2(n609), .IN3(RxBufferAlmostEmpty), .Q(n143)
         );
  OA221X1 U112 ( .IN1(n144), .IN2(n640), .IN3(n765), .IN4(r_RxEn), .IN5(n145), 
        .Q(n1788) );
  OA21X1 U113 ( .IN1(n676), .IN2(RxAbortSync3), .IN3(n687), .Q(n145) );
  AO22X1 U114 ( .IN1(n535), .IN2(n697), .IN3(n8), .IN4(n146), .Q(n1787) );
  AO21X1 U115 ( .IN1(n532), .IN2(RxAbortSync3), .IN3(n147), .Q(n146) );
  INVX0 U116 ( .INP(n148), .ZN(n147) );
  AO222X1 U117 ( .IN1(r_TxBDNum[0]), .IN2(n149), .IN3(n148), .IN4(
        RxBDAddress[1]), .IN5(N807), .IN6(n150), .Q(n1786) );
  AO222X1 U118 ( .IN1(r_TxBDNum[1]), .IN2(n149), .IN3(n148), .IN4(
        RxBDAddress[2]), .IN5(N808), .IN6(n150), .Q(n1785) );
  AO222X1 U119 ( .IN1(r_TxBDNum[2]), .IN2(n149), .IN3(n148), .IN4(
        RxBDAddress[3]), .IN5(N809), .IN6(n150), .Q(n1784) );
  AO222X1 U120 ( .IN1(r_TxBDNum[3]), .IN2(n149), .IN3(n148), .IN4(
        RxBDAddress[4]), .IN5(N810), .IN6(n150), .Q(n1783) );
  AO222X1 U121 ( .IN1(r_TxBDNum[4]), .IN2(n149), .IN3(n148), .IN4(
        RxBDAddress[5]), .IN5(N811), .IN6(n150), .Q(n1782) );
  AO222X1 U122 ( .IN1(r_TxBDNum[5]), .IN2(n149), .IN3(n148), .IN4(
        RxBDAddress[6]), .IN5(N812), .IN6(n150), .Q(n1781) );
  AO222X1 U123 ( .IN1(r_TxBDNum[6]), .IN2(n149), .IN3(n148), .IN4(
        RxBDAddress[7]), .IN5(N813), .IN6(n150), .Q(n1780) );
  NOR3X0 U124 ( .IN1(n151), .IN2(n638), .IN3(n92), .QN(n150) );
  NOR2X0 U125 ( .IN1(n151), .IN2(n152), .QN(n148) );
  AO21X1 U126 ( .IN1(n638), .IN2(n152), .IN3(n151), .Q(n149) );
  AND2X1 U127 ( .IN1(r_RxEn), .IN2(n765), .Q(n151) );
  AO22X1 U128 ( .IN1(n697), .IN2(n637), .IN3(n722), .IN4(n153), .Q(n1779) );
  NOR2X0 U129 ( .IN1(n1429), .IN2(n154), .QN(n1778) );
  INVX0 U130 ( .INP(n155), .ZN(n154) );
  MUX21X1 U131 ( .IN1(n704), .IN2(WB_DAT_O[1]), .S(n144), .Q(n155) );
  MUX21X1 U132 ( .IN1(n625), .IN2(RxData[0]), .S(n156), .Q(n1777) );
  MUX21X1 U133 ( .IN1(n624), .IN2(RxData[7]), .S(n156), .Q(n1776) );
  MUX21X1 U134 ( .IN1(n623), .IN2(RxData[6]), .S(n156), .Q(n1775) );
  MUX21X1 U135 ( .IN1(n622), .IN2(RxData[5]), .S(n156), .Q(n1774) );
  MUX21X1 U136 ( .IN1(n621), .IN2(RxData[4]), .S(n156), .Q(n1773) );
  MUX21X1 U137 ( .IN1(n620), .IN2(RxData[3]), .S(n156), .Q(n1772) );
  MUX21X1 U138 ( .IN1(n619), .IN2(RxData[2]), .S(n156), .Q(n1771) );
  MUX21X1 U139 ( .IN1(n618), .IN2(RxData[1]), .S(n156), .Q(n1770) );
  AOI221X1 U140 ( .IN1(n157), .IN2(n702), .IN3(n158), .IN4(n159), .IN5(n160), 
        .QN(n156) );
  MUX21X1 U141 ( .IN1(n618), .IN2(RxDataLatched2[25]), .S(n161), .Q(n1769) );
  NAND2X0 U142 ( .IN1(n162), .IN2(n163), .QN(n1768) );
  NAND3X0 U143 ( .IN1(n164), .IN2(n635), .IN3(n165), .QN(n163) );
  NOR2X0 U144 ( .IN1(n1429), .IN2(n166), .QN(n1767) );
  MUX21X1 U145 ( .IN1(n549), .IN2(n167), .S(n144), .Q(n166) );
  INVX0 U146 ( .INP(WB_DAT_O[0]), .ZN(n167) );
  AO21X1 U147 ( .IN1(n168), .IN2(n158), .IN3(n169), .Q(n1766) );
  MUX21X1 U148 ( .IN1(n170), .IN2(n171), .S(n985), .Q(n169) );
  NOR2X0 U149 ( .IN1(n548), .IN2(n172), .QN(n171) );
  MUX21X1 U150 ( .IN1(n173), .IN2(n548), .S(n174), .Q(n170) );
  NOR2X0 U151 ( .IN1(n168), .IN2(n175), .QN(n173) );
  OA21X1 U152 ( .IN1(n176), .IN2(n177), .IN3(n104), .Q(n1765) );
  NOR2X0 U153 ( .IN1(n679), .IN2(WriteRxDataToFifoSync2), .QN(n176) );
  NOR2X0 U154 ( .IN1(RxAbort), .IN2(n178), .QN(n1764) );
  OA22X1 U155 ( .IN1(n847), .IN2(n179), .IN3(n161), .IN4(n180), .Q(n178) );
  INVX0 U156 ( .INP(n181), .ZN(n180) );
  NOR2X0 U157 ( .IN1(n848), .IN2(n849), .QN(n179) );
  AO21X1 U158 ( .IN1(n168), .IN2(n549), .IN3(n182), .Q(n1763) );
  MUX21X1 U159 ( .IN1(n183), .IN2(n174), .S(n548), .Q(n182) );
  NOR3X0 U160 ( .IN1(n175), .IN2(n168), .IN3(n174), .QN(n183) );
  INVX0 U161 ( .INP(n172), .ZN(n174) );
  NAND3X0 U162 ( .IN1(n184), .IN2(n185), .IN3(n186), .QN(n172) );
  NAND2X0 U163 ( .IN1(n552), .IN2(n187), .QN(n185) );
  NOR2X0 U164 ( .IN1(n175), .IN2(n184), .QN(n168) );
  OA21X1 U165 ( .IN1(n181), .IN2(n636), .IN3(n186), .Q(n1762) );
  INVX0 U166 ( .INP(n175), .ZN(n186) );
  NAND2X0 U167 ( .IN1(n847), .IN2(n104), .QN(n175) );
  NAND2X0 U168 ( .IN1(n552), .IN2(n188), .QN(n181) );
  NAND4X0 U169 ( .IN1(RxEndFrm), .IN2(n189), .IN3(RxValid), .IN4(n685), .QN(
        n188) );
  OA21X1 U170 ( .IN1(n190), .IN2(n191), .IN3(n104), .Q(n1761) );
  INVX0 U171 ( .INP(RxAbort), .ZN(n104) );
  AOI21X1 U172 ( .IN1(n636), .IN2(n189), .IN3(n552), .QN(n191) );
  NOR3X0 U173 ( .IN1(n103), .IN2(n189), .IN3(n187), .QN(n190) );
  INVX0 U174 ( .INP(RxEndFrm), .ZN(n103) );
  MUX21X1 U175 ( .IN1(n625), .IN2(RxDataLatched2[24]), .S(n161), .Q(n1760) );
  MUX21X1 U176 ( .IN1(n619), .IN2(RxDataLatched2[26]), .S(n161), .Q(n1759) );
  MUX21X1 U177 ( .IN1(n620), .IN2(RxDataLatched2[27]), .S(n161), .Q(n1758) );
  MUX21X1 U178 ( .IN1(n621), .IN2(RxDataLatched2[28]), .S(n161), .Q(n1757) );
  MUX21X1 U179 ( .IN1(n622), .IN2(RxDataLatched2[29]), .S(n161), .Q(n1756) );
  MUX21X1 U180 ( .IN1(n623), .IN2(RxDataLatched2[30]), .S(n161), .Q(n1755) );
  MUX21X1 U181 ( .IN1(n624), .IN2(RxDataLatched2[31]), .S(n161), .Q(n1754) );
  MUX21X1 U182 ( .IN1(n617), .IN2(RxData[0]), .S(n192), .Q(n1753) );
  MUX21X1 U183 ( .IN1(n616), .IN2(RxData[1]), .S(n192), .Q(n1752) );
  MUX21X1 U184 ( .IN1(n615), .IN2(RxData[2]), .S(n192), .Q(n1751) );
  MUX21X1 U185 ( .IN1(n614), .IN2(RxData[3]), .S(n192), .Q(n1750) );
  MUX21X1 U186 ( .IN1(n613), .IN2(RxData[4]), .S(n192), .Q(n1749) );
  MUX21X1 U187 ( .IN1(n612), .IN2(RxData[5]), .S(n192), .Q(n1748) );
  MUX21X1 U188 ( .IN1(n611), .IN2(RxData[6]), .S(n192), .Q(n1747) );
  MUX21X1 U189 ( .IN1(n610), .IN2(RxData[7]), .S(n192), .Q(n1746) );
  AND2X1 U190 ( .IN1(n193), .IN2(n194), .Q(n192) );
  OAI22X1 U191 ( .IN1(n159), .IN2(n985), .IN3(n157), .IN4(n987), .QN(n194) );
  MUX21X1 U192 ( .IN1(n548), .IN2(n549), .S(RxStartFrm), .Q(n193) );
  MUX21X1 U193 ( .IN1(n633), .IN2(RxData[0]), .S(n195), .Q(n1745) );
  MUX21X1 U194 ( .IN1(n632), .IN2(RxData[7]), .S(n195), .Q(n1744) );
  MUX21X1 U195 ( .IN1(n631), .IN2(RxData[6]), .S(n195), .Q(n1743) );
  MUX21X1 U196 ( .IN1(n630), .IN2(RxData[5]), .S(n195), .Q(n1742) );
  MUX21X1 U197 ( .IN1(n629), .IN2(RxData[4]), .S(n195), .Q(n1741) );
  MUX21X1 U198 ( .IN1(n628), .IN2(RxData[3]), .S(n195), .Q(n1740) );
  MUX21X1 U199 ( .IN1(n627), .IN2(RxData[2]), .S(n195), .Q(n1739) );
  MUX21X1 U200 ( .IN1(n626), .IN2(RxData[1]), .S(n195), .Q(n1738) );
  AOI221X1 U201 ( .IN1(n548), .IN2(n157), .IN3(n549), .IN4(n159), .IN5(n160), 
        .QN(n195) );
  AO21X1 U202 ( .IN1(n157), .IN2(n159), .IN3(n196), .Q(n160) );
  INVX0 U203 ( .INP(n197), .ZN(n196) );
  MUX21X1 U204 ( .IN1(n985), .IN2(n987), .S(RxStartFrm), .Q(n197) );
  NAND2X0 U205 ( .IN1(n198), .IN2(n640), .QN(n159) );
  NAND2X0 U206 ( .IN1(n199), .IN2(n552), .QN(n157) );
  AO21X1 U207 ( .IN1(n549), .IN2(n200), .IN3(n201), .Q(n1737) );
  MUX21X1 U208 ( .IN1(n202), .IN2(n198), .S(n9), .Q(n201) );
  NOR2X0 U209 ( .IN1(n198), .IN2(n200), .QN(n202) );
  AO21X1 U210 ( .IN1(n200), .IN2(n158), .IN3(n203), .Q(n1736) );
  MUX21X1 U211 ( .IN1(n204), .IN2(n205), .S(n547), .Q(n203) );
  NOR2X0 U212 ( .IN1(n9), .IN2(n206), .QN(n205) );
  MUX21X1 U213 ( .IN1(n207), .IN2(n9), .S(n198), .Q(n204) );
  INVX0 U214 ( .INP(n206), .ZN(n198) );
  NAND4X0 U215 ( .IN1(n552), .IN2(RxValid), .IN3(n101), .IN4(n685), .QN(n206)
         );
  INVX0 U216 ( .INP(RxStartFrm), .ZN(n101) );
  XOR2X1 U217 ( .IN1(n987), .IN2(n549), .Q(n158) );
  AO22X1 U218 ( .IN1(n161), .IN2(RxDataLatched2[0]), .IN3(n208), .IN4(
        RxData[0]), .Q(n1735) );
  AO22X1 U219 ( .IN1(n161), .IN2(RxDataLatched2[1]), .IN3(n208), .IN4(
        RxData[1]), .Q(n1734) );
  AO22X1 U220 ( .IN1(n161), .IN2(RxDataLatched2[2]), .IN3(n208), .IN4(
        RxData[2]), .Q(n1733) );
  AO22X1 U221 ( .IN1(n161), .IN2(RxDataLatched2[3]), .IN3(n208), .IN4(
        RxData[3]), .Q(n1732) );
  AO22X1 U222 ( .IN1(n161), .IN2(RxDataLatched2[4]), .IN3(n208), .IN4(
        RxData[4]), .Q(n1731) );
  AO22X1 U223 ( .IN1(n161), .IN2(RxDataLatched2[5]), .IN3(n208), .IN4(
        RxData[5]), .Q(n1730) );
  AO22X1 U224 ( .IN1(n161), .IN2(RxDataLatched2[6]), .IN3(n208), .IN4(
        RxData[6]), .Q(n1729) );
  AO22X1 U225 ( .IN1(n161), .IN2(RxDataLatched2[7]), .IN3(n208), .IN4(
        RxData[7]), .Q(n1728) );
  INVX0 U226 ( .INP(n209), .ZN(n208) );
  AO22X1 U227 ( .IN1(n161), .IN2(RxDataLatched2[8]), .IN3(n210), .IN4(n617), 
        .Q(n1727) );
  AO22X1 U228 ( .IN1(n161), .IN2(RxDataLatched2[9]), .IN3(n210), .IN4(n616), 
        .Q(n1726) );
  AO22X1 U229 ( .IN1(n161), .IN2(RxDataLatched2[10]), .IN3(n210), .IN4(n615), 
        .Q(n1725) );
  AO22X1 U230 ( .IN1(n161), .IN2(RxDataLatched2[11]), .IN3(n210), .IN4(n614), 
        .Q(n1724) );
  AO22X1 U231 ( .IN1(n161), .IN2(RxDataLatched2[12]), .IN3(n210), .IN4(n613), 
        .Q(n1723) );
  AO22X1 U232 ( .IN1(n161), .IN2(RxDataLatched2[13]), .IN3(n210), .IN4(n612), 
        .Q(n1722) );
  AO22X1 U233 ( .IN1(n161), .IN2(RxDataLatched2[14]), .IN3(n210), .IN4(n611), 
        .Q(n1721) );
  AO22X1 U234 ( .IN1(n161), .IN2(RxDataLatched2[15]), .IN3(n210), .IN4(n610), 
        .Q(n1720) );
  NAND2X0 U235 ( .IN1(n209), .IN2(n211), .QN(n210) );
  OR3X1 U236 ( .IN1(n9), .IN2(n547), .IN3(n161), .Q(n211) );
  NAND2X0 U237 ( .IN1(n177), .IN2(n212), .QN(n209) );
  AO21X1 U238 ( .IN1(n547), .IN2(n9), .IN3(n652), .Q(n212) );
  AO22X1 U239 ( .IN1(n161), .IN2(RxDataLatched2[16]), .IN3(n213), .IN4(n633), 
        .Q(n1719) );
  AO22X1 U240 ( .IN1(n161), .IN2(RxDataLatched2[17]), .IN3(n213), .IN4(n626), 
        .Q(n1718) );
  AO22X1 U241 ( .IN1(n161), .IN2(RxDataLatched2[18]), .IN3(n213), .IN4(n627), 
        .Q(n1717) );
  AO22X1 U242 ( .IN1(n161), .IN2(RxDataLatched2[19]), .IN3(n213), .IN4(n628), 
        .Q(n1716) );
  AO22X1 U243 ( .IN1(n161), .IN2(RxDataLatched2[20]), .IN3(n213), .IN4(n629), 
        .Q(n1715) );
  AO22X1 U244 ( .IN1(n161), .IN2(RxDataLatched2[21]), .IN3(n213), .IN4(n630), 
        .Q(n1714) );
  AO22X1 U245 ( .IN1(n161), .IN2(RxDataLatched2[22]), .IN3(n213), .IN4(n631), 
        .Q(n1713) );
  AO22X1 U246 ( .IN1(n161), .IN2(RxDataLatched2[23]), .IN3(n213), .IN4(n632), 
        .Q(n1712) );
  AND2X1 U247 ( .IN1(n214), .IN2(n177), .Q(n213) );
  NAND3X0 U248 ( .IN1(n700), .IN2(n636), .IN3(n547), .QN(n214) );
  INVX0 U249 ( .INP(n177), .ZN(n161) );
  AO22X1 U250 ( .IN1(n189), .IN2(n215), .IN3(n216), .IN4(n199), .Q(n177) );
  INVX0 U251 ( .INP(n184), .ZN(n199) );
  NAND2X0 U252 ( .IN1(n200), .IN2(n640), .QN(n184) );
  NOR2X0 U253 ( .IN1(n549), .IN2(n987), .QN(n216) );
  OAI22X1 U254 ( .IN1(n552), .IN2(n652), .IN3(n187), .IN4(RxStartFrm), .QN(
        n215) );
  NAND3X0 U255 ( .IN1(n640), .IN2(n685), .IN3(RxValid), .QN(n187) );
  NOR2X0 U256 ( .IN1(n985), .IN2(n548), .QN(n189) );
  AO22X1 U257 ( .IN1(n217), .IN2(n218), .IN3(rx_burst_en), .IN4(n219), .Q(
        n1711) );
  AO21X1 U258 ( .IN1(n220), .IN2(n221), .IN3(n222), .Q(n219) );
  NAND3X0 U259 ( .IN1(rx_burst_cnt[1]), .IN2(n1), .IN3(rx_burst_cnt[0]), .QN(
        n221) );
  OR3X1 U260 ( .IN1(rxfifo_cnt[4]), .IN2(rxfifo_cnt[3]), .IN3(n223), .Q(n217)
         );
  OA21X1 U261 ( .IN1(n551), .IN2(n224), .IN3(rxfifo_cnt[2]), .Q(n223) );
  OR2X1 U262 ( .IN1(rxfifo_cnt[1]), .IN2(rxfifo_cnt[0]), .Q(n224) );
  NAND2X0 U263 ( .IN1(n225), .IN2(n226), .QN(n1710) );
  NAND3X0 U264 ( .IN1(n164), .IN2(n727), .IN3(n165), .QN(n226) );
  OA22X1 U265 ( .IN1(n995), .IN2(TxDone_wb), .IN3(n753), .IN4(n651), .Q(n1709)
         );
  MUX21X1 U266 ( .IN1(n227), .IN2(n650), .S(n228), .Q(n1708) );
  OA21X1 U267 ( .IN1(n996), .IN2(TxRetry_wb), .IN3(n14), .Q(n228) );
  OR2X1 U268 ( .IN1(TxRetry_wb), .IN2(n996), .Q(n227) );
  OA21X1 U269 ( .IN1(N848), .IN2(n726), .IN3(n140), .Q(n1707) );
  NAND2X0 U270 ( .IN1(n229), .IN2(n230), .QN(n1706) );
  NAND4X0 U271 ( .IN1(n222), .IN2(n231), .IN3(n232), .IN4(n728), .QN(n230) );
  AO22X1 U272 ( .IN1(n233), .IN2(n126), .IN3(tx_burst_cnt[0]), .IN4(n127), .Q(
        n1705) );
  AO22X1 U273 ( .IN1(n126), .IN2(n234), .IN3(tx_burst_cnt[1]), .IN4(n127), .Q(
        n1704) );
  AND2X1 U274 ( .IN1(n130), .IN2(n235), .Q(n127) );
  OA21X1 U275 ( .IN1(n236), .IN2(n237), .IN3(n229), .Q(n130) );
  AO22X1 U276 ( .IN1(n233), .IN2(n238), .IN3(n222), .IN4(rx_burst_cnt[0]), .Q(
        n1703) );
  AO22X1 U277 ( .IN1(n222), .IN2(rx_burst_cnt[1]), .IN3(n238), .IN4(n234), .Q(
        n1702) );
  XOR2X1 U278 ( .IN1(n233), .IN2(n239), .Q(n234) );
  AO22X1 U279 ( .IN1(n125), .IN2(n238), .IN3(n222), .IN4(rx_burst_cnt[2]), .Q(
        n1701) );
  NOR2X0 U280 ( .IN1(n218), .IN2(n238), .QN(n222) );
  XOR2X1 U281 ( .IN1(n240), .IN2(n241), .Q(n125) );
  OR2X1 U282 ( .IN1(n233), .IN2(n239), .Q(n240) );
  AO21X1 U283 ( .IN1(n165), .IN2(m_wb_we_o), .IN3(n242), .Q(n1700) );
  AO21X1 U284 ( .IN1(n220), .IN2(m_wb_cyc_o), .IN3(n243), .Q(n1699) );
  NAND2X0 U285 ( .IN1(n705), .IN2(n165), .QN(n1698) );
  AO221X1 U286 ( .IN1(n165), .IN2(m_wb_sel_o[1]), .IN3(n549), .IN4(n242), 
        .IN5(n244), .Q(n1697) );
  AO21X1 U287 ( .IN1(n165), .IN2(m_wb_sel_o[2]), .IN3(n244), .Q(n1696) );
  AO21X1 U288 ( .IN1(n987), .IN2(n242), .IN3(n245), .Q(n244) );
  AO221X1 U289 ( .IN1(n246), .IN2(n549), .IN3(n165), .IN4(m_wb_sel_o[3]), 
        .IN5(n245), .Q(n1695) );
  NOR2X0 U290 ( .IN1(n162), .IN2(n704), .QN(n246) );
  NAND2X0 U291 ( .IN1(n225), .IN2(n247), .QN(n1694) );
  NAND3X0 U292 ( .IN1(n165), .IN2(n634), .IN3(n220), .QN(n247) );
  INVX0 U293 ( .INP(n218), .ZN(n220) );
  NAND2X0 U294 ( .IN1(n164), .IN2(n229), .QN(n218) );
  NAND4X0 U295 ( .IN1(n248), .IN2(n249), .IN3(n250), .IN4(n251), .QN(n229) );
  OR2X1 U296 ( .IN1(n117), .IN2(n252), .Q(n250) );
  MUX21X1 U297 ( .IN1(n253), .IN2(n254), .S(n237), .Q(n248) );
  NAND2X0 U298 ( .IN1(tx_burst_en), .IN2(n727), .QN(n254) );
  NAND3X0 U299 ( .IN1(n255), .IN2(n256), .IN3(RxBufferEmpty), .QN(n164) );
  INVX0 U300 ( .INP(n237), .ZN(n256) );
  AO21X1 U301 ( .IN1(n252), .IN2(n251), .IN3(n257), .Q(n255) );
  OA21X1 U302 ( .IN1(n553), .IN2(n634), .IN3(n258), .Q(n1693) );
  AO22X1 U303 ( .IN1(n95), .IN2(n732), .IN3(n259), .IN4(r_RxEn), .Q(n1692) );
  NOR2X0 U304 ( .IN1(n142), .IN2(n640), .QN(n259) );
  AO22X1 U305 ( .IN1(n644), .IN2(n260), .IN3(BDCs[0]), .IN4(n261), .Q(n1691)
         );
  AO22X1 U306 ( .IN1(n643), .IN2(n260), .IN3(BDCs[1]), .IN4(n261), .Q(n1690)
         );
  AO22X1 U307 ( .IN1(n642), .IN2(n260), .IN3(BDCs[2]), .IN4(n261), .Q(n1689)
         );
  AO22X1 U308 ( .IN1(n641), .IN2(n260), .IN3(BDCs[3]), .IN4(n261), .Q(n1688)
         );
  AND2X1 U309 ( .IN1(WB_WE_I), .IN2(n107), .Q(n261) );
  MUX21X1 U310 ( .IN1(n608), .IN2(n262), .S(n107), .Q(n1687) );
  NOR2X0 U311 ( .IN1(WB_WE_I), .IN2(n263), .QN(n262) );
  NOR4X0 U312 ( .IN1(BDCs[3]), .IN2(BDCs[2]), .IN3(BDCs[1]), .IN4(BDCs[0]), 
        .QN(n263) );
  NAND2X0 U313 ( .IN1(n260), .IN2(n264), .QN(n1686) );
  NAND3X0 U314 ( .IN1(n265), .IN2(WbEn), .IN3(n106), .QN(n264) );
  NOR2X0 U315 ( .IN1(n722), .IN2(n266), .QN(n1685) );
  INVX0 U316 ( .INP(n267), .ZN(n266) );
  MUX21X1 U317 ( .IN1(n637), .IN2(WB_DAT_O[15]), .S(n97), .Q(n267) );
  AO22X1 U318 ( .IN1(n687), .IN2(n609), .IN3(n1465), .IN4(ShiftEndedSync1), 
        .Q(n1684) );
  AO221X1 U319 ( .IN1(ram_di[0]), .IN2(n106), .IN3(WB_DAT_I[0]), .IN4(n107), 
        .IN5(n268), .Q(n1683) );
  AO22X1 U320 ( .IN1(CarrierSenseLost), .IN2(n109), .IN3(n658), .IN4(n110), 
        .Q(n268) );
  AO221X1 U321 ( .IN1(ram_di[1]), .IN2(n106), .IN3(WB_DAT_I[1]), .IN4(n107), 
        .IN5(n269), .Q(n1682) );
  AO22X1 U322 ( .IN1(DeferLatched), .IN2(n109), .IN3(n659), .IN4(n110), .Q(
        n269) );
  AO221X1 U323 ( .IN1(ram_di[2]), .IN2(n106), .IN3(WB_DAT_I[2]), .IN4(n107), 
        .IN5(n270), .Q(n1681) );
  AO22X1 U324 ( .IN1(LateCollLatched), .IN2(n109), .IN3(n660), .IN4(n110), .Q(
        n270) );
  AO221X1 U325 ( .IN1(ram_di[3]), .IN2(n106), .IN3(WB_DAT_I[3]), .IN4(n107), 
        .IN5(n271), .Q(n1680) );
  AO22X1 U326 ( .IN1(RetryLimit), .IN2(n109), .IN3(n661), .IN4(n110), .Q(n271)
         );
  AO221X1 U327 ( .IN1(ram_di[4]), .IN2(n106), .IN3(WB_DAT_I[4]), .IN4(n107), 
        .IN5(n272), .Q(n1679) );
  AO22X1 U328 ( .IN1(RetryCntLatched[0]), .IN2(n109), .IN3(n662), .IN4(n110), 
        .Q(n272) );
  AO221X1 U329 ( .IN1(ram_di[5]), .IN2(n106), .IN3(WB_DAT_I[5]), .IN4(n107), 
        .IN5(n273), .Q(n1678) );
  AO22X1 U330 ( .IN1(RetryCntLatched[1]), .IN2(n109), .IN3(n663), .IN4(n110), 
        .Q(n273) );
  AO221X1 U331 ( .IN1(ram_di[6]), .IN2(n106), .IN3(WB_DAT_I[6]), .IN4(n107), 
        .IN5(n274), .Q(n1677) );
  AO22X1 U332 ( .IN1(RetryCntLatched[2]), .IN2(n109), .IN3(n656), .IN4(n110), 
        .Q(n274) );
  AO221X1 U333 ( .IN1(ram_di[7]), .IN2(n106), .IN3(WB_DAT_I[7]), .IN4(n107), 
        .IN5(n275), .Q(n1676) );
  AO22X1 U334 ( .IN1(RetryCntLatched[3]), .IN2(n109), .IN3(n664), .IN4(n110), 
        .Q(n275) );
  AO221X1 U335 ( .IN1(ram_di[8]), .IN2(n106), .IN3(WB_DAT_I[8]), .IN4(n107), 
        .IN5(n276), .Q(n1675) );
  AO22X1 U336 ( .IN1(n109), .IN2(TxUnderRun), .IN3(n665), .IN4(n110), .Q(n276)
         );
  AO22X1 U337 ( .IN1(WB_DAT_I[9]), .IN2(n107), .IN3(ram_di[9]), .IN4(n106), 
        .Q(n1674) );
  AO22X1 U338 ( .IN1(WB_DAT_I[10]), .IN2(n107), .IN3(ram_di[10]), .IN4(n106), 
        .Q(n1673) );
  AO222X1 U339 ( .IN1(WB_DAT_I[11]), .IN2(n107), .IN3(ram_di[11]), .IN4(n106), 
        .IN5(n109), .IN6(PerPacketCrcEn), .Q(n1672) );
  AO222X1 U340 ( .IN1(WB_DAT_I[12]), .IN2(n107), .IN3(ram_di[12]), .IN4(n106), 
        .IN5(n109), .IN6(PerPacketPad), .Q(n1671) );
  AO221X1 U341 ( .IN1(ram_di[13]), .IN2(n106), .IN3(WB_DAT_I[13]), .IN4(n107), 
        .IN5(n277), .Q(n1670) );
  AO22X1 U342 ( .IN1(n647), .IN2(n109), .IN3(n638), .IN4(n110), .Q(n277) );
  AO221X1 U343 ( .IN1(ram_di[14]), .IN2(n106), .IN3(WB_DAT_I[14]), .IN4(n107), 
        .IN5(n278), .Q(n1669) );
  AO22X1 U344 ( .IN1(n646), .IN2(n109), .IN3(n110), .IN4(n639), .Q(n278) );
  AO22X1 U345 ( .IN1(WB_DAT_I[15]), .IN2(n107), .IN3(ram_di[15]), .IN4(n106), 
        .Q(n1668) );
  AO221X1 U346 ( .IN1(ram_di[16]), .IN2(n106), .IN3(WB_DAT_I[16]), .IN4(n107), 
        .IN5(n279), .Q(n1667) );
  AO22X1 U347 ( .IN1(n592), .IN2(n109), .IN3(n666), .IN4(n110), .Q(n279) );
  AO221X1 U348 ( .IN1(ram_di[17]), .IN2(n106), .IN3(WB_DAT_I[17]), .IN4(n107), 
        .IN5(n280), .Q(n1666) );
  AO22X1 U349 ( .IN1(n593), .IN2(n109), .IN3(n667), .IN4(n110), .Q(n280) );
  AO221X1 U350 ( .IN1(ram_di[18]), .IN2(n106), .IN3(WB_DAT_I[18]), .IN4(n107), 
        .IN5(n281), .Q(n1665) );
  AO22X1 U351 ( .IN1(n594), .IN2(n109), .IN3(n668), .IN4(n110), .Q(n281) );
  AO221X1 U352 ( .IN1(ram_di[19]), .IN2(n106), .IN3(WB_DAT_I[19]), .IN4(n107), 
        .IN5(n282), .Q(n1664) );
  AO22X1 U353 ( .IN1(n595), .IN2(n109), .IN3(n669), .IN4(n110), .Q(n282) );
  AO221X1 U354 ( .IN1(ram_di[20]), .IN2(n106), .IN3(WB_DAT_I[20]), .IN4(n107), 
        .IN5(n283), .Q(n1663) );
  AO22X1 U355 ( .IN1(n596), .IN2(n109), .IN3(n670), .IN4(n110), .Q(n283) );
  AO221X1 U356 ( .IN1(ram_di[21]), .IN2(n106), .IN3(WB_DAT_I[21]), .IN4(n107), 
        .IN5(n284), .Q(n1662) );
  AO22X1 U357 ( .IN1(n597), .IN2(n109), .IN3(n671), .IN4(n110), .Q(n284) );
  AO221X1 U358 ( .IN1(ram_di[22]), .IN2(n106), .IN3(WB_DAT_I[22]), .IN4(n107), 
        .IN5(n285), .Q(n1661) );
  AO22X1 U359 ( .IN1(n598), .IN2(n109), .IN3(n672), .IN4(n110), .Q(n285) );
  AO221X1 U360 ( .IN1(ram_di[23]), .IN2(n106), .IN3(WB_DAT_I[23]), .IN4(n107), 
        .IN5(n286), .Q(n1660) );
  AO22X1 U361 ( .IN1(n599), .IN2(n109), .IN3(n673), .IN4(n110), .Q(n286) );
  AO221X1 U362 ( .IN1(ram_di[24]), .IN2(n106), .IN3(WB_DAT_I[24]), .IN4(n107), 
        .IN5(n287), .Q(n1659) );
  AO22X1 U363 ( .IN1(n600), .IN2(n109), .IN3(n675), .IN4(n110), .Q(n287) );
  AO221X1 U364 ( .IN1(ram_di[25]), .IN2(n106), .IN3(WB_DAT_I[25]), .IN4(n107), 
        .IN5(n288), .Q(n1658) );
  AO22X1 U365 ( .IN1(n601), .IN2(n109), .IN3(n677), .IN4(n110), .Q(n288) );
  AO221X1 U366 ( .IN1(ram_di[26]), .IN2(n106), .IN3(WB_DAT_I[26]), .IN4(n107), 
        .IN5(n289), .Q(n1657) );
  AO22X1 U367 ( .IN1(n602), .IN2(n109), .IN3(n678), .IN4(n110), .Q(n289) );
  AO221X1 U368 ( .IN1(ram_di[27]), .IN2(n106), .IN3(WB_DAT_I[27]), .IN4(n107), 
        .IN5(n290), .Q(n1656) );
  AO22X1 U369 ( .IN1(n603), .IN2(n109), .IN3(n680), .IN4(n110), .Q(n290) );
  AO221X1 U370 ( .IN1(ram_di[28]), .IN2(n106), .IN3(WB_DAT_I[28]), .IN4(n107), 
        .IN5(n291), .Q(n1655) );
  AO22X1 U371 ( .IN1(n604), .IN2(n109), .IN3(n681), .IN4(n110), .Q(n291) );
  AO221X1 U372 ( .IN1(ram_di[29]), .IN2(n106), .IN3(WB_DAT_I[29]), .IN4(n107), 
        .IN5(n292), .Q(n1654) );
  AO22X1 U373 ( .IN1(n605), .IN2(n109), .IN3(n682), .IN4(n110), .Q(n292) );
  AO221X1 U374 ( .IN1(ram_di[30]), .IN2(n106), .IN3(WB_DAT_I[30]), .IN4(n107), 
        .IN5(n293), .Q(n1653) );
  AO22X1 U375 ( .IN1(n606), .IN2(n109), .IN3(n683), .IN4(n110), .Q(n293) );
  MUX21X1 U376 ( .IN1(n294), .IN2(n295), .S(n111), .Q(n1652) );
  OA21X1 U377 ( .IN1(n296), .IN2(n297), .IN3(WB_DAT_O[15]), .Q(n295) );
  NAND4X0 U378 ( .IN1(n298), .IN2(n299), .IN3(n300), .IN4(n301), .QN(n297) );
  NOR4X0 U379 ( .IN1(WB_DAT_O[24]), .IN2(WB_DAT_O[23]), .IN3(WB_DAT_O[22]), 
        .IN4(WB_DAT_O[21]), .QN(n301) );
  OAI21X1 U380 ( .IN1(WB_DAT_O[17]), .IN2(WB_DAT_O[16]), .IN3(WB_DAT_O[18]), 
        .QN(n300) );
  INVX0 U381 ( .INP(WB_DAT_O[20]), .ZN(n299) );
  INVX0 U382 ( .INP(WB_DAT_O[19]), .ZN(n298) );
  OR4X1 U383 ( .IN1(WB_DAT_O[26]), .IN2(WB_DAT_O[27]), .IN3(WB_DAT_O[25]), 
        .IN4(n302), .Q(n296) );
  OR4X1 U384 ( .IN1(WB_DAT_O[31]), .IN2(WB_DAT_O[30]), .IN3(WB_DAT_O[29]), 
        .IN4(WB_DAT_O[28]), .Q(n302) );
  NOR2X0 U385 ( .IN1(n746), .IN2(n303), .QN(n294) );
  MUX21X1 U386 ( .IN1(N857), .IN2(n138), .S(n735), .Q(n1651) );
  INVX0 U387 ( .INP(n304), .ZN(n138) );
  MUX21X1 U388 ( .IN1(n305), .IN2(WB_DAT_O[0]), .S(n306), .Q(n1650) );
  NOR2X0 U389 ( .IN1(n840), .IN2(n767), .QN(n305) );
  MUX21X1 U390 ( .IN1(n307), .IN2(WB_DAT_O[1]), .S(n306), .Q(n1649) );
  NOR2X0 U391 ( .IN1(n989), .IN2(n767), .QN(n307) );
  AO222X1 U392 ( .IN1(n113), .IN2(n308), .IN3(n309), .IN4(n35), .IN5(
        WB_DAT_O[16]), .IN6(n111), .Q(n1648) );
  AO21X1 U393 ( .IN1(n113), .IN2(n840), .IN3(n310), .Q(n309) );
  AO222X1 U394 ( .IN1(n310), .IN2(n38), .IN3(n311), .IN4(n113), .IN5(
        WB_DAT_O[17]), .IN6(n111), .Q(n1647) );
  XOR3X1 U395 ( .IN1(n721), .IN2(n308), .IN3(n312), .Q(n311) );
  AO222X1 U396 ( .IN1(n310), .IN2(n33), .IN3(n313), .IN4(n113), .IN5(
        WB_DAT_O[18]), .IN6(n111), .Q(n1646) );
  XOR3X1 U397 ( .IN1(n33), .IN2(n314), .IN3(n315), .Q(n313) );
  AO21X1 U398 ( .IN1(WB_DAT_O[19]), .IN2(n111), .IN3(n316), .Q(n1645) );
  MUX21X1 U399 ( .IN1(n317), .IN2(n318), .S(n708), .Q(n316) );
  NOR2X0 U400 ( .IN1(n319), .IN2(n320), .QN(n318) );
  AO222X1 U401 ( .IN1(n113), .IN2(n321), .IN3(n322), .IN4(n30), .IN5(
        WB_DAT_O[20]), .IN6(n111), .Q(n1644) );
  AO21X1 U402 ( .IN1(n113), .IN2(n11), .IN3(n317), .Q(n322) );
  AO21X1 U403 ( .IN1(n113), .IN2(n319), .IN3(n310), .Q(n317) );
  AO21X1 U404 ( .IN1(WB_DAT_O[21]), .IN2(n111), .IN3(n323), .Q(n1643) );
  MUX21X1 U405 ( .IN1(n324), .IN2(n325), .S(n710), .Q(n323) );
  NOR2X0 U406 ( .IN1(n326), .IN2(n320), .QN(n325) );
  AO222X1 U407 ( .IN1(n113), .IN2(n327), .IN3(n328), .IN4(n50), .IN5(
        WB_DAT_O[22]), .IN6(n111), .Q(n1642) );
  AO21X1 U408 ( .IN1(n113), .IN2(n29), .IN3(n324), .Q(n328) );
  AO21X1 U409 ( .IN1(n113), .IN2(n326), .IN3(n310), .Q(n324) );
  INVX0 U410 ( .INP(n321), .ZN(n326) );
  AO21X1 U411 ( .IN1(WB_DAT_O[23]), .IN2(n111), .IN3(n329), .Q(n1641) );
  MUX21X1 U412 ( .IN1(n330), .IN2(n331), .S(n712), .Q(n329) );
  NOR2X0 U413 ( .IN1(n332), .IN2(n320), .QN(n331) );
  AO222X1 U414 ( .IN1(n113), .IN2(n333), .IN3(n334), .IN4(n37), .IN5(
        WB_DAT_O[24]), .IN6(n111), .Q(n1640) );
  AO21X1 U415 ( .IN1(n113), .IN2(n12), .IN3(n330), .Q(n334) );
  AO21X1 U416 ( .IN1(n113), .IN2(n332), .IN3(n310), .Q(n330) );
  AO21X1 U417 ( .IN1(WB_DAT_O[25]), .IN2(n111), .IN3(n335), .Q(n1639) );
  MUX21X1 U418 ( .IN1(n336), .IN2(n337), .S(n714), .Q(n335) );
  NOR2X0 U419 ( .IN1(n338), .IN2(n320), .QN(n337) );
  AO221X1 U420 ( .IN1(n339), .IN2(n36), .IN3(WB_DAT_O[26]), .IN4(n111), .IN5(
        n340), .Q(n1638) );
  AO21X1 U421 ( .IN1(n113), .IN2(n3), .IN3(n336), .Q(n339) );
  AO21X1 U422 ( .IN1(n113), .IN2(n338), .IN3(n310), .Q(n336) );
  AO21X1 U423 ( .IN1(WB_DAT_O[27]), .IN2(n111), .IN3(n341), .Q(n1637) );
  MUX21X1 U424 ( .IN1(n342), .IN2(n340), .S(n716), .Q(n341) );
  AO221X1 U425 ( .IN1(n343), .IN2(n19), .IN3(WB_DAT_O[28]), .IN4(n111), .IN5(
        n344), .Q(n1636) );
  AO21X1 U426 ( .IN1(n113), .IN2(n4), .IN3(n342), .Q(n343) );
  AO21X1 U427 ( .IN1(WB_DAT_O[29]), .IN2(n111), .IN3(n345), .Q(n1635) );
  MUX21X1 U428 ( .IN1(n346), .IN2(n344), .S(n718), .Q(n345) );
  AO21X1 U429 ( .IN1(WB_DAT_O[30]), .IN2(n111), .IN3(n347), .Q(n1634) );
  MUX21X1 U430 ( .IN1(n114), .IN2(n348), .S(n719), .Q(n347) );
  AND2X1 U431 ( .IN1(n718), .IN2(n344), .Q(n348) );
  NOR2X0 U432 ( .IN1(n349), .IN2(n350), .QN(n344) );
  INVX0 U433 ( .INP(n340), .ZN(n349) );
  NOR2X0 U434 ( .IN1(n351), .IN2(n320), .QN(n340) );
  AO21X1 U435 ( .IN1(n113), .IN2(n43), .IN3(n346), .Q(n114) );
  AO21X1 U436 ( .IN1(n113), .IN2(n350), .IN3(n342), .Q(n346) );
  AO21X1 U437 ( .IN1(n113), .IN2(n351), .IN3(n310), .Q(n342) );
  NOR2X0 U438 ( .IN1(n767), .IN2(n111), .QN(n310) );
  NAND3X0 U439 ( .IN1(n715), .IN2(n714), .IN3(n333), .QN(n351) );
  INVX0 U440 ( .INP(n338), .ZN(n333) );
  NAND3X0 U441 ( .IN1(n713), .IN2(n712), .IN3(n327), .QN(n338) );
  INVX0 U442 ( .INP(n332), .ZN(n327) );
  NAND3X0 U443 ( .IN1(n711), .IN2(n710), .IN3(n321), .QN(n332) );
  NOR3X0 U444 ( .IN1(n30), .IN2(n11), .IN3(n319), .QN(n321) );
  AO21X1 U445 ( .IN1(n315), .IN2(n314), .IN3(n33), .Q(n319) );
  AO22X1 U446 ( .IN1(n352), .IN2(n312), .IN3(n353), .IN4(n38), .Q(n315) );
  NAND2X0 U447 ( .IN1(n354), .IN2(n308), .QN(n353) );
  INVX0 U448 ( .INP(n354), .ZN(n312) );
  OA21X1 U449 ( .IN1(n989), .IN2(n840), .IN3(n314), .Q(n354) );
  NAND2X0 U450 ( .IN1(n989), .IN2(n840), .QN(n314) );
  INVX0 U451 ( .INP(n308), .ZN(n352) );
  NOR2X0 U452 ( .IN1(n35), .IN2(n840), .QN(n308) );
  INVX0 U453 ( .INP(n320), .ZN(n113) );
  NAND3X0 U454 ( .IN1(n355), .IN2(n94), .IN3(n767), .QN(n320) );
  AND2X1 U455 ( .IN1(m_wb_ack_i), .IN2(n727), .Q(n767) );
  NOR3X0 U456 ( .IN1(n356), .IN2(n357), .IN3(n358), .QN(n1633) );
  AND2X1 U457 ( .IN1(n93), .IN2(n533), .Q(n358) );
  MUX21X1 U458 ( .IN1(n359), .IN2(n360), .S(n361), .Q(n1632) );
  NOR2X0 U459 ( .IN1(n720), .IN2(n355), .QN(n360) );
  NOR2X0 U460 ( .IN1(n990), .IN2(n303), .QN(n359) );
  MUX21X1 U461 ( .IN1(n362), .IN2(n363), .S(n361), .Q(n1631) );
  AND2X1 U462 ( .IN1(LatchValidBytes), .IN2(n1435), .Q(n361) );
  NOR2X0 U463 ( .IN1(n721), .IN2(n355), .QN(n363) );
  NOR2X0 U464 ( .IN1(n991), .IN2(n303), .QN(n362) );
  NOR2X0 U465 ( .IN1(n100), .IN2(n364), .QN(n1630) );
  MUX21X1 U466 ( .IN1(n686), .IN2(n365), .S(n1445), .Q(n364) );
  NAND3X0 U467 ( .IN1(n686), .IN2(n692), .IN3(n366), .QN(n365) );
  MUX41X1 U468 ( .IN1(n367), .IN3(n368), .IN2(n369), .IN4(n370), .S0(n991), 
        .S1(n990), .Q(n366) );
  NAND2X0 U469 ( .IN1(n536), .IN2(n371), .QN(n100) );
  INVX0 U470 ( .INP(TxAbort), .ZN(n371) );
  MUX21X1 U471 ( .IN1(n372), .IN2(n589), .S(n373), .Q(n1629) );
  NOR4X0 U472 ( .IN1(TxRetry), .IN2(TxAbort), .IN3(TxEndFrm), .IN4(n374), .QN(
        n373) );
  OA21X1 U473 ( .IN1(n375), .IN2(n749), .IN3(n692), .Q(n372) );
  NOR3X0 U474 ( .IN1(TxEndFrm), .IN2(TxRetry), .IN3(TxAbort), .QN(n375) );
  AO221X1 U475 ( .IN1(n376), .IN2(ReadTxDataFromFifo_tck), .IN3(n748), .IN4(
        n377), .IN5(n378), .Q(n1628) );
  NAND2X0 U476 ( .IN1(ReadTxDataFromFifo_syncb2), .IN2(n1448), .QN(n376) );
  AO22X1 U477 ( .IN1(n379), .IN2(n589), .IN3(n380), .IN4(TxBufferAlmostEmpty), 
        .Q(n1627) );
  NOR2X0 U478 ( .IN1(n381), .IN2(n382), .QN(n380) );
  INVX0 U479 ( .INP(n303), .ZN(n379) );
  AO22X1 U480 ( .IN1(n723), .IN2(TxStartFrm_wb), .IN3(n383), .IN4(n994), .Q(
        n1626) );
  OA21X1 U481 ( .IN1(n357), .IN2(TxBufferFull), .IN3(n733), .Q(n383) );
  INVX0 U482 ( .INP(n382), .ZN(n357) );
  NAND3X0 U483 ( .IN1(n721), .IN2(n720), .IN3(n119), .QN(n382) );
  INVX0 U484 ( .INP(n355), .ZN(n119) );
  NAND2X0 U485 ( .IN1(n1433), .IN2(n384), .QN(n1625) );
  AO221X1 U486 ( .IN1(n537), .IN2(TxAbort), .IN3(TxRetry), .IN4(n536), .IN5(
        n385), .Q(n384) );
  NAND2X0 U487 ( .IN1(TxStartFrm), .IN2(n724), .QN(n385) );
  AO21X1 U488 ( .IN1(n545), .IN2(n386), .IN3(n387), .Q(n1624) );
  MUX21X1 U489 ( .IN1(n388), .IN2(n389), .S(n544), .Q(n387) );
  NOR3X0 U490 ( .IN1(n390), .IN2(n386), .IN3(n389), .QN(n388) );
  NAND2X0 U491 ( .IN1(n391), .IN2(n392), .QN(n1623) );
  OAI21X1 U492 ( .IN1(n393), .IN2(n394), .IN3(n386), .QN(n392) );
  INVX0 U493 ( .INP(n395), .ZN(n386) );
  MUX21X1 U494 ( .IN1(n396), .IN2(n397), .S(n389), .Q(n391) );
  AND2X1 U495 ( .IN1(n398), .IN2(n98), .Q(n389) );
  NOR2X0 U496 ( .IN1(n369), .IN2(n367), .QN(n397) );
  NAND3X0 U497 ( .IN1(n395), .IN2(n694), .IN3(n398), .QN(n396) );
  NAND3X0 U498 ( .IN1(n381), .IN2(TxStartFrm), .IN3(n398), .QN(n395) );
  INVX0 U499 ( .INP(n390), .ZN(n398) );
  NAND2X0 U500 ( .IN1(n537), .IN2(n536), .QN(n390) );
  OAI21X1 U501 ( .IN1(n303), .IN2(n994), .IN3(n993), .QN(n1622) );
  AO21X1 U502 ( .IN1(n995), .IN2(TxDone_wb), .IN3(n356), .Q(n303) );
  AO21X1 U503 ( .IN1(n996), .IN2(TxRetry_wb), .IN3(n399), .Q(n356) );
  MUX21X1 U504 ( .IN1(TxData_wb[0]), .IN2(n588), .S(n400), .Q(n1621) );
  MUX21X1 U505 ( .IN1(TxData_wb[1]), .IN2(n587), .S(n400), .Q(n1620) );
  MUX21X1 U506 ( .IN1(TxData_wb[2]), .IN2(n586), .S(n400), .Q(n1619) );
  MUX21X1 U507 ( .IN1(TxData_wb[3]), .IN2(n585), .S(n400), .Q(n1618) );
  MUX21X1 U508 ( .IN1(TxData_wb[4]), .IN2(n584), .S(n400), .Q(n1617) );
  MUX21X1 U509 ( .IN1(TxData_wb[5]), .IN2(n583), .S(n400), .Q(n1616) );
  MUX21X1 U510 ( .IN1(TxData_wb[6]), .IN2(n582), .S(n400), .Q(n1615) );
  MUX21X1 U511 ( .IN1(TxData_wb[7]), .IN2(n581), .S(n400), .Q(n1614) );
  MUX21X1 U512 ( .IN1(TxData_wb[8]), .IN2(n580), .S(n400), .Q(n1613) );
  MUX21X1 U513 ( .IN1(TxData_wb[9]), .IN2(n579), .S(n400), .Q(n1612) );
  MUX21X1 U514 ( .IN1(TxData_wb[10]), .IN2(n578), .S(n400), .Q(n1611) );
  MUX21X1 U515 ( .IN1(TxData_wb[11]), .IN2(n577), .S(n400), .Q(n1610) );
  MUX21X1 U516 ( .IN1(TxData_wb[12]), .IN2(n576), .S(n400), .Q(n1609) );
  MUX21X1 U517 ( .IN1(TxData_wb[13]), .IN2(n575), .S(n400), .Q(n1608) );
  MUX21X1 U518 ( .IN1(TxData_wb[14]), .IN2(n574), .S(n400), .Q(n1607) );
  MUX21X1 U519 ( .IN1(TxData_wb[15]), .IN2(n573), .S(n400), .Q(n1606) );
  MUX21X1 U520 ( .IN1(TxData_wb[16]), .IN2(n572), .S(n400), .Q(n1605) );
  MUX21X1 U521 ( .IN1(TxData_wb[17]), .IN2(n571), .S(n400), .Q(n1604) );
  MUX21X1 U522 ( .IN1(TxData_wb[18]), .IN2(n570), .S(n400), .Q(n1603) );
  MUX21X1 U523 ( .IN1(TxData_wb[19]), .IN2(n569), .S(n400), .Q(n1602) );
  MUX21X1 U524 ( .IN1(TxData_wb[20]), .IN2(n568), .S(n400), .Q(n1601) );
  MUX21X1 U525 ( .IN1(TxData_wb[21]), .IN2(n567), .S(n400), .Q(n1600) );
  MUX21X1 U526 ( .IN1(TxData_wb[22]), .IN2(n566), .S(n400), .Q(n1599) );
  MUX21X1 U527 ( .IN1(TxData_wb[23]), .IN2(n565), .S(n400), .Q(n1598) );
  MUX21X1 U528 ( .IN1(TxData_wb[24]), .IN2(n564), .S(n400), .Q(n1597) );
  MUX21X1 U529 ( .IN1(TxData_wb[25]), .IN2(n563), .S(n400), .Q(n1596) );
  MUX21X1 U530 ( .IN1(TxData_wb[26]), .IN2(n562), .S(n400), .Q(n1595) );
  MUX21X1 U531 ( .IN1(TxData_wb[27]), .IN2(n561), .S(n400), .Q(n1594) );
  MUX21X1 U532 ( .IN1(TxData_wb[28]), .IN2(n560), .S(n400), .Q(n1593) );
  MUX21X1 U533 ( .IN1(TxData_wb[29]), .IN2(n559), .S(n400), .Q(n1592) );
  MUX21X1 U534 ( .IN1(TxData_wb[30]), .IN2(n558), .S(n400), .Q(n1591) );
  MUX21X1 U535 ( .IN1(TxData_wb[31]), .IN2(n557), .S(n400), .Q(n1590) );
  INVX0 U536 ( .INP(n374), .ZN(n377) );
  NAND2X0 U537 ( .IN1(n98), .IN2(n370), .QN(n374) );
  NAND2X0 U538 ( .IN1(n401), .IN2(n402), .QN(n378) );
  NAND3X0 U539 ( .IN1(n98), .IN2(TxStartFrm), .IN3(n368), .QN(n402) );
  AO221X1 U540 ( .IN1(TxData_wb[24]), .IN2(n403), .IN3(n404), .IN4(TxData[0]), 
        .IN5(n405), .Q(n1589) );
  AO22X1 U541 ( .IN1(n406), .IN2(n407), .IN3(n408), .IN4(n409), .Q(n405) );
  AO221X1 U542 ( .IN1(n588), .IN2(n370), .IN3(n368), .IN4(n564), .IN5(n410), 
        .Q(n409) );
  AO22X1 U543 ( .IN1(n367), .IN2(n580), .IN3(n369), .IN4(n572), .Q(n410) );
  AO222X1 U544 ( .IN1(n393), .IN2(TxData_wb[8]), .IN3(n394), .IN4(
        TxData_wb[16]), .IN5(n411), .IN6(TxData_wb[0]), .Q(n407) );
  AO221X1 U545 ( .IN1(TxData_wb[25]), .IN2(n403), .IN3(n404), .IN4(TxData[1]), 
        .IN5(n412), .Q(n1588) );
  AO22X1 U546 ( .IN1(n406), .IN2(n413), .IN3(n408), .IN4(n414), .Q(n412) );
  AO221X1 U547 ( .IN1(n369), .IN2(n571), .IN3(n367), .IN4(n579), .IN5(n415), 
        .Q(n414) );
  AO22X1 U548 ( .IN1(n563), .IN2(n368), .IN3(n587), .IN4(n370), .Q(n415) );
  AO222X1 U549 ( .IN1(n393), .IN2(TxData_wb[9]), .IN3(n394), .IN4(
        TxData_wb[17]), .IN5(n411), .IN6(TxData_wb[1]), .Q(n413) );
  AO221X1 U550 ( .IN1(TxData_wb[26]), .IN2(n403), .IN3(n404), .IN4(TxData[2]), 
        .IN5(n416), .Q(n1587) );
  AO22X1 U551 ( .IN1(n406), .IN2(n417), .IN3(n408), .IN4(n418), .Q(n416) );
  AO221X1 U552 ( .IN1(n369), .IN2(n570), .IN3(n367), .IN4(n578), .IN5(n419), 
        .Q(n418) );
  AO22X1 U553 ( .IN1(n562), .IN2(n368), .IN3(n586), .IN4(n370), .Q(n419) );
  AO222X1 U554 ( .IN1(n393), .IN2(TxData_wb[10]), .IN3(n394), .IN4(
        TxData_wb[18]), .IN5(n411), .IN6(TxData_wb[2]), .Q(n417) );
  AO221X1 U555 ( .IN1(TxData_wb[27]), .IN2(n403), .IN3(n404), .IN4(TxData[3]), 
        .IN5(n420), .Q(n1586) );
  AO22X1 U556 ( .IN1(n406), .IN2(n421), .IN3(n408), .IN4(n422), .Q(n420) );
  AO221X1 U557 ( .IN1(n369), .IN2(n569), .IN3(n367), .IN4(n577), .IN5(n423), 
        .Q(n422) );
  AO22X1 U558 ( .IN1(n561), .IN2(n368), .IN3(n585), .IN4(n370), .Q(n423) );
  AO222X1 U559 ( .IN1(n393), .IN2(TxData_wb[11]), .IN3(n394), .IN4(
        TxData_wb[19]), .IN5(n411), .IN6(TxData_wb[3]), .Q(n421) );
  AO221X1 U560 ( .IN1(TxData_wb[28]), .IN2(n403), .IN3(n404), .IN4(TxData[4]), 
        .IN5(n424), .Q(n1585) );
  AO22X1 U561 ( .IN1(n406), .IN2(n425), .IN3(n408), .IN4(n426), .Q(n424) );
  AO221X1 U562 ( .IN1(n369), .IN2(n568), .IN3(n367), .IN4(n576), .IN5(n427), 
        .Q(n426) );
  AO22X1 U563 ( .IN1(n560), .IN2(n368), .IN3(n584), .IN4(n370), .Q(n427) );
  AO222X1 U564 ( .IN1(n393), .IN2(TxData_wb[12]), .IN3(n394), .IN4(
        TxData_wb[20]), .IN5(n411), .IN6(TxData_wb[4]), .Q(n425) );
  AO221X1 U565 ( .IN1(TxData_wb[29]), .IN2(n403), .IN3(n404), .IN4(TxData[5]), 
        .IN5(n428), .Q(n1584) );
  AO22X1 U566 ( .IN1(n406), .IN2(n429), .IN3(n408), .IN4(n430), .Q(n428) );
  AO221X1 U567 ( .IN1(n369), .IN2(n567), .IN3(n367), .IN4(n575), .IN5(n431), 
        .Q(n430) );
  AO22X1 U568 ( .IN1(n559), .IN2(n368), .IN3(n583), .IN4(n370), .Q(n431) );
  AO222X1 U569 ( .IN1(n393), .IN2(TxData_wb[13]), .IN3(n394), .IN4(
        TxData_wb[21]), .IN5(n411), .IN6(TxData_wb[5]), .Q(n429) );
  AO221X1 U570 ( .IN1(TxData_wb[30]), .IN2(n403), .IN3(n404), .IN4(TxData[6]), 
        .IN5(n432), .Q(n1583) );
  AO22X1 U571 ( .IN1(n406), .IN2(n433), .IN3(n408), .IN4(n434), .Q(n432) );
  AO221X1 U572 ( .IN1(n369), .IN2(n566), .IN3(n367), .IN4(n574), .IN5(n435), 
        .Q(n434) );
  AO22X1 U573 ( .IN1(n558), .IN2(n368), .IN3(n582), .IN4(n370), .Q(n435) );
  AO222X1 U574 ( .IN1(n393), .IN2(TxData_wb[14]), .IN3(n394), .IN4(
        TxData_wb[22]), .IN5(n411), .IN6(TxData_wb[6]), .Q(n433) );
  AO221X1 U575 ( .IN1(TxData_wb[31]), .IN2(n403), .IN3(n404), .IN4(TxData[7]), 
        .IN5(n436), .Q(n1582) );
  AO22X1 U576 ( .IN1(n406), .IN2(n437), .IN3(n408), .IN4(n438), .Q(n436) );
  AO221X1 U577 ( .IN1(n369), .IN2(n565), .IN3(n367), .IN4(n573), .IN5(n439), 
        .Q(n438) );
  AO22X1 U578 ( .IN1(n557), .IN2(n368), .IN3(n581), .IN4(n370), .Q(n439) );
  NOR2X0 U579 ( .IN1(n544), .IN2(n543), .QN(n370) );
  NOR2X0 U580 ( .IN1(n694), .IN2(n693), .QN(n368) );
  NOR2X0 U581 ( .IN1(n693), .IN2(n543), .QN(n367) );
  NOR2X0 U582 ( .IN1(n694), .IN2(n544), .QN(n369) );
  INVX0 U583 ( .INP(n440), .ZN(n408) );
  AO222X1 U584 ( .IN1(n393), .IN2(TxData_wb[15]), .IN3(n394), .IN4(
        TxData_wb[23]), .IN5(n411), .IN6(TxData_wb[7]), .Q(n437) );
  NOR2X0 U585 ( .IN1(n688), .IN2(n545), .QN(n394) );
  NOR2X0 U586 ( .IN1(n689), .IN2(n546), .QN(n393) );
  AND3X1 U587 ( .IN1(n441), .IN2(n401), .IN3(n440), .Q(n404) );
  NAND3X0 U588 ( .IN1(n441), .IN2(n401), .IN3(n98), .QN(n440) );
  NOR2X0 U589 ( .IN1(n381), .IN2(n749), .QN(n98) );
  INVX0 U590 ( .INP(TxUsedData), .ZN(n381) );
  INVX0 U591 ( .INP(n406), .ZN(n401) );
  NAND2X0 U592 ( .IN1(n441), .IN2(n442), .QN(n403) );
  NAND3X0 U593 ( .IN1(n546), .IN2(n545), .IN3(n406), .QN(n442) );
  NOR2X0 U594 ( .IN1(TxStartFrm), .IN2(n1433), .QN(n406) );
  NAND3X0 U595 ( .IN1(TxUsedData), .IN2(TxStartFrm), .IN3(n411), .QN(n441) );
  NOR2X0 U596 ( .IN1(n546), .IN2(n545), .QN(n411) );
  OA21X1 U597 ( .IN1(n443), .IN2(n654), .IN3(n444), .Q(n1581) );
  INVX0 U598 ( .INP(n399), .ZN(n444) );
  NOR2X0 U599 ( .IN1(n696), .IN2(n1452), .QN(n399) );
  NOR2X0 U600 ( .IN1(n123), .IN2(n445), .QN(n443) );
  INVX0 U601 ( .INP(TxBufferEmpty), .ZN(n445) );
  OAI21X1 U602 ( .IN1(n746), .IN2(n542), .IN3(n140), .QN(n1580) );
  NAND3X0 U603 ( .IN1(n746), .IN2(n446), .IN3(n542), .QN(n140) );
  NAND2X0 U604 ( .IN1(n541), .IN2(n91), .QN(n446) );
  AO22X1 U605 ( .IN1(n447), .IN2(TxBDAddress[1]), .IN3(N800), .IN4(n448), .Q(
        n1579) );
  AO22X1 U606 ( .IN1(n447), .IN2(TxBDAddress[2]), .IN3(N801), .IN4(n448), .Q(
        n1578) );
  AO22X1 U607 ( .IN1(n447), .IN2(TxBDAddress[3]), .IN3(N802), .IN4(n448), .Q(
        n1577) );
  AO22X1 U608 ( .IN1(n447), .IN2(TxBDAddress[4]), .IN3(N803), .IN4(n448), .Q(
        n1576) );
  AO22X1 U609 ( .IN1(n447), .IN2(TxBDAddress[5]), .IN3(N804), .IN4(n448), .Q(
        n1575) );
  AO22X1 U610 ( .IN1(n447), .IN2(TxBDAddress[6]), .IN3(N805), .IN4(n448), .Q(
        n1574) );
  AO22X1 U611 ( .IN1(n447), .IN2(TxBDAddress[7]), .IN3(N806), .IN4(n448), .Q(
        n1573) );
  NOR2X0 U612 ( .IN1(n449), .IN2(n647), .QN(n448) );
  AND2X1 U613 ( .IN1(n450), .IN2(n449), .Q(n447) );
  NAND2X0 U614 ( .IN1(n451), .IN2(n450), .QN(n449) );
  NAND2X0 U615 ( .IN1(n766), .IN2(r_TxEn), .QN(n450) );
  AO221X1 U616 ( .IN1(ram_addr[0]), .IN2(n106), .IN3(WB_ADR_I[2]), .IN4(n107), 
        .IN5(n452), .Q(n1572) );
  AO22X1 U617 ( .IN1(n109), .IN2(n725), .IN3(n110), .IN4(n722), .Q(n452) );
  AO221X1 U618 ( .IN1(ram_addr[1]), .IN2(n106), .IN3(WB_ADR_I[3]), .IN4(n107), 
        .IN5(n453), .Q(n1571) );
  AO22X1 U619 ( .IN1(n109), .IN2(TxBDAddress[1]), .IN3(n110), .IN4(
        RxBDAddress[1]), .Q(n453) );
  AO221X1 U620 ( .IN1(ram_addr[2]), .IN2(n106), .IN3(WB_ADR_I[4]), .IN4(n107), 
        .IN5(n454), .Q(n1570) );
  AO22X1 U621 ( .IN1(n109), .IN2(TxBDAddress[2]), .IN3(n110), .IN4(
        RxBDAddress[2]), .Q(n454) );
  AO221X1 U622 ( .IN1(ram_addr[3]), .IN2(n106), .IN3(WB_ADR_I[5]), .IN4(n107), 
        .IN5(n455), .Q(n1569) );
  AO22X1 U623 ( .IN1(n109), .IN2(TxBDAddress[3]), .IN3(n110), .IN4(
        RxBDAddress[3]), .Q(n455) );
  AO221X1 U624 ( .IN1(ram_addr[4]), .IN2(n106), .IN3(WB_ADR_I[6]), .IN4(n107), 
        .IN5(n456), .Q(n1568) );
  AO22X1 U625 ( .IN1(n109), .IN2(TxBDAddress[4]), .IN3(n110), .IN4(
        RxBDAddress[4]), .Q(n456) );
  AO221X1 U626 ( .IN1(ram_addr[5]), .IN2(n106), .IN3(WB_ADR_I[7]), .IN4(n107), 
        .IN5(n457), .Q(n1567) );
  AO22X1 U627 ( .IN1(n109), .IN2(TxBDAddress[5]), .IN3(n110), .IN4(
        RxBDAddress[5]), .Q(n457) );
  AO221X1 U628 ( .IN1(ram_addr[6]), .IN2(n106), .IN3(WB_ADR_I[8]), .IN4(n107), 
        .IN5(n458), .Q(n1566) );
  AO22X1 U629 ( .IN1(n109), .IN2(TxBDAddress[6]), .IN3(n110), .IN4(
        RxBDAddress[6]), .Q(n458) );
  AO221X1 U630 ( .IN1(ram_addr[7]), .IN2(n106), .IN3(WB_ADR_I[9]), .IN4(n107), 
        .IN5(n459), .Q(n1565) );
  AO22X1 U631 ( .IN1(n109), .IN2(TxBDAddress[7]), .IN3(n110), .IN4(
        RxBDAddress[7]), .Q(n459) );
  NOR3X0 U632 ( .IN1(n110), .IN2(n109), .IN3(n107), .QN(n106) );
  INVX0 U633 ( .INP(n260), .ZN(n107) );
  NAND2X0 U634 ( .IN1(n460), .IN2(n744), .QN(n260) );
  MUX21X1 U635 ( .IN1(n737), .IN2(n461), .S(n745), .Q(n460) );
  OA21X1 U636 ( .IN1(n743), .IN2(n757), .IN3(n538), .Q(n461) );
  AND3X1 U637 ( .IN1(n745), .IN2(n645), .IN3(n462), .Q(n109) );
  MUX21X1 U638 ( .IN1(n463), .IN2(n757), .S(n744), .Q(n462) );
  NOR2X0 U639 ( .IN1(n732), .IN2(n757), .QN(n463) );
  NOR2X0 U640 ( .IN1(n265), .IN2(n743), .QN(n110) );
  NAND3X0 U641 ( .IN1(n737), .IN2(n734), .IN3(n745), .QN(n265) );
  AOI22X1 U642 ( .IN1(n91), .IN2(n1419), .IN3(n1452), .IN4(n1451), .QN(n1564)
         );
  AO21X1 U643 ( .IN1(n648), .IN2(n1420), .IN3(n654), .Q(n1563) );
  OA21X1 U644 ( .IN1(n648), .IN2(TxUnderRun), .IN3(n1420), .Q(n1562) );
  AO222X1 U645 ( .IN1(N350), .IN2(n464), .IN3(n465), .IN4(TxPointerMSB[2]), 
        .IN5(WB_DAT_O[2]), .IN6(n306), .Q(n1561) );
  AO222X1 U646 ( .IN1(N351), .IN2(n464), .IN3(n465), .IN4(TxPointerMSB[3]), 
        .IN5(WB_DAT_O[3]), .IN6(n306), .Q(n1560) );
  AO222X1 U647 ( .IN1(N352), .IN2(n464), .IN3(n465), .IN4(TxPointerMSB[4]), 
        .IN5(WB_DAT_O[4]), .IN6(n306), .Q(n1559) );
  AO222X1 U648 ( .IN1(N353), .IN2(n464), .IN3(n465), .IN4(TxPointerMSB[5]), 
        .IN5(WB_DAT_O[5]), .IN6(n306), .Q(n1558) );
  AO222X1 U649 ( .IN1(N354), .IN2(n464), .IN3(n465), .IN4(TxPointerMSB[6]), 
        .IN5(WB_DAT_O[6]), .IN6(n306), .Q(n1557) );
  AO222X1 U650 ( .IN1(N355), .IN2(n464), .IN3(n465), .IN4(TxPointerMSB[7]), 
        .IN5(WB_DAT_O[7]), .IN6(n306), .Q(n1556) );
  AO222X1 U651 ( .IN1(N356), .IN2(n464), .IN3(n465), .IN4(TxPointerMSB[8]), 
        .IN5(WB_DAT_O[8]), .IN6(n306), .Q(n1555) );
  AO222X1 U652 ( .IN1(N357), .IN2(n464), .IN3(n465), .IN4(TxPointerMSB[9]), 
        .IN5(WB_DAT_O[9]), .IN6(n306), .Q(n1554) );
  AO222X1 U653 ( .IN1(N358), .IN2(n464), .IN3(n465), .IN4(TxPointerMSB[10]), 
        .IN5(WB_DAT_O[10]), .IN6(n306), .Q(n1553) );
  AO222X1 U654 ( .IN1(N359), .IN2(n464), .IN3(n465), .IN4(TxPointerMSB[11]), 
        .IN5(WB_DAT_O[11]), .IN6(n306), .Q(n1552) );
  AO222X1 U655 ( .IN1(N360), .IN2(n464), .IN3(n465), .IN4(TxPointerMSB[12]), 
        .IN5(WB_DAT_O[12]), .IN6(n306), .Q(n1551) );
  AO222X1 U656 ( .IN1(N361), .IN2(n464), .IN3(n465), .IN4(TxPointerMSB[13]), 
        .IN5(WB_DAT_O[13]), .IN6(n306), .Q(n1550) );
  AO222X1 U657 ( .IN1(N362), .IN2(n464), .IN3(n465), .IN4(TxPointerMSB[14]), 
        .IN5(WB_DAT_O[14]), .IN6(n306), .Q(n1549) );
  AO222X1 U658 ( .IN1(N363), .IN2(n464), .IN3(n465), .IN4(TxPointerMSB[15]), 
        .IN5(n306), .IN6(WB_DAT_O[15]), .Q(n1548) );
  AO222X1 U659 ( .IN1(N364), .IN2(n464), .IN3(n465), .IN4(TxPointerMSB[16]), 
        .IN5(WB_DAT_O[16]), .IN6(n306), .Q(n1547) );
  AO222X1 U660 ( .IN1(N365), .IN2(n464), .IN3(n465), .IN4(TxPointerMSB[17]), 
        .IN5(WB_DAT_O[17]), .IN6(n306), .Q(n1546) );
  AO222X1 U661 ( .IN1(N366), .IN2(n464), .IN3(n465), .IN4(TxPointerMSB[18]), 
        .IN5(n306), .IN6(WB_DAT_O[18]), .Q(n1545) );
  AO222X1 U662 ( .IN1(N367), .IN2(n464), .IN3(n465), .IN4(TxPointerMSB[19]), 
        .IN5(WB_DAT_O[19]), .IN6(n306), .Q(n1544) );
  AO222X1 U663 ( .IN1(N368), .IN2(n464), .IN3(n465), .IN4(TxPointerMSB[20]), 
        .IN5(WB_DAT_O[20]), .IN6(n306), .Q(n1543) );
  AO222X1 U664 ( .IN1(N369), .IN2(n464), .IN3(n465), .IN4(TxPointerMSB[21]), 
        .IN5(WB_DAT_O[21]), .IN6(n306), .Q(n1542) );
  AO222X1 U665 ( .IN1(N370), .IN2(n464), .IN3(n465), .IN4(TxPointerMSB[22]), 
        .IN5(WB_DAT_O[22]), .IN6(n306), .Q(n1541) );
  AO222X1 U666 ( .IN1(N371), .IN2(n464), .IN3(n465), .IN4(TxPointerMSB[23]), 
        .IN5(WB_DAT_O[23]), .IN6(n306), .Q(n1540) );
  AO222X1 U667 ( .IN1(N372), .IN2(n464), .IN3(n465), .IN4(TxPointerMSB[24]), 
        .IN5(WB_DAT_O[24]), .IN6(n306), .Q(n1539) );
  AO222X1 U668 ( .IN1(N373), .IN2(n464), .IN3(n465), .IN4(TxPointerMSB[25]), 
        .IN5(WB_DAT_O[25]), .IN6(n306), .Q(n1538) );
  AO222X1 U669 ( .IN1(N374), .IN2(n464), .IN3(n465), .IN4(TxPointerMSB[26]), 
        .IN5(WB_DAT_O[26]), .IN6(n306), .Q(n1537) );
  AO222X1 U670 ( .IN1(N375), .IN2(n464), .IN3(n465), .IN4(TxPointerMSB[27]), 
        .IN5(WB_DAT_O[27]), .IN6(n306), .Q(n1536) );
  AO222X1 U671 ( .IN1(N376), .IN2(n464), .IN3(n465), .IN4(TxPointerMSB[28]), 
        .IN5(WB_DAT_O[28]), .IN6(n306), .Q(n1535) );
  AO222X1 U672 ( .IN1(N377), .IN2(n464), .IN3(n465), .IN4(TxPointerMSB[29]), 
        .IN5(WB_DAT_O[29]), .IN6(n306), .Q(n1534) );
  AO222X1 U673 ( .IN1(N378), .IN2(n464), .IN3(n465), .IN4(TxPointerMSB[30]), 
        .IN5(WB_DAT_O[30]), .IN6(n306), .Q(n1533) );
  AO222X1 U674 ( .IN1(N379), .IN2(n464), .IN3(n465), .IN4(TxPointerMSB[31]), 
        .IN5(n306), .IN6(WB_DAT_O[31]), .Q(n1532) );
  NOR2X0 U675 ( .IN1(n464), .IN2(n306), .QN(n465) );
  NOR3X0 U676 ( .IN1(n553), .IN2(n539), .IN3(n306), .QN(n464) );
  AO222X1 U677 ( .IN1(N998), .IN2(n466), .IN3(n467), .IN4(RxPointerMSB[2]), 
        .IN5(WB_DAT_O[2]), .IN6(n144), .Q(n1531) );
  AO222X1 U678 ( .IN1(N999), .IN2(n466), .IN3(n467), .IN4(RxPointerMSB[3]), 
        .IN5(WB_DAT_O[3]), .IN6(n144), .Q(n1530) );
  AO222X1 U679 ( .IN1(N1000), .IN2(n466), .IN3(n467), .IN4(RxPointerMSB[4]), 
        .IN5(WB_DAT_O[4]), .IN6(n144), .Q(n1529) );
  AO222X1 U680 ( .IN1(N1001), .IN2(n466), .IN3(n467), .IN4(RxPointerMSB[5]), 
        .IN5(WB_DAT_O[5]), .IN6(n144), .Q(n1528) );
  AO222X1 U681 ( .IN1(N1002), .IN2(n466), .IN3(n467), .IN4(RxPointerMSB[6]), 
        .IN5(WB_DAT_O[6]), .IN6(n144), .Q(n1527) );
  AO222X1 U682 ( .IN1(N1003), .IN2(n466), .IN3(n467), .IN4(RxPointerMSB[7]), 
        .IN5(WB_DAT_O[7]), .IN6(n144), .Q(n1526) );
  AO222X1 U683 ( .IN1(N1004), .IN2(n466), .IN3(n467), .IN4(RxPointerMSB[8]), 
        .IN5(WB_DAT_O[8]), .IN6(n144), .Q(n1525) );
  AO222X1 U684 ( .IN1(N1005), .IN2(n466), .IN3(n467), .IN4(RxPointerMSB[9]), 
        .IN5(WB_DAT_O[9]), .IN6(n144), .Q(n1524) );
  AO222X1 U685 ( .IN1(N1006), .IN2(n466), .IN3(n467), .IN4(RxPointerMSB[10]), 
        .IN5(WB_DAT_O[10]), .IN6(n144), .Q(n1523) );
  AO222X1 U686 ( .IN1(N1007), .IN2(n466), .IN3(n467), .IN4(RxPointerMSB[11]), 
        .IN5(WB_DAT_O[11]), .IN6(n144), .Q(n1522) );
  AO222X1 U687 ( .IN1(N1008), .IN2(n466), .IN3(n467), .IN4(RxPointerMSB[12]), 
        .IN5(WB_DAT_O[12]), .IN6(n144), .Q(n1521) );
  AO222X1 U688 ( .IN1(N1009), .IN2(n466), .IN3(n467), .IN4(RxPointerMSB[13]), 
        .IN5(WB_DAT_O[13]), .IN6(n144), .Q(n1520) );
  AO222X1 U689 ( .IN1(N1010), .IN2(n466), .IN3(n467), .IN4(RxPointerMSB[14]), 
        .IN5(WB_DAT_O[14]), .IN6(n144), .Q(n1519) );
  AO222X1 U690 ( .IN1(N1011), .IN2(n466), .IN3(n467), .IN4(RxPointerMSB[15]), 
        .IN5(WB_DAT_O[15]), .IN6(n144), .Q(n1518) );
  AO222X1 U691 ( .IN1(N1012), .IN2(n466), .IN3(n467), .IN4(RxPointerMSB[16]), 
        .IN5(WB_DAT_O[16]), .IN6(n144), .Q(n1517) );
  AO222X1 U692 ( .IN1(N1013), .IN2(n466), .IN3(n467), .IN4(RxPointerMSB[17]), 
        .IN5(WB_DAT_O[17]), .IN6(n144), .Q(n1516) );
  AO222X1 U693 ( .IN1(N1014), .IN2(n466), .IN3(n467), .IN4(RxPointerMSB[18]), 
        .IN5(WB_DAT_O[18]), .IN6(n144), .Q(n1515) );
  AO222X1 U694 ( .IN1(N1015), .IN2(n466), .IN3(n467), .IN4(RxPointerMSB[19]), 
        .IN5(WB_DAT_O[19]), .IN6(n144), .Q(n1514) );
  AO222X1 U695 ( .IN1(N1016), .IN2(n466), .IN3(n467), .IN4(RxPointerMSB[20]), 
        .IN5(WB_DAT_O[20]), .IN6(n144), .Q(n1513) );
  AO222X1 U696 ( .IN1(N1017), .IN2(n466), .IN3(n467), .IN4(RxPointerMSB[21]), 
        .IN5(WB_DAT_O[21]), .IN6(n144), .Q(n1512) );
  AO222X1 U697 ( .IN1(N1018), .IN2(n466), .IN3(n467), .IN4(RxPointerMSB[22]), 
        .IN5(WB_DAT_O[22]), .IN6(n144), .Q(n1511) );
  AO222X1 U698 ( .IN1(N1019), .IN2(n466), .IN3(n467), .IN4(RxPointerMSB[23]), 
        .IN5(WB_DAT_O[23]), .IN6(n144), .Q(n1510) );
  AO222X1 U699 ( .IN1(N1020), .IN2(n466), .IN3(n467), .IN4(RxPointerMSB[24]), 
        .IN5(WB_DAT_O[24]), .IN6(n144), .Q(n1509) );
  AO222X1 U700 ( .IN1(N1021), .IN2(n466), .IN3(n467), .IN4(RxPointerMSB[25]), 
        .IN5(WB_DAT_O[25]), .IN6(n144), .Q(n1508) );
  AO222X1 U701 ( .IN1(N1022), .IN2(n466), .IN3(n467), .IN4(RxPointerMSB[26]), 
        .IN5(WB_DAT_O[26]), .IN6(n144), .Q(n1507) );
  AO222X1 U702 ( .IN1(N1023), .IN2(n466), .IN3(n467), .IN4(RxPointerMSB[27]), 
        .IN5(WB_DAT_O[27]), .IN6(n144), .Q(n1506) );
  AO222X1 U703 ( .IN1(N1024), .IN2(n466), .IN3(n467), .IN4(RxPointerMSB[28]), 
        .IN5(WB_DAT_O[28]), .IN6(n144), .Q(n1505) );
  AO222X1 U704 ( .IN1(N1025), .IN2(n466), .IN3(n467), .IN4(RxPointerMSB[29]), 
        .IN5(WB_DAT_O[29]), .IN6(n144), .Q(n1504) );
  AO222X1 U705 ( .IN1(N1026), .IN2(n466), .IN3(n467), .IN4(RxPointerMSB[30]), 
        .IN5(WB_DAT_O[30]), .IN6(n144), .Q(n1503) );
  AO222X1 U706 ( .IN1(N1027), .IN2(n466), .IN3(n467), .IN4(RxPointerMSB[31]), 
        .IN5(n144), .IN6(WB_DAT_O[31]), .Q(n1502) );
  NOR2X0 U707 ( .IN1(n466), .IN2(n144), .QN(n467) );
  INVX0 U708 ( .INP(n95), .ZN(n144) );
  AND2X1 U709 ( .IN1(n1429), .IN2(n95), .Q(n466) );
  NAND2X0 U710 ( .IN1(n722), .IN2(n468), .QN(n95) );
  AO221X1 U711 ( .IN1(n165), .IN2(m_wb_adr_o[0]), .IN3(n469), .IN4(
        TxPointerMSB[2]), .IN5(n470), .Q(n1501) );
  AO22X1 U712 ( .IN1(n471), .IN2(RxPointerMSB[2]), .IN3(N651), .IN4(n472), .Q(
        n470) );
  AO221X1 U713 ( .IN1(n165), .IN2(m_wb_adr_o[1]), .IN3(n469), .IN4(
        TxPointerMSB[3]), .IN5(n473), .Q(n1500) );
  AO22X1 U714 ( .IN1(n471), .IN2(RxPointerMSB[3]), .IN3(N652), .IN4(n472), .Q(
        n473) );
  AO221X1 U715 ( .IN1(n165), .IN2(m_wb_adr_o[2]), .IN3(n469), .IN4(
        TxPointerMSB[4]), .IN5(n474), .Q(n1499) );
  AO22X1 U716 ( .IN1(n471), .IN2(RxPointerMSB[4]), .IN3(N653), .IN4(n472), .Q(
        n474) );
  AO221X1 U717 ( .IN1(n165), .IN2(m_wb_adr_o[3]), .IN3(n469), .IN4(
        TxPointerMSB[5]), .IN5(n475), .Q(n1498) );
  AO22X1 U718 ( .IN1(n471), .IN2(RxPointerMSB[5]), .IN3(N654), .IN4(n472), .Q(
        n475) );
  AO221X1 U719 ( .IN1(n165), .IN2(m_wb_adr_o[4]), .IN3(n469), .IN4(
        TxPointerMSB[6]), .IN5(n476), .Q(n1497) );
  AO22X1 U720 ( .IN1(n471), .IN2(RxPointerMSB[6]), .IN3(N655), .IN4(n472), .Q(
        n476) );
  AO221X1 U721 ( .IN1(n165), .IN2(m_wb_adr_o[5]), .IN3(n469), .IN4(
        TxPointerMSB[7]), .IN5(n477), .Q(n1496) );
  AO22X1 U722 ( .IN1(n471), .IN2(RxPointerMSB[7]), .IN3(N656), .IN4(n472), .Q(
        n477) );
  AO221X1 U723 ( .IN1(n165), .IN2(m_wb_adr_o[6]), .IN3(n469), .IN4(
        TxPointerMSB[8]), .IN5(n478), .Q(n1495) );
  AO22X1 U724 ( .IN1(n471), .IN2(RxPointerMSB[8]), .IN3(N657), .IN4(n472), .Q(
        n478) );
  AO221X1 U725 ( .IN1(n165), .IN2(m_wb_adr_o[7]), .IN3(n469), .IN4(
        TxPointerMSB[9]), .IN5(n479), .Q(n1494) );
  AO22X1 U726 ( .IN1(n471), .IN2(RxPointerMSB[9]), .IN3(N658), .IN4(n472), .Q(
        n479) );
  AO221X1 U727 ( .IN1(n165), .IN2(m_wb_adr_o[8]), .IN3(n469), .IN4(
        TxPointerMSB[10]), .IN5(n480), .Q(n1493) );
  AO22X1 U728 ( .IN1(n471), .IN2(RxPointerMSB[10]), .IN3(N659), .IN4(n472), 
        .Q(n480) );
  AO221X1 U729 ( .IN1(n165), .IN2(m_wb_adr_o[9]), .IN3(n469), .IN4(
        TxPointerMSB[11]), .IN5(n481), .Q(n1492) );
  AO22X1 U730 ( .IN1(n471), .IN2(RxPointerMSB[11]), .IN3(N660), .IN4(n472), 
        .Q(n481) );
  AO221X1 U731 ( .IN1(n165), .IN2(m_wb_adr_o[10]), .IN3(n469), .IN4(
        TxPointerMSB[12]), .IN5(n482), .Q(n1491) );
  AO22X1 U732 ( .IN1(n471), .IN2(RxPointerMSB[12]), .IN3(N661), .IN4(n472), 
        .Q(n482) );
  AO221X1 U733 ( .IN1(n165), .IN2(m_wb_adr_o[11]), .IN3(n469), .IN4(
        TxPointerMSB[13]), .IN5(n483), .Q(n1490) );
  AO22X1 U734 ( .IN1(n471), .IN2(RxPointerMSB[13]), .IN3(N662), .IN4(n472), 
        .Q(n483) );
  AO221X1 U735 ( .IN1(n165), .IN2(m_wb_adr_o[12]), .IN3(n469), .IN4(
        TxPointerMSB[14]), .IN5(n484), .Q(n1489) );
  AO22X1 U736 ( .IN1(n471), .IN2(RxPointerMSB[14]), .IN3(N663), .IN4(n472), 
        .Q(n484) );
  AO221X1 U737 ( .IN1(n165), .IN2(m_wb_adr_o[13]), .IN3(n469), .IN4(
        TxPointerMSB[15]), .IN5(n485), .Q(n1488) );
  AO22X1 U738 ( .IN1(n471), .IN2(RxPointerMSB[15]), .IN3(N664), .IN4(n472), 
        .Q(n485) );
  AO221X1 U739 ( .IN1(n165), .IN2(m_wb_adr_o[14]), .IN3(n469), .IN4(
        TxPointerMSB[16]), .IN5(n486), .Q(n1487) );
  AO22X1 U740 ( .IN1(n471), .IN2(RxPointerMSB[16]), .IN3(N665), .IN4(n472), 
        .Q(n486) );
  AO221X1 U741 ( .IN1(n165), .IN2(m_wb_adr_o[15]), .IN3(n469), .IN4(
        TxPointerMSB[17]), .IN5(n487), .Q(n1486) );
  AO22X1 U742 ( .IN1(n471), .IN2(RxPointerMSB[17]), .IN3(N666), .IN4(n472), 
        .Q(n487) );
  AO221X1 U743 ( .IN1(n165), .IN2(m_wb_adr_o[16]), .IN3(n469), .IN4(
        TxPointerMSB[18]), .IN5(n488), .Q(n1485) );
  AO22X1 U744 ( .IN1(n471), .IN2(RxPointerMSB[18]), .IN3(N667), .IN4(n472), 
        .Q(n488) );
  AO221X1 U745 ( .IN1(n165), .IN2(m_wb_adr_o[17]), .IN3(n469), .IN4(
        TxPointerMSB[19]), .IN5(n489), .Q(n1484) );
  AO22X1 U746 ( .IN1(n471), .IN2(RxPointerMSB[19]), .IN3(N668), .IN4(n472), 
        .Q(n489) );
  AO221X1 U747 ( .IN1(n165), .IN2(m_wb_adr_o[18]), .IN3(n469), .IN4(
        TxPointerMSB[20]), .IN5(n490), .Q(n1483) );
  AO22X1 U748 ( .IN1(n471), .IN2(RxPointerMSB[20]), .IN3(N669), .IN4(n472), 
        .Q(n490) );
  AO221X1 U749 ( .IN1(n165), .IN2(m_wb_adr_o[19]), .IN3(n469), .IN4(
        TxPointerMSB[21]), .IN5(n491), .Q(n1482) );
  AO22X1 U750 ( .IN1(n471), .IN2(RxPointerMSB[21]), .IN3(N670), .IN4(n472), 
        .Q(n491) );
  AO221X1 U751 ( .IN1(n165), .IN2(m_wb_adr_o[20]), .IN3(n469), .IN4(
        TxPointerMSB[22]), .IN5(n492), .Q(n1481) );
  AO22X1 U752 ( .IN1(n471), .IN2(RxPointerMSB[22]), .IN3(N671), .IN4(n472), 
        .Q(n492) );
  AO221X1 U753 ( .IN1(n165), .IN2(m_wb_adr_o[21]), .IN3(n469), .IN4(
        TxPointerMSB[23]), .IN5(n493), .Q(n1480) );
  AO22X1 U754 ( .IN1(n471), .IN2(RxPointerMSB[23]), .IN3(N672), .IN4(n472), 
        .Q(n493) );
  AO221X1 U755 ( .IN1(n165), .IN2(m_wb_adr_o[22]), .IN3(n469), .IN4(
        TxPointerMSB[24]), .IN5(n494), .Q(n1479) );
  AO22X1 U756 ( .IN1(n471), .IN2(RxPointerMSB[24]), .IN3(N673), .IN4(n472), 
        .Q(n494) );
  AO221X1 U757 ( .IN1(n165), .IN2(m_wb_adr_o[23]), .IN3(n469), .IN4(
        TxPointerMSB[25]), .IN5(n495), .Q(n1478) );
  AO22X1 U758 ( .IN1(n471), .IN2(RxPointerMSB[25]), .IN3(N674), .IN4(n472), 
        .Q(n495) );
  AO221X1 U759 ( .IN1(n165), .IN2(m_wb_adr_o[24]), .IN3(n469), .IN4(
        TxPointerMSB[26]), .IN5(n496), .Q(n1477) );
  AO22X1 U760 ( .IN1(n471), .IN2(RxPointerMSB[26]), .IN3(N675), .IN4(n472), 
        .Q(n496) );
  AO221X1 U761 ( .IN1(n165), .IN2(m_wb_adr_o[25]), .IN3(n469), .IN4(
        TxPointerMSB[27]), .IN5(n497), .Q(n1476) );
  AO22X1 U762 ( .IN1(n471), .IN2(RxPointerMSB[27]), .IN3(N676), .IN4(n472), 
        .Q(n497) );
  AO221X1 U763 ( .IN1(n165), .IN2(m_wb_adr_o[26]), .IN3(n469), .IN4(
        TxPointerMSB[28]), .IN5(n498), .Q(n1475) );
  AO22X1 U764 ( .IN1(n471), .IN2(RxPointerMSB[28]), .IN3(N677), .IN4(n472), 
        .Q(n498) );
  AO221X1 U765 ( .IN1(n165), .IN2(m_wb_adr_o[27]), .IN3(n469), .IN4(
        TxPointerMSB[29]), .IN5(n499), .Q(n1474) );
  AO22X1 U766 ( .IN1(n471), .IN2(RxPointerMSB[29]), .IN3(N678), .IN4(n472), 
        .Q(n499) );
  AO221X1 U767 ( .IN1(n165), .IN2(m_wb_adr_o[28]), .IN3(n469), .IN4(
        TxPointerMSB[30]), .IN5(n500), .Q(n1473) );
  AO22X1 U768 ( .IN1(n471), .IN2(RxPointerMSB[30]), .IN3(N679), .IN4(n472), 
        .Q(n500) );
  AO221X1 U769 ( .IN1(n165), .IN2(m_wb_adr_o[29]), .IN3(n469), .IN4(
        TxPointerMSB[31]), .IN5(n501), .Q(n1472) );
  AO22X1 U770 ( .IN1(n471), .IN2(RxPointerMSB[31]), .IN3(N680), .IN4(n472), 
        .Q(n501) );
  NAND3X0 U771 ( .IN1(n233), .IN2(n241), .IN3(n239), .QN(n472) );
  OA22X1 U772 ( .IN1(n5), .IN2(n235), .IN3(n2), .IN4(n502), .Q(n239) );
  AOI22X1 U773 ( .IN1(n126), .IN2(tx_burst_cnt[2]), .IN3(rx_burst_cnt[2]), 
        .IN4(n238), .QN(n241) );
  OA21X1 U774 ( .IN1(n7), .IN2(n502), .IN3(n132), .Q(n233) );
  NAND2X0 U775 ( .IN1(tx_burst_cnt[0]), .IN2(n126), .QN(n132) );
  INVX0 U776 ( .INP(n235), .ZN(n126) );
  NAND2X0 U777 ( .IN1(n503), .IN2(n504), .QN(n471) );
  NAND4X0 U778 ( .IN1(n238), .IN2(n7), .IN3(n2), .IN4(n1), .QN(n504) );
  INVX0 U779 ( .INP(n502), .ZN(n238) );
  NAND2X0 U780 ( .IN1(n505), .IN2(n506), .QN(n469) );
  OR4X1 U781 ( .IN1(n235), .IN2(tx_burst_cnt[0]), .IN3(tx_burst_cnt[1]), .IN4(
        tx_burst_cnt[2]), .Q(n506) );
  INVX0 U782 ( .INP(n243), .ZN(n165) );
  NAND2X0 U783 ( .IN1(n162), .IN2(n225), .QN(n243) );
  INVX0 U784 ( .INP(n245), .ZN(n225) );
  NAND2X0 U785 ( .IN1(n505), .IN2(n235), .QN(n245) );
  NAND3X0 U786 ( .IN1(n237), .IN2(n507), .IN3(tx_burst_en), .QN(n235) );
  NAND3X0 U787 ( .IN1(n236), .IN2(n232), .IN3(n508), .QN(n507) );
  NAND3X0 U788 ( .IN1(n117), .IN2(n251), .IN3(n551), .QN(n508) );
  NOR2X0 U789 ( .IN1(n728), .IN2(n550), .QN(n117) );
  NAND3X0 U790 ( .IN1(n509), .IN2(n6), .IN3(n237), .QN(n505) );
  NAND2X0 U791 ( .IN1(n236), .IN2(n232), .QN(n509) );
  NAND3X0 U792 ( .IN1(n249), .IN2(n510), .IN3(n257), .QN(n232) );
  NAND2X0 U793 ( .IN1(n253), .IN2(n727), .QN(n510) );
  OR2X1 U794 ( .IN1(n511), .IN2(n253), .Q(n236) );
  INVX0 U795 ( .INP(n242), .ZN(n162) );
  NAND2X0 U796 ( .IN1(n503), .IN2(n502), .QN(n242) );
  NAND3X0 U797 ( .IN1(rx_burst_en), .IN2(n253), .IN3(n512), .QN(n502) );
  MUX21X1 U798 ( .IN1(n513), .IN2(n514), .S(n550), .Q(n512) );
  AO22X1 U799 ( .IN1(n515), .IN2(n540), .IN3(n516), .IN4(n257), .Q(n514) );
  NOR2X0 U800 ( .IN1(n551), .IN2(n237), .QN(n516) );
  XOR2X1 U801 ( .IN1(n251), .IN2(n551), .Q(n515) );
  AND2X1 U802 ( .IN1(n551), .IN2(n257), .Q(n513) );
  OA21X1 U803 ( .IN1(n511), .IN2(RxBufferEmpty), .IN3(n231), .Q(n503) );
  NAND4X0 U804 ( .IN1(n257), .IN2(n249), .IN3(n517), .IN4(n518), .QN(n231) );
  NAND2X0 U805 ( .IN1(n237), .IN2(n550), .QN(n518) );
  NOR2X0 U806 ( .IN1(n533), .IN2(n653), .QN(n237) );
  NOR2X0 U807 ( .IN1(rx_burst_en), .IN2(RxBufferEmpty), .QN(n517) );
  XOR2X1 U808 ( .IN1(n551), .IN2(n550), .Q(n249) );
  NOR2X0 U809 ( .IN1(n251), .IN2(n540), .QN(n257) );
  INVX0 U810 ( .INP(n258), .ZN(n251) );
  NAND4X0 U811 ( .IN1(n258), .IN2(n252), .IN3(n551), .IN4(n550), .QN(n511) );
  AOI21X1 U812 ( .IN1(rx_burst_en), .IN2(n253), .IN3(n728), .QN(n252) );
  INVX0 U813 ( .INP(RxBufferEmpty), .ZN(n253) );
  OA21X1 U814 ( .IN1(n152), .IN2(RxStatusWriteLatched), .IN3(n860), .Q(n1471)
         );
  AO22X1 U815 ( .IN1(n1469), .IN2(Busy_IRQ_rck), .IN3(n200), .IN4(n8), .Q(
        n1470) );
  INVX0 U816 ( .INP(n207), .ZN(n200) );
  NAND2X0 U817 ( .IN1(RxStartFrm), .IN2(RxValid), .QN(n207) );
  AND2X1 U818 ( .IN1(m_wb_ack_i), .IN2(n635), .Q(n1429) );
  MUX21X1 U819 ( .IN1(n684), .IN2(RxLength[15]), .S(LoadRxStatus), .Q(n1384)
         );
  MUX21X1 U820 ( .IN1(n683), .IN2(RxLength[14]), .S(LoadRxStatus), .Q(n1382)
         );
  MUX21X1 U821 ( .IN1(n682), .IN2(RxLength[13]), .S(LoadRxStatus), .Q(n1380)
         );
  MUX21X1 U822 ( .IN1(n681), .IN2(RxLength[12]), .S(LoadRxStatus), .Q(n1378)
         );
  MUX21X1 U823 ( .IN1(n680), .IN2(RxLength[11]), .S(LoadRxStatus), .Q(n1376)
         );
  MUX21X1 U824 ( .IN1(n678), .IN2(RxLength[10]), .S(LoadRxStatus), .Q(n1374)
         );
  MUX21X1 U825 ( .IN1(n677), .IN2(RxLength[9]), .S(LoadRxStatus), .Q(n1372) );
  MUX21X1 U826 ( .IN1(n675), .IN2(RxLength[8]), .S(LoadRxStatus), .Q(n1370) );
  MUX21X1 U827 ( .IN1(n673), .IN2(RxLength[7]), .S(LoadRxStatus), .Q(n1368) );
  MUX21X1 U828 ( .IN1(n672), .IN2(RxLength[6]), .S(LoadRxStatus), .Q(n1366) );
  MUX21X1 U829 ( .IN1(n671), .IN2(RxLength[5]), .S(LoadRxStatus), .Q(n1364) );
  MUX21X1 U830 ( .IN1(n670), .IN2(RxLength[4]), .S(LoadRxStatus), .Q(n1362) );
  MUX21X1 U831 ( .IN1(n669), .IN2(RxLength[3]), .S(LoadRxStatus), .Q(n1360) );
  MUX21X1 U832 ( .IN1(n668), .IN2(RxLength[2]), .S(LoadRxStatus), .Q(n1358) );
  MUX21X1 U833 ( .IN1(n667), .IN2(RxLength[1]), .S(LoadRxStatus), .Q(n1356) );
  MUX21X1 U834 ( .IN1(n666), .IN2(RxLength[0]), .S(LoadRxStatus), .Q(n1354) );
  MUX21X1 U835 ( .IN1(n665), .IN2(ReceivedPauseFrm), .S(LoadRxStatus), .Q(
        n1352) );
  MUX21X1 U836 ( .IN1(n664), .IN2(AddressMiss), .S(LoadRxStatus), .Q(n1350) );
  MUX21X1 U837 ( .IN1(n663), .IN2(InvalidSymbol), .S(LoadRxStatus), .Q(n1348)
         );
  MUX21X1 U838 ( .IN1(n662), .IN2(DribbleNibble), .S(LoadRxStatus), .Q(n1346)
         );
  MUX21X1 U839 ( .IN1(n661), .IN2(ReceivedPacketTooBig), .S(LoadRxStatus), .Q(
        n1344) );
  MUX21X1 U840 ( .IN1(n660), .IN2(ShortFrame), .S(LoadRxStatus), .Q(n1342) );
  MUX21X1 U841 ( .IN1(n659), .IN2(LatchedCrcError), .S(LoadRxStatus), .Q(n1340) );
  MUX21X1 U842 ( .IN1(n658), .IN2(RxLateCollision), .S(LoadRxStatus), .Q(n1338) );
  MUX21X1 U843 ( .IN1(n656), .IN2(n657), .S(LoadRxStatus), .Q(n1335) );
  MUX21X1 U844 ( .IN1(PerPacketCrcEn), .IN2(WB_DAT_O[11]), .S(n111), .Q(n1301)
         );
  MUX21X1 U845 ( .IN1(PerPacketPad), .IN2(WB_DAT_O[12]), .S(n111), .Q(n1299)
         );
  MUX21X1 U846 ( .IN1(n647), .IN2(WB_DAT_O[13]), .S(n111), .Q(n1297) );
  MUX21X1 U847 ( .IN1(n646), .IN2(WB_DAT_O[14]), .S(n111), .Q(n1288) );
  MUX21X1 U848 ( .IN1(n639), .IN2(WB_DAT_O[14]), .S(n97), .Q(n1266) );
  MUX21X1 U849 ( .IN1(n638), .IN2(WB_DAT_O[13]), .S(n97), .Q(n1264) );
  AND2X1 U850 ( .IN1(n697), .IN2(n468), .Q(n97) );
  INVX0 U851 ( .INP(n153), .ZN(n468) );
  NOR2X0 U852 ( .IN1(n730), .IN2(n729), .QN(n124) );
  MUX21X1 U853 ( .IN1(n688), .IN2(WB_DAT_O[1]), .S(n306), .Q(n1159) );
  MUX21X1 U854 ( .IN1(n689), .IN2(WB_DAT_O[0]), .S(n306), .Q(n1157) );
  INVX0 U855 ( .INP(n93), .ZN(n306) );
  NAND2X0 U856 ( .IN1(n725), .IN2(n304), .QN(n93) );
  MUX21X1 U857 ( .IN1(n607), .IN2(WB_DAT_O[31]), .S(n111), .Q(n1133) );
  MUX21X1 U858 ( .IN1(n606), .IN2(WB_DAT_O[30]), .S(n111), .Q(n1130) );
  MUX21X1 U859 ( .IN1(n605), .IN2(WB_DAT_O[29]), .S(n111), .Q(n1127) );
  MUX21X1 U860 ( .IN1(n604), .IN2(WB_DAT_O[28]), .S(n111), .Q(n1124) );
  MUX21X1 U861 ( .IN1(n603), .IN2(WB_DAT_O[27]), .S(n111), .Q(n1121) );
  MUX21X1 U862 ( .IN1(n602), .IN2(WB_DAT_O[26]), .S(n111), .Q(n1118) );
  MUX21X1 U863 ( .IN1(n601), .IN2(WB_DAT_O[25]), .S(n111), .Q(n1115) );
  MUX21X1 U864 ( .IN1(n600), .IN2(WB_DAT_O[24]), .S(n111), .Q(n1112) );
  MUX21X1 U865 ( .IN1(n599), .IN2(WB_DAT_O[23]), .S(n111), .Q(n1109) );
  MUX21X1 U866 ( .IN1(n598), .IN2(WB_DAT_O[22]), .S(n111), .Q(n1106) );
  MUX21X1 U867 ( .IN1(n597), .IN2(WB_DAT_O[21]), .S(n111), .Q(n1103) );
  MUX21X1 U868 ( .IN1(n596), .IN2(WB_DAT_O[20]), .S(n111), .Q(n1100) );
  MUX21X1 U869 ( .IN1(n595), .IN2(WB_DAT_O[19]), .S(n111), .Q(n1097) );
  MUX21X1 U870 ( .IN1(n594), .IN2(WB_DAT_O[18]), .S(n111), .Q(n1094) );
  MUX21X1 U871 ( .IN1(n593), .IN2(WB_DAT_O[17]), .S(n111), .Q(n1091) );
  MUX21X1 U872 ( .IN1(n592), .IN2(WB_DAT_O[16]), .S(n111), .Q(n1088) );
  NAND2X0 U873 ( .IN1(n731), .IN2(n304), .QN(n94) );
  NOR3X0 U874 ( .IN1(n556), .IN2(n1463), .IN3(RxBufferFull), .QN(_2_net_) );
  NOR2X0 U875 ( .IN1(TxBufferEmpty), .IN2(n123), .QN(_1_net_) );
  NAND2X0 U876 ( .IN1(ReadTxDataFromFifo_sync2), .IN2(n1449), .QN(n123) );
  NOR2X0 U877 ( .IN1(n1420), .IN2(BlockingTxStatusWrite_sync3), .QN(
        RstDeferLatched) );
  NOR3X0 U878 ( .IN1(n519), .IN2(n1451), .IN3(n651), .QN(N857) );
  NOR3X0 U879 ( .IN1(n1450), .IN2(n650), .IN3(n519), .QN(N848) );
  NOR3X0 U880 ( .IN1(n1452), .IN2(n649), .IN3(n519), .QN(N837) );
  OA21X1 U881 ( .IN1(tx_burst_en), .IN2(n258), .IN3(n727), .Q(n519) );
  NOR2X0 U882 ( .IN1(m_wb_err_i), .IN2(m_wb_ack_i), .QN(n258) );
  NOR2X0 U883 ( .IN1(n746), .IN2(n355), .QN(N792) );
  NAND4X0 U884 ( .IN1(n709), .IN2(n708), .IN3(n707), .IN4(n133), .QN(n355) );
  INVX0 U885 ( .INP(n122), .ZN(n133) );
  NAND4X0 U886 ( .IN1(n712), .IN2(n711), .IN3(n520), .IN4(n521), .QN(n122) );
  NOR4X0 U887 ( .IN1(n36), .IN2(n522), .IN3(n43), .IN4(n32), .QN(n521) );
  NAND2X0 U888 ( .IN1(n714), .IN2(n713), .QN(n522) );
  NOR3X0 U889 ( .IN1(n29), .IN2(n350), .IN3(n54), .QN(n520) );
  NAND2X0 U890 ( .IN1(n717), .IN2(n716), .QN(n350) );
  AO22X1 U891 ( .IN1(n89), .IN2(n523), .IN3(n524), .IN4(n608), .Q(N76) );
  INVX0 U892 ( .INP(n142), .ZN(n524) );
  NAND2X0 U893 ( .IN1(n744), .IN2(WbEn), .QN(n142) );
  OR4X1 U894 ( .IN1(n641), .IN2(n642), .IN3(n643), .IN4(n644), .Q(n523) );
  NOR2X0 U895 ( .IN1(n838), .IN2(n744), .QN(n89) );
  NOR4X0 U896 ( .IN1(n674), .IN2(n525), .IN3(n526), .IN4(n92), .QN(N1268) );
  NOR4X0 U897 ( .IN1(n527), .IN2(n92), .IN3(n674), .IN4(n526), .QN(N1265) );
  OA21X1 U898 ( .IN1(n528), .IN2(r_RxFlow), .IN3(ReceivedPauseFrm), .Q(n526)
         );
  INVX0 U899 ( .INP(r_PassAll), .ZN(n528) );
  INVX0 U900 ( .INP(n152), .ZN(n92) );
  NOR2X0 U901 ( .IN1(n153), .IN2(n687), .QN(n152) );
  NAND2X0 U902 ( .IN1(n757), .IN2(RxEn), .QN(n153) );
  NAND2X0 U903 ( .IN1(ReceivedPacketGood), .IN2(n525), .QN(n527) );
  NOR4X0 U904 ( .IN1(n658), .IN2(n659), .IN3(n656), .IN4(n529), .QN(n525) );
  OR3X1 U905 ( .IN1(n661), .IN2(n663), .IN3(n662), .Q(n529) );
  NOR3X0 U906 ( .IN1(n91), .IN2(n530), .IN3(n10), .QN(N1261) );
  AND3X1 U907 ( .IN1(n530), .IN2(n646), .IN3(n451), .Q(N1258) );
  INVX0 U908 ( .INP(n91), .ZN(n451) );
  NAND3X0 U909 ( .IN1(n304), .IN2(n531), .IN3(n1419), .QN(n91) );
  NAND2X0 U910 ( .IN1(n747), .IN2(n13), .QN(n531) );
  NOR2X0 U911 ( .IN1(n883), .IN2(n745), .QN(n304) );
  NOR4X0 U912 ( .IN1(TxUnderRun), .IN2(CarrierSenseLost), .IN3(LateCollLatched), .IN4(RetryLimit), .QN(n530) );
  NOR2X0 U913 ( .IN1(n1468), .IN2(Busy_IRQ_sync3), .QN(Busy_IRQ) );
endmodule


module eth_macstatus_test_1 ( MRxClk, Reset, ReceivedLengthOK, ReceiveEnd, 
        ReceivedPacketGood, RxCrcError, MRxErr, MRxDV, RxStateSFD, RxStateData, 
        RxStatePreamble, RxStateIdle, Transmitting, RxByteCnt, RxByteCntEq0, 
        RxByteCntGreat2, RxByteCntMaxFrame, InvalidSymbol, MRxD, 
        LatchedCrcError, Collision, CollValid, RxLateCollision, r_RecSmall, 
        r_MinFL, r_MaxFL, ShortFrame, DribbleNibble, ReceivedPacketTooBig, 
        r_HugEn, LoadRxStatus, StartTxDone, StartTxAbort, RetryCnt, 
        RetryCntLatched, MTxClk, MaxCollisionOccured, RetryLimit, 
        LateCollision, LateCollLatched, DeferIndication, DeferLatched, 
        RstDeferLatched, TxStartFrm, StatePreamble, StateData, CarrierSense, 
        CarrierSenseLost, TxUsedData, LatchedMRxErr, Loopback, r_FullD, 
        eth_top_test_point_11887_in, test_si, test_se );
  input [1:0] RxStateData;
  input [15:0] RxByteCnt;
  input [3:0] MRxD;
  input [5:0] CollValid;
  input [15:0] r_MinFL;
  input [15:0] r_MaxFL;
  input [3:0] RetryCnt;
  output [3:0] RetryCntLatched;
  input [1:0] StateData;
  input MRxClk, Reset, RxCrcError, MRxErr, MRxDV, RxStateSFD, RxStatePreamble,
         RxStateIdle, Transmitting, RxByteCntEq0, RxByteCntGreat2,
         RxByteCntMaxFrame, Collision, r_RecSmall, r_HugEn, StartTxDone,
         StartTxAbort, MTxClk, MaxCollisionOccured, LateCollision,
         DeferIndication, RstDeferLatched, TxStartFrm, StatePreamble,
         CarrierSense, TxUsedData, Loopback, r_FullD,
         eth_top_test_point_11887_in, test_si, test_se;
  output ReceivedLengthOK, ReceiveEnd, ReceivedPacketGood, InvalidSymbol,
         LatchedCrcError, RxLateCollision, ShortFrame, DribbleNibble,
         ReceivedPacketTooBig, LoadRxStatus, RetryLimit, LateCollLatched,
         DeferLatched, CarrierSenseLost, LatchedMRxErr;
  wire   N7, TakeSample, n42, n43, n44, n45, n50, n52, n54, n56, n58, n60, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n138, n139, n140, n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n46, n47, n48, n49,
         n51, n53, n55, n57, n59, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120;

  SDFFARX1 LatchedCrcError_reg ( .D(n82), .SI(InvalidSymbol), .SE(test_se), 
        .CLK(MRxClk), .RSTB(n120), .Q(LatchedCrcError), .QN(ReceivedPacketGood) );
  SDFFARX1 LatchedMRxErr_reg ( .D(N7), .SI(LatchedCrcError), .SE(test_se), 
        .CLK(MRxClk), .RSTB(n120), .Q(LatchedMRxErr) );
  SDFFARX1 LoadRxStatus_reg ( .D(TakeSample), .SI(LateCollLatched), .SE(
        test_se), .CLK(MRxClk), .RSTB(n120), .Q(LoadRxStatus), .QN(n73) );
  SDFFARX1 ReceiveEnd_reg ( .D(LoadRxStatus), .SI(LoadRxStatus), .SE(test_se), 
        .CLK(MRxClk), .RSTB(n120), .Q(ReceiveEnd) );
  SDFFARX1 InvalidSymbol_reg ( .D(n81), .SI(DribbleNibble), .SE(test_se), 
        .CLK(MRxClk), .RSTB(n120), .Q(InvalidSymbol), .QN(n42) );
  SDFFASX1 RxColWindow_reg ( .D(n80), .SI(RetryLimit), .SE(test_se), .CLK(
        MRxClk), .SETB(n120), .Q(n138), .QN(n119) );
  SDFFARX1 RxLateCollision_reg ( .D(n79), .SI(n138), .SE(test_se), .CLK(MRxClk), .RSTB(n120), .Q(RxLateCollision) );
  SDFFARX1 ShortFrame_reg ( .D(n78), .SI(RxLateCollision), .SE(test_se), .CLK(
        MRxClk), .RSTB(n120), .Q(ShortFrame), .QN(n140) );
  SDFFARX1 DribbleNibble_reg ( .D(n77), .SI(DeferLatched), .SE(test_se), .CLK(
        MRxClk), .RSTB(n120), .Q(DribbleNibble), .QN(n43) );
  SDFFARX1 ReceivedPacketTooBig_reg ( .D(n76), .SI(ReceiveEnd), .SE(test_se), 
        .CLK(MRxClk), .RSTB(n120), .Q(ReceivedPacketTooBig), .QN(n139) );
  SDFFARX1 \RetryCntLatched_reg[3]  ( .D(n60), .SI(RetryCntLatched[2]), .SE(
        test_se), .CLK(MTxClk), .RSTB(n120), .Q(RetryCntLatched[3]) );
  SDFFARX1 \RetryCntLatched_reg[2]  ( .D(n58), .SI(RetryCntLatched[1]), .SE(
        test_se), .CLK(MTxClk), .RSTB(n120), .Q(RetryCntLatched[2]) );
  SDFFARX1 \RetryCntLatched_reg[1]  ( .D(n56), .SI(RetryCntLatched[0]), .SE(
        test_se), .CLK(MTxClk), .RSTB(n120), .Q(RetryCntLatched[1]) );
  SDFFARX1 \RetryCntLatched_reg[0]  ( .D(n54), .SI(ReceivedPacketTooBig), .SE(
        test_se), .CLK(MTxClk), .RSTB(n120), .Q(RetryCntLatched[0]) );
  SDFFARX1 RetryLimit_reg ( .D(n52), .SI(RetryCntLatched[3]), .SE(test_se), 
        .CLK(MTxClk), .RSTB(n120), .Q(RetryLimit) );
  SDFFARX1 LateCollLatched_reg ( .D(n50), .SI(LatchedMRxErr), .SE(test_se), 
        .CLK(MTxClk), .RSTB(n120), .Q(LateCollLatched) );
  SDFFARX1 DeferLatched_reg ( .D(n75), .SI(CarrierSenseLost), .SE(test_se), 
        .CLK(MTxClk), .RSTB(n120), .Q(DeferLatched), .QN(n44) );
  SDFFARX1 CarrierSenseLost_reg ( .D(n74), .SI(test_si), .SE(test_se), .CLK(
        MTxClk), .RSTB(n120), .Q(CarrierSenseLost), .QN(n45) );
  INVX0 U3 ( .INP(eth_top_test_point_11887_in), .ZN(n120) );
  NOR2X0 U4 ( .IN1(RxStateSFD), .IN2(n1), .QN(n82) );
  MUX21X1 U5 ( .IN1(ReceivedPacketGood), .IN2(n2), .S(RxStateData[0]), .Q(n1)
         );
  NAND2X0 U6 ( .IN1(RxCrcError), .IN2(n3), .QN(n2) );
  INVX0 U7 ( .INP(RxByteCntEq0), .ZN(n3) );
  OAI22X1 U8 ( .IN1(n42), .IN2(n4), .IN3(n5), .IN4(n6), .QN(n81) );
  NAND3X0 U9 ( .IN1(MRxD[3]), .IN2(MRxD[2]), .IN3(MRxErr), .QN(n6) );
  NAND2X0 U10 ( .IN1(n7), .IN2(MRxD[1]), .QN(n5) );
  NOR2X0 U11 ( .IN1(MRxD[0]), .IN2(n8), .QN(n7) );
  OA22X1 U12 ( .IN1(n9), .IN2(n10), .IN3(RxStateIdle), .IN4(n138), .Q(n80) );
  NAND4X0 U13 ( .IN1(n11), .IN2(n12), .IN3(n13), .IN4(n14), .QN(n10) );
  XOR2X1 U14 ( .IN1(n15), .IN2(CollValid[2]), .Q(n14) );
  XOR2X1 U15 ( .IN1(n16), .IN2(CollValid[3]), .Q(n13) );
  XOR2X1 U16 ( .IN1(n17), .IN2(CollValid[4]), .Q(n12) );
  XOR2X1 U17 ( .IN1(n18), .IN2(CollValid[5]), .Q(n11) );
  NAND4X0 U18 ( .IN1(n19), .IN2(n20), .IN3(RxStateData[1]), .IN4(n21), .QN(n9)
         );
  XOR2X1 U19 ( .IN1(n22), .IN2(CollValid[0]), .Q(n20) );
  XOR2X1 U20 ( .IN1(n23), .IN2(CollValid[1]), .Q(n19) );
  OA21X1 U21 ( .IN1(n24), .IN2(RxLateCollision), .IN3(n73), .Q(n79) );
  NOR3X0 U22 ( .IN1(n21), .IN2(r_FullD), .IN3(n25), .QN(n24) );
  NOR2X0 U23 ( .IN1(n119), .IN2(r_RecSmall), .QN(n25) );
  INVX0 U24 ( .INP(Collision), .ZN(n21) );
  NOR2X0 U25 ( .IN1(n4), .IN2(n26), .QN(n78) );
  MUX21X1 U26 ( .IN1(n140), .IN2(n27), .S(TakeSample), .Q(n26) );
  NOR2X0 U27 ( .IN1(RxStateSFD), .IN2(n28), .QN(n77) );
  OA21X1 U28 ( .IN1(MRxDV), .IN2(n29), .IN3(n43), .Q(n28) );
  INVX0 U29 ( .INP(RxStateData[1]), .ZN(n29) );
  NOR2X0 U30 ( .IN1(n4), .IN2(n30), .QN(n76) );
  MUX21X1 U31 ( .IN1(n139), .IN2(n31), .S(TakeSample), .Q(n30) );
  OR2X1 U32 ( .IN1(r_HugEn), .IN2(n32), .Q(n31) );
  INVX0 U33 ( .INP(n73), .ZN(n4) );
  OR2X1 U34 ( .IN1(n33), .IN2(DeferIndication), .Q(n75) );
  NOR2X0 U35 ( .IN1(n44), .IN2(RstDeferLatched), .QN(n33) );
  OAI21X1 U36 ( .IN1(n45), .IN2(TxStartFrm), .IN3(n34), .QN(n74) );
  OR4X1 U37 ( .IN1(CarrierSense), .IN2(n35), .IN3(Collision), .IN4(n36), .Q(
        n34) );
  OR2X1 U38 ( .IN1(r_FullD), .IN2(Loopback), .Q(n36) );
  NOR3X0 U39 ( .IN1(StateData[0]), .IN2(StatePreamble), .IN3(StateData[1]), 
        .QN(n35) );
  MUX21X1 U40 ( .IN1(RetryCnt[3]), .IN2(RetryCntLatched[3]), .S(n37), .Q(n60)
         );
  MUX21X1 U41 ( .IN1(RetryCnt[2]), .IN2(RetryCntLatched[2]), .S(n37), .Q(n58)
         );
  MUX21X1 U42 ( .IN1(RetryCnt[1]), .IN2(RetryCntLatched[1]), .S(n37), .Q(n56)
         );
  MUX21X1 U43 ( .IN1(RetryCnt[0]), .IN2(RetryCntLatched[0]), .S(n37), .Q(n54)
         );
  MUX21X1 U44 ( .IN1(MaxCollisionOccured), .IN2(RetryLimit), .S(n37), .Q(n52)
         );
  MUX21X1 U45 ( .IN1(LateCollision), .IN2(LateCollLatched), .S(n37), .Q(n50)
         );
  NOR2X0 U46 ( .IN1(StartTxDone), .IN2(StartTxAbort), .QN(n37) );
  AO22X1 U47 ( .IN1(RxByteCntMaxFrame), .IN2(RxStateData[0]), .IN3(n38), .IN4(
        n8), .Q(TakeSample) );
  INVX0 U48 ( .INP(MRxDV), .ZN(n8) );
  AND2X1 U49 ( .IN1(n27), .IN2(n32), .Q(ReceivedLengthOK) );
  AO21X1 U50 ( .IN1(r_MaxFL[15]), .IN2(n39), .IN3(n40), .Q(n32) );
  OA22X1 U51 ( .IN1(r_MaxFL[15]), .IN2(n39), .IN3(n41), .IN4(n46), .Q(n40) );
  AND2X1 U52 ( .IN1(n47), .IN2(r_MaxFL[14]), .Q(n46) );
  OA221X1 U53 ( .IN1(r_MaxFL[13]), .IN2(n48), .IN3(r_MaxFL[14]), .IN4(n47), 
        .IN5(n49), .Q(n41) );
  AO221X1 U54 ( .IN1(r_MaxFL[12]), .IN2(n51), .IN3(r_MaxFL[13]), .IN4(n48), 
        .IN5(n53), .Q(n49) );
  OA221X1 U55 ( .IN1(r_MaxFL[12]), .IN2(n51), .IN3(r_MaxFL[11]), .IN4(n55), 
        .IN5(n57), .Q(n53) );
  AO221X1 U56 ( .IN1(r_MaxFL[10]), .IN2(n59), .IN3(r_MaxFL[11]), .IN4(n55), 
        .IN5(n61), .Q(n57) );
  OA221X1 U57 ( .IN1(r_MaxFL[10]), .IN2(n59), .IN3(r_MaxFL[9]), .IN4(n62), 
        .IN5(n63), .Q(n61) );
  AO221X1 U58 ( .IN1(r_MaxFL[8]), .IN2(n64), .IN3(r_MaxFL[9]), .IN4(n62), 
        .IN5(n65), .Q(n63) );
  OA221X1 U59 ( .IN1(r_MaxFL[8]), .IN2(n64), .IN3(r_MaxFL[7]), .IN4(n66), 
        .IN5(n67), .Q(n65) );
  AO221X1 U60 ( .IN1(r_MaxFL[6]), .IN2(n68), .IN3(r_MaxFL[7]), .IN4(n66), 
        .IN5(n69), .Q(n67) );
  OA221X1 U61 ( .IN1(r_MaxFL[6]), .IN2(n68), .IN3(r_MaxFL[5]), .IN4(n18), 
        .IN5(n70), .Q(n69) );
  AO221X1 U62 ( .IN1(r_MaxFL[4]), .IN2(n17), .IN3(r_MaxFL[5]), .IN4(n18), 
        .IN5(n71), .Q(n70) );
  OA221X1 U63 ( .IN1(r_MaxFL[4]), .IN2(n17), .IN3(r_MaxFL[3]), .IN4(n16), 
        .IN5(n72), .Q(n71) );
  AO222X1 U64 ( .IN1(n83), .IN2(n15), .IN3(r_MaxFL[2]), .IN4(n84), .IN5(
        r_MaxFL[3]), .IN6(n16), .Q(n72) );
  OR2X1 U65 ( .IN1(n83), .IN2(n15), .Q(n84) );
  AO21X1 U66 ( .IN1(r_MaxFL[1]), .IN2(n23), .IN3(n85), .Q(n83) );
  OA22X1 U67 ( .IN1(r_MaxFL[1]), .IN2(n23), .IN3(r_MaxFL[0]), .IN4(n22), .Q(
        n85) );
  INVX0 U68 ( .INP(RxByteCnt[7]), .ZN(n66) );
  INVX0 U69 ( .INP(RxByteCnt[8]), .ZN(n64) );
  INVX0 U70 ( .INP(RxByteCnt[9]), .ZN(n62) );
  INVX0 U71 ( .INP(RxByteCnt[10]), .ZN(n59) );
  INVX0 U72 ( .INP(RxByteCnt[11]), .ZN(n55) );
  INVX0 U73 ( .INP(RxByteCnt[12]), .ZN(n51) );
  INVX0 U74 ( .INP(RxByteCnt[13]), .ZN(n48) );
  INVX0 U75 ( .INP(RxByteCnt[15]), .ZN(n39) );
  AO21X1 U76 ( .IN1(RxByteCnt[15]), .IN2(n86), .IN3(n87), .Q(n27) );
  OA22X1 U77 ( .IN1(RxByteCnt[15]), .IN2(n86), .IN3(n88), .IN4(n89), .Q(n87)
         );
  OA221X1 U78 ( .IN1(RxByteCnt[14]), .IN2(n90), .IN3(RxByteCnt[13]), .IN4(n91), 
        .IN5(n92), .Q(n89) );
  AO221X1 U79 ( .IN1(RxByteCnt[13]), .IN2(n91), .IN3(RxByteCnt[12]), .IN4(n93), 
        .IN5(n94), .Q(n92) );
  OA221X1 U80 ( .IN1(RxByteCnt[12]), .IN2(n93), .IN3(RxByteCnt[11]), .IN4(n95), 
        .IN5(n96), .Q(n94) );
  AO221X1 U81 ( .IN1(RxByteCnt[11]), .IN2(n95), .IN3(RxByteCnt[10]), .IN4(n97), 
        .IN5(n98), .Q(n96) );
  OA221X1 U82 ( .IN1(RxByteCnt[9]), .IN2(n99), .IN3(RxByteCnt[10]), .IN4(n97), 
        .IN5(n100), .Q(n98) );
  AO221X1 U83 ( .IN1(RxByteCnt[9]), .IN2(n99), .IN3(RxByteCnt[8]), .IN4(n101), 
        .IN5(n102), .Q(n100) );
  OA221X1 U84 ( .IN1(RxByteCnt[8]), .IN2(n101), .IN3(RxByteCnt[7]), .IN4(n103), 
        .IN5(n104), .Q(n102) );
  AO221X1 U85 ( .IN1(RxByteCnt[7]), .IN2(n103), .IN3(RxByteCnt[6]), .IN4(n105), 
        .IN5(n106), .Q(n104) );
  AOI222X1 U86 ( .IN1(r_MinFL[6]), .IN2(n68), .IN3(r_MinFL[5]), .IN4(n107), 
        .IN5(n108), .IN6(n18), .QN(n106) );
  OR2X1 U87 ( .IN1(n108), .IN2(n18), .Q(n107) );
  INVX0 U88 ( .INP(RxByteCnt[5]), .ZN(n18) );
  AO22X1 U89 ( .IN1(n109), .IN2(n17), .IN3(r_MinFL[4]), .IN4(n110), .Q(n108)
         );
  OR2X1 U90 ( .IN1(n109), .IN2(n17), .Q(n110) );
  INVX0 U91 ( .INP(RxByteCnt[4]), .ZN(n17) );
  AO22X1 U92 ( .IN1(n111), .IN2(n16), .IN3(r_MinFL[3]), .IN4(n112), .Q(n109)
         );
  OR2X1 U93 ( .IN1(n111), .IN2(n16), .Q(n112) );
  INVX0 U94 ( .INP(RxByteCnt[3]), .ZN(n16) );
  AO22X1 U95 ( .IN1(n113), .IN2(n15), .IN3(r_MinFL[2]), .IN4(n114), .Q(n111)
         );
  OR2X1 U96 ( .IN1(n113), .IN2(n15), .Q(n114) );
  INVX0 U97 ( .INP(RxByteCnt[2]), .ZN(n15) );
  AO22X1 U98 ( .IN1(r_MinFL[1]), .IN2(n23), .IN3(n115), .IN4(r_MinFL[0]), .Q(
        n113) );
  OA21X1 U99 ( .IN1(r_MinFL[1]), .IN2(n23), .IN3(n22), .Q(n115) );
  INVX0 U100 ( .INP(RxByteCnt[0]), .ZN(n22) );
  INVX0 U101 ( .INP(RxByteCnt[1]), .ZN(n23) );
  INVX0 U102 ( .INP(RxByteCnt[6]), .ZN(n68) );
  INVX0 U103 ( .INP(r_MinFL[6]), .ZN(n105) );
  INVX0 U104 ( .INP(r_MinFL[7]), .ZN(n103) );
  INVX0 U105 ( .INP(r_MinFL[8]), .ZN(n101) );
  INVX0 U106 ( .INP(r_MinFL[9]), .ZN(n99) );
  INVX0 U107 ( .INP(r_MinFL[10]), .ZN(n97) );
  INVX0 U108 ( .INP(r_MinFL[11]), .ZN(n95) );
  INVX0 U109 ( .INP(r_MinFL[12]), .ZN(n93) );
  INVX0 U110 ( .INP(r_MinFL[13]), .ZN(n91) );
  INVX0 U111 ( .INP(r_MinFL[14]), .ZN(n90) );
  NOR2X0 U112 ( .IN1(r_MinFL[14]), .IN2(n47), .QN(n88) );
  INVX0 U113 ( .INP(RxByteCnt[14]), .ZN(n47) );
  INVX0 U114 ( .INP(r_MinFL[15]), .ZN(n86) );
  AND3X1 U115 ( .IN1(MRxErr), .IN2(n116), .IN3(MRxDV), .Q(N7) );
  OR4X1 U116 ( .IN1(RxStateSFD), .IN2(RxStatePreamble), .IN3(n117), .IN4(n38), 
        .Q(n116) );
  OR2X1 U117 ( .IN1(RxStateData[1]), .IN2(RxStateData[0]), .Q(n38) );
  NOR2X0 U118 ( .IN1(Transmitting), .IN2(n118), .QN(n117) );
  INVX0 U119 ( .INP(RxStateIdle), .ZN(n118) );
endmodule


module eth_top ( wb_clk_i, wb_rst_i, wb_dat_i, wb_dat_o, wb_adr_i, wb_sel_i, 
        wb_we_i, wb_cyc_i, wb_stb_i, wb_ack_o, wb_err_o, m_wb_adr_o, 
        m_wb_sel_o, m_wb_we_o, m_wb_dat_o, m_wb_dat_i, m_wb_cyc_o, m_wb_stb_o, 
        m_wb_ack_i, m_wb_err_i, mtx_clk_pad_i, mtxd_pad_o, mtxen_pad_o, 
        mtxerr_pad_o, mrx_clk_pad_i, mrxd_pad_i, mrxdv_pad_i, mrxerr_pad_i, 
        mcoll_pad_i, mcrs_pad_i, mdc_pad_o, md_pad_i, md_pad_o, md_padoe_o, 
        int_o, data_source, test_mode, data_sourcea, test_si1, test_si2, 
        test_so2, test_si3, test_so3, test_si4, test_so4, test_si5, test_so5, 
        test_si6, test_so6, test_si7, test_so7, test_si8, test_se );
  input [31:0] wb_dat_i;
  output [31:0] wb_dat_o;
  input [11:2] wb_adr_i;
  input [3:0] wb_sel_i;
  output [31:0] m_wb_adr_o;
  output [3:0] m_wb_sel_o;
  output [31:0] m_wb_dat_o;
  input [31:0] m_wb_dat_i;
  output [3:0] mtxd_pad_o;
  input [3:0] mrxd_pad_i;
  input wb_clk_i, wb_rst_i, wb_we_i, wb_cyc_i, wb_stb_i, m_wb_ack_i,
         m_wb_err_i, mtx_clk_pad_i, mrx_clk_pad_i, mrxdv_pad_i, mrxerr_pad_i,
         mcoll_pad_i, mcrs_pad_i, md_pad_i, data_source, test_mode,
         data_sourcea, test_si1, test_si2, test_si3, test_si4, test_si5,
         test_si6, test_si7, test_si8, test_se;
  output wb_ack_o, wb_err_o, m_wb_we_o, m_wb_cyc_o, m_wb_stb_o, mtxen_pad_o,
         mtxerr_pad_o, mdc_pad_o, md_pad_o, md_padoe_o, int_o, test_so2,
         test_so3, test_so4, test_so5, test_so6, test_so7;
  wire   r_MiiNoPre, r_WCtrlData, r_RStat, r_ScanStat, Busy_stat, LinkFail,
         NValid_stat, WCtrlDataStart, RStatStart, UpdateMIIRX_DATAReg, BDAck,
         N9, N10, r_RecSmall, r_Pad, r_HugEn, r_CrcEn, r_DlyCrcEn, r_FullD,
         r_ExDfrEn, r_NoBckof, r_LoopBck, r_IFG, r_Pro, r_Bro, r_TxEn, r_RxEn,
         Busy_IRQ, RxE_IRQ, RxB_IRQ, TxE_IRQ, TxB_IRQ, r_TxFlow, r_RxFlow,
         r_PassAll, r_TxPauseRq, RstTxPauseRq, TxCtrlEndFrm, StartTxDone,
         SetPauseTimer, TPauseRq, TxStartFrm, TxEndFrm, TxUsedDataIn, TxDoneIn,
         TxAbortIn, RxValid, RxStartFrm, RxEndFrm, ReceiveEnd,
         ReceivedPacketGood, _0_net_, PadOut, _1_net_, CrcEnOut,
         ReceivedLengthOK, TxStartFrmOut, TxEndFrmOut, TxUsedData, TxDone,
         TxAbort, WillSendControlFrame, ReceivedPauseFrm, ControlFrmAddressOK,
         RxStatusWriteLatched_sync2, PerPacketCrcEn, PerPacketPad, MRxDV_Lb,
         MRxErr_Lb, TxCarrierSense, Collision, TxUnderRun, TxRetry,
         WillTransmit, ResetCollision, StartTxAbort, MaxCollisionOccured,
         LateCollision, DeferIndication, StatePreamble, Transmitting,
         RxByteCntEq0, RxByteCntGreat2, RxByteCntMaxFrame, RxCrcError,
         RxStateIdle, RxStatePreamble, RxStateSFD, RxAbort, AddressMiss,
         CarrierSense_Tx2, CarrierSense_Tx1, Collision_Tx1, WillTransmit_q,
         WillSendControlFrame_sync1, WillSendControlFrame_sync2,
         WillSendControlFrame_sync3, N23, N24, TxPauseRq_sync1,
         TxPauseRq_sync3, TxPauseRq_sync2, N25, RxAbort_latch, ShortFrame,
         LatchedMRxErr, InvalidSymbol, RxAbort_wb, RxAbort_sync1,
         RxAbortRst_sync1, LatchedCrcError, RxLateCollision, DribbleNibble,
         ReceivedPacketTooBig, LoadRxStatus, RetryLimit, LateCollLatched,
         DeferLatched, RstDeferLatched, CarrierSenseLost, n26, n27, n28, n29,
         n30, n33, n35, n36, n37, n89, n90, n91, n92, n94, n122, n123, n144,
         n145, n146, n147, n148, n150, n152, n154, n164, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242;
  wire   [7:0] r_ClkDiv;
  wire   [15:0] r_CtrlData;
  wire   [4:0] r_RGAD;
  wire   [4:0] r_FIAD;
  wire   [15:0] Prsd;
  wire   [3:0] BDCs;
  wire   [31:0] temp_wb_dat_o;
  wire   [31:0] RegDataOut;
  wire   [6:0] r_IPGT;
  wire   [6:0] r_IPGR1;
  wire   [6:0] r_IPGR2;
  wire   [15:0] r_MinFL;
  wire   [15:0] r_MaxFL;
  wire   [3:0] r_MaxRet;
  wire   [5:0] r_CollValid;
  wire   [47:0] r_MAC;
  wire   [7:0] r_TxBDNum;
  wire   [31:0] r_HASH0;
  wire   [31:0] r_HASH1;
  wire   [15:0] r_TxPauseTV;
  wire   [7:0] TxData;
  wire   [7:0] RxData;
  wire   [7:0] TxDataOut;
  wire   [3:0] MRxD_Lb;
  wire   [3:0] RetryCnt;
  wire   [1:0] StateData;
  wire   [15:0] RxByteCnt;
  wire   [1:0] RxStateData;
  wire   [3:0] RetryCntLatched;
  tri   [31:0] BD_WB_DAT_O;
  assign m_wb_adr_o[0] = 1'b0;
  assign m_wb_adr_o[1] = 1'b0;

  SDFFARX1 temp_wb_err_o_reg_reg ( .D(N10), .SI(wb_dat_o[31]), .SE(test_se), 
        .CLK(n164), .RSTB(n242), .Q(wb_err_o) );
  SDFFARX1 CarrierSense_Tx1_reg ( .D(mcrs_pad_i), .SI(test_si1), .SE(test_se), 
        .CLK(n154), .RSTB(n242), .Q(CarrierSense_Tx1) );
  SDFFARX1 CarrierSense_Tx2_reg ( .D(CarrierSense_Tx1), .SI(CarrierSense_Tx1), 
        .SE(test_se), .CLK(n154), .RSTB(n242), .Q(CarrierSense_Tx2), .QN(n27)
         );
  SDFFARX1 Collision_Tx1_reg ( .D(mcoll_pad_i), .SI(CarrierSense_Tx2), .SE(
        test_se), .CLK(n154), .RSTB(n242), .Q(Collision_Tx1) );
  SDFFARX1 RxAbortRst_reg ( .D(RxAbortRst_sync1), .SI(RstTxPauseRq), .SE(
        test_se), .CLK(n152), .RSTB(n242), .Q(n148), .QN(n33) );
  SDFFARX1 RxAbort_sync1_reg ( .D(RxAbort_latch), .SI(RxAbort_latch), .SE(
        test_se), .CLK(n164), .RSTB(n242), .Q(RxAbort_sync1) );
  SDFFARX1 RxAbort_wb_reg ( .D(RxAbort_sync1), .SI(RxAbort_sync1), .SE(test_se), .CLK(n164), .RSTB(n242), .Q(RxAbort_wb) );
  SDFFARX1 RxAbortRst_sync1_reg ( .D(RxAbort_wb), .SI(n148), .SE(test_se), 
        .CLK(n152), .RSTB(n242), .Q(RxAbortRst_sync1) );
  SDFFARX1 WillSendControlFrame_sync1_reg ( .D(WillSendControlFrame), .SI(
        TxPauseRq_sync3), .SE(test_se), .CLK(n164), .RSTB(n242), .Q(
        WillSendControlFrame_sync1) );
  SDFFARX1 WillSendControlFrame_sync2_reg ( .D(WillSendControlFrame_sync1), 
        .SI(WillSendControlFrame_sync1), .SE(test_se), .CLK(n164), .RSTB(n242), 
        .Q(WillSendControlFrame_sync2), .QN(n29) );
  SDFFARX1 WillSendControlFrame_sync3_reg ( .D(WillSendControlFrame_sync2), 
        .SI(WillSendControlFrame_sync2), .SE(test_se), .CLK(n164), .RSTB(n242), 
        .Q(WillSendControlFrame_sync3) );
  SDFFARX1 RstTxPauseRq_reg ( .D(N23), .SI(n123), .SE(test_se), .CLK(n164), 
        .RSTB(n242), .Q(RstTxPauseRq) );
  SDFFARX1 TxPauseRq_sync1_reg ( .D(N24), .SI(TPauseRq), .SE(test_se), .CLK(
        n154), .RSTB(n242), .Q(TxPauseRq_sync1) );
  SDFFARX1 TxPauseRq_sync2_reg ( .D(TxPauseRq_sync1), .SI(TxPauseRq_sync1), 
        .SE(test_se), .CLK(n154), .RSTB(n242), .Q(TxPauseRq_sync2), .QN(n28)
         );
  SDFFARX1 TxPauseRq_sync3_reg ( .D(TxPauseRq_sync2), .SI(TxPauseRq_sync2), 
        .SE(test_se), .CLK(n154), .RSTB(n242), .Q(TxPauseRq_sync3) );
  SDFFARX1 TPauseRq_reg ( .D(N25), .SI(n122), .SE(test_se), .CLK(n154), .RSTB(
        n242), .Q(TPauseRq) );
  SDFFX1 WillTransmit_q_reg ( .D(WillTransmit), .SI(n147), .SE(test_se), .CLK(
        n152), .Q(WillTransmit_q) );
  SDFFX1 WillTransmit_q2_reg ( .D(WillTransmit_q), .SI(
        WillSendControlFrame_sync3), .SE(test_se), .CLK(n152), .Q(n147), .QN(
        n26) );
  SDFFARX1 temp_wb_ack_o_reg_reg ( .D(N9), .SI(RxStateSFD), .SE(test_se), 
        .CLK(n164), .RSTB(n242), .Q(wb_ack_o), .QN(n30) );
  SDFFARX1 \temp_wb_dat_o_reg_reg[0]  ( .D(temp_wb_dat_o[0]), .SI(wb_ack_o), 
        .SE(test_se), .CLK(n164), .RSTB(n242), .Q(wb_dat_o[0]) );
  SDFFARX1 \temp_wb_dat_o_reg_reg[1]  ( .D(temp_wb_dat_o[1]), .SI(wb_dat_o[0]), 
        .SE(test_se), .CLK(n164), .RSTB(n242), .Q(wb_dat_o[1]) );
  SDFFARX1 \temp_wb_dat_o_reg_reg[2]  ( .D(temp_wb_dat_o[2]), .SI(wb_dat_o[1]), 
        .SE(test_se), .CLK(n164), .RSTB(n242), .Q(wb_dat_o[2]) );
  SDFFARX1 \temp_wb_dat_o_reg_reg[3]  ( .D(temp_wb_dat_o[3]), .SI(wb_dat_o[2]), 
        .SE(test_se), .CLK(n164), .RSTB(n242), .Q(wb_dat_o[3]) );
  SDFFARX1 \temp_wb_dat_o_reg_reg[4]  ( .D(temp_wb_dat_o[4]), .SI(wb_dat_o[3]), 
        .SE(test_se), .CLK(n164), .RSTB(n242), .Q(wb_dat_o[4]) );
  SDFFARX1 \temp_wb_dat_o_reg_reg[5]  ( .D(temp_wb_dat_o[5]), .SI(wb_dat_o[4]), 
        .SE(test_se), .CLK(n164), .RSTB(n242), .Q(wb_dat_o[5]) );
  SDFFARX1 \temp_wb_dat_o_reg_reg[6]  ( .D(temp_wb_dat_o[6]), .SI(wb_dat_o[5]), 
        .SE(test_se), .CLK(n164), .RSTB(n242), .Q(wb_dat_o[6]) );
  SDFFARX1 \temp_wb_dat_o_reg_reg[7]  ( .D(temp_wb_dat_o[7]), .SI(wb_dat_o[6]), 
        .SE(test_se), .CLK(n164), .RSTB(n242), .Q(wb_dat_o[7]) );
  SDFFARX1 \temp_wb_dat_o_reg_reg[8]  ( .D(temp_wb_dat_o[8]), .SI(wb_dat_o[7]), 
        .SE(test_se), .CLK(n164), .RSTB(n242), .Q(wb_dat_o[8]) );
  SDFFARX1 \temp_wb_dat_o_reg_reg[9]  ( .D(temp_wb_dat_o[9]), .SI(wb_dat_o[8]), 
        .SE(test_se), .CLK(n164), .RSTB(n242), .Q(wb_dat_o[9]) );
  SDFFARX1 \temp_wb_dat_o_reg_reg[10]  ( .D(temp_wb_dat_o[10]), .SI(
        wb_dat_o[9]), .SE(test_se), .CLK(n164), .RSTB(n242), .Q(wb_dat_o[10])
         );
  SDFFARX1 \temp_wb_dat_o_reg_reg[11]  ( .D(temp_wb_dat_o[11]), .SI(
        wb_dat_o[10]), .SE(test_se), .CLK(n164), .RSTB(n242), .Q(wb_dat_o[11])
         );
  SDFFARX1 \temp_wb_dat_o_reg_reg[12]  ( .D(temp_wb_dat_o[12]), .SI(
        wb_dat_o[11]), .SE(test_se), .CLK(n164), .RSTB(n242), .Q(wb_dat_o[12])
         );
  SDFFARX1 \temp_wb_dat_o_reg_reg[13]  ( .D(temp_wb_dat_o[13]), .SI(
        wb_dat_o[12]), .SE(test_se), .CLK(n164), .RSTB(n242), .Q(wb_dat_o[13])
         );
  SDFFARX1 \temp_wb_dat_o_reg_reg[14]  ( .D(temp_wb_dat_o[14]), .SI(
        wb_dat_o[13]), .SE(test_se), .CLK(n164), .RSTB(n242), .Q(wb_dat_o[14])
         );
  SDFFARX1 \temp_wb_dat_o_reg_reg[15]  ( .D(temp_wb_dat_o[15]), .SI(
        wb_dat_o[14]), .SE(test_se), .CLK(n164), .RSTB(n242), .Q(wb_dat_o[15])
         );
  SDFFARX1 \temp_wb_dat_o_reg_reg[16]  ( .D(temp_wb_dat_o[16]), .SI(
        wb_dat_o[15]), .SE(test_se), .CLK(n164), .RSTB(n242), .Q(wb_dat_o[16])
         );
  SDFFARX1 \temp_wb_dat_o_reg_reg[17]  ( .D(temp_wb_dat_o[17]), .SI(
        wb_dat_o[16]), .SE(test_se), .CLK(n164), .RSTB(n242), .Q(wb_dat_o[17])
         );
  SDFFARX1 \temp_wb_dat_o_reg_reg[18]  ( .D(temp_wb_dat_o[18]), .SI(
        wb_dat_o[17]), .SE(test_se), .CLK(n164), .RSTB(n242), .Q(wb_dat_o[18])
         );
  SDFFARX1 \temp_wb_dat_o_reg_reg[19]  ( .D(temp_wb_dat_o[19]), .SI(
        wb_dat_o[18]), .SE(test_se), .CLK(n164), .RSTB(n242), .Q(wb_dat_o[19])
         );
  SDFFARX1 \temp_wb_dat_o_reg_reg[20]  ( .D(temp_wb_dat_o[20]), .SI(
        wb_dat_o[19]), .SE(test_se), .CLK(n164), .RSTB(n242), .Q(wb_dat_o[20])
         );
  SDFFARX1 \temp_wb_dat_o_reg_reg[21]  ( .D(temp_wb_dat_o[21]), .SI(
        wb_dat_o[20]), .SE(test_se), .CLK(n164), .RSTB(n242), .Q(wb_dat_o[21])
         );
  SDFFARX1 \temp_wb_dat_o_reg_reg[22]  ( .D(temp_wb_dat_o[22]), .SI(
        wb_dat_o[21]), .SE(test_se), .CLK(n164), .RSTB(n242), .Q(wb_dat_o[22])
         );
  SDFFARX1 \temp_wb_dat_o_reg_reg[23]  ( .D(temp_wb_dat_o[23]), .SI(
        wb_dat_o[22]), .SE(test_se), .CLK(n164), .RSTB(n242), .Q(wb_dat_o[23])
         );
  SDFFARX1 \temp_wb_dat_o_reg_reg[24]  ( .D(temp_wb_dat_o[24]), .SI(
        wb_dat_o[23]), .SE(test_se), .CLK(n164), .RSTB(n242), .Q(wb_dat_o[24])
         );
  SDFFARX1 \temp_wb_dat_o_reg_reg[25]  ( .D(temp_wb_dat_o[25]), .SI(
        wb_dat_o[24]), .SE(test_se), .CLK(n164), .RSTB(n242), .Q(wb_dat_o[25])
         );
  SDFFARX1 \temp_wb_dat_o_reg_reg[26]  ( .D(temp_wb_dat_o[26]), .SI(
        wb_dat_o[25]), .SE(test_se), .CLK(n164), .RSTB(n242), .Q(wb_dat_o[26])
         );
  SDFFARX1 \temp_wb_dat_o_reg_reg[27]  ( .D(temp_wb_dat_o[27]), .SI(
        wb_dat_o[26]), .SE(test_se), .CLK(n164), .RSTB(n242), .Q(wb_dat_o[27])
         );
  SDFFARX1 \temp_wb_dat_o_reg_reg[28]  ( .D(temp_wb_dat_o[28]), .SI(
        wb_dat_o[27]), .SE(test_se), .CLK(n164), .RSTB(n242), .Q(wb_dat_o[28])
         );
  SDFFARX1 \temp_wb_dat_o_reg_reg[29]  ( .D(temp_wb_dat_o[29]), .SI(
        wb_dat_o[28]), .SE(test_se), .CLK(n164), .RSTB(n242), .Q(wb_dat_o[29])
         );
  SDFFARX1 \temp_wb_dat_o_reg_reg[30]  ( .D(temp_wb_dat_o[30]), .SI(
        wb_dat_o[29]), .SE(test_se), .CLK(n164), .RSTB(n242), .Q(wb_dat_o[30])
         );
  SDFFARX1 \temp_wb_dat_o_reg_reg[31]  ( .D(temp_wb_dat_o[31]), .SI(
        wb_dat_o[30]), .SE(test_se), .CLK(n164), .RSTB(n242), .Q(wb_dat_o[31])
         );
  SDFFARX1 RxAbort_latch_reg ( .D(n37), .SI(RxAbortRst_sync1), .SE(test_se), 
        .CLK(n152), .RSTB(n242), .Q(RxAbort_latch) );
  SDFFARX1 RxEnSync_reg ( .D(n36), .SI(RxAbort_wb), .SE(test_se), .CLK(n152), 
        .RSTB(n242), .Q(n122) );
  SDFFARX1 Collision_Tx2_reg ( .D(n35), .SI(Collision_Tx1), .SE(test_se), 
        .CLK(n154), .RSTB(n242), .Q(n123), .QN(n94) );
  eth_miim_test_1 miim1 ( .Clk(n164), .Reset(wb_rst_i), .Divider(r_ClkDiv), 
        .NoPre(r_MiiNoPre), .CtrlData(r_CtrlData), .Rgad(r_RGAD), .Fiad(r_FIAD), .WCtrlData(r_WCtrlData), .RStat(r_RStat), .ScanStat(r_ScanStat), .Mdi(
        md_pad_i), .Mdo(md_pad_o), .MdoEn(md_padoe_o), .Mdc(mdc_pad_o), .Busy(
        Busy_stat), .Prsd(Prsd), .LinkFail(LinkFail), .Nvalid(NValid_stat), 
        .WCtrlDataStart(WCtrlDataStart), .RStatStart(RStatStart), 
        .UpdateMIIRX_DATAReg(UpdateMIIRX_DATAReg), 
        .eth_top_test_point_11887_in(n218), .test_si(ShortFrame), .test_so(
        n145), .test_se(test_se) );
  eth_registers_test_1 ethreg1 ( .DataIn(wb_dat_i), .Address(wb_adr_i[9:2]), 
        .Rw(wb_we_i), .Cs({n92, n91, n90, n89}), .Clk(n164), .Reset(wb_rst_i), 
        .DataOut(RegDataOut), .r_RecSmall(r_RecSmall), .r_Pad(r_Pad), 
        .r_HugEn(r_HugEn), .r_CrcEn(r_CrcEn), .r_DlyCrcEn(r_DlyCrcEn), 
        .r_FullD(r_FullD), .r_ExDfrEn(r_ExDfrEn), .r_NoBckof(r_NoBckof), 
        .r_LoopBck(r_LoopBck), .r_IFG(r_IFG), .r_Pro(r_Pro), .r_Bro(r_Bro), 
        .r_TxEn(r_TxEn), .r_RxEn(r_RxEn), .TxB_IRQ(TxB_IRQ), .TxE_IRQ(TxE_IRQ), 
        .RxB_IRQ(RxB_IRQ), .RxE_IRQ(RxE_IRQ), .Busy_IRQ(Busy_IRQ), .r_IPGT(
        r_IPGT), .r_IPGR1(r_IPGR1), .r_IPGR2(r_IPGR2), .r_MinFL(r_MinFL), 
        .r_MaxFL(r_MaxFL), .r_MaxRet(r_MaxRet), .r_CollValid(r_CollValid), 
        .r_TxFlow(r_TxFlow), .r_RxFlow(r_RxFlow), .r_PassAll(r_PassAll), 
        .r_MiiNoPre(r_MiiNoPre), .r_ClkDiv(r_ClkDiv), .r_WCtrlData(r_WCtrlData), .r_RStat(r_RStat), .r_ScanStat(r_ScanStat), .r_RGAD(r_RGAD), .r_FIAD(r_FIAD), 
        .r_CtrlData(r_CtrlData), .NValid_stat(NValid_stat), .Busy_stat(
        Busy_stat), .LinkFail(LinkFail), .r_MAC(r_MAC), .WCtrlDataStart(
        WCtrlDataStart), .RStatStart(RStatStart), .UpdateMIIRX_DATAReg(
        UpdateMIIRX_DATAReg), .Prsd(Prsd), .r_TxBDNum(r_TxBDNum), .int_o(int_o), .r_HASH0(r_HASH0), .r_HASH1(r_HASH1), .r_TxPauseTV(r_TxPauseTV), 
        .r_TxPauseRq(r_TxPauseRq), .RstTxPauseRq(RstTxPauseRq), .TxCtrlEndFrm(
        TxCtrlEndFrm), .StartTxDone(StartTxDone), .TxClk(n154), .RxClk(n152), 
        .SetPauseTimer(SetPauseTimer), .eth_top_test_point_11887_in(n217), 
        .test_si(WillTransmit_q), .test_so(n146), .test_se(test_se) );
  eth_maccontrol_test_1 maccontrol1 ( .MTxClk(n154), .MRxClk(n152), .TxReset(
        wb_rst_i), .RxReset(wb_rst_i), .TPauseRq(TPauseRq), .TxDataIn(TxData), 
        .TxStartFrmIn(TxStartFrm), .TxUsedDataIn(TxUsedDataIn), .TxEndFrmIn(
        TxEndFrm), .TxDoneIn(TxDoneIn), .TxAbortIn(TxAbortIn), .RxData(RxData), 
        .RxValid(RxValid), .RxStartFrm(RxStartFrm), .RxEndFrm(RxEndFrm), 
        .ReceiveEnd(ReceiveEnd), .ReceivedPacketGood(ReceivedPacketGood), 
        .ReceivedLengthOK(ReceivedLengthOK), .TxFlow(r_TxFlow), .RxFlow(
        r_RxFlow), .DlyCrcEn(r_DlyCrcEn), .TxPauseTV(r_TxPauseTV), .MAC(r_MAC), 
        .PadIn(_0_net_), .PadOut(PadOut), .CrcEnIn(_1_net_), .CrcEnOut(
        CrcEnOut), .TxDataOut(TxDataOut), .TxStartFrmOut(TxStartFrmOut), 
        .TxEndFrmOut(TxEndFrmOut), .TxDoneOut(TxDone), .TxAbortOut(TxAbort), 
        .TxUsedDataOut(TxUsedData), .WillSendControlFrame(WillSendControlFrame), .TxCtrlEndFrm(TxCtrlEndFrm), .ReceivedPauseFrm(ReceivedPauseFrm), 
        .ControlFrmAddressOK(ControlFrmAddressOK), .SetPauseTimer(
        SetPauseTimer), .r_PassAll(r_PassAll), .RxStatusWriteLatched_sync2(
        RxStatusWriteLatched_sync2), .eth_top_data_sourcea_in(data_sourcea), 
        .eth_top_test_mode_in(test_mode), .eth_top_test_point_11887_in(n218), 
        .test_si(n146), .test_se(test_se) );
  eth_txethmac_test_1 txethmac1 ( .MTxClk(n154), .Reset(wb_rst_i), 
        .TxStartFrm(TxStartFrmOut), .TxEndFrm(TxEndFrmOut), .TxUnderRun(
        TxUnderRun), .TxData(TxDataOut), .CarrierSense(TxCarrierSense), 
        .Collision(Collision), .Pad(PadOut), .CrcEn(CrcEnOut), .FullD(r_FullD), 
        .HugEn(r_HugEn), .DlyCrcEn(r_DlyCrcEn), .MinFL(r_MinFL), .MaxFL(
        r_MaxFL), .IPGT(r_IPGT), .IPGR1(r_IPGR1), .IPGR2(r_IPGR2), .CollValid(
        r_CollValid), .MaxRet(r_MaxRet), .NoBckof(r_NoBckof), .ExDfrEn(
        r_ExDfrEn), .MTxD(mtxd_pad_o), .MTxEn(mtxen_pad_o), .MTxErr(
        mtxerr_pad_o), .TxDone(TxDoneIn), .TxRetry(TxRetry), .TxAbort(
        TxAbortIn), .TxUsedData(TxUsedDataIn), .WillTransmit(WillTransmit), 
        .ResetCollision(ResetCollision), .RetryCnt(RetryCnt), .StartTxDone(
        StartTxDone), .StartTxAbort(StartTxAbort), .MaxCollisionOccured(
        MaxCollisionOccured), .LateCollision(LateCollision), .DeferIndication(
        DeferIndication), .StatePreamble(StatePreamble), .StateData(StateData), 
        .eth_top_test_point_11887_in(n150), .test_si2(n144), .test_si1(
        wb_err_o), .test_se(test_se) );
  eth_rxethmac_test_1 rxethmac1 ( .MRxClk(n152), .MRxDV(MRxDV_Lb), .MRxD(
        MRxD_Lb), .Reset(wb_rst_i), .Transmitting(Transmitting), .MaxFL(
        r_MaxFL), .r_IFG(r_IFG), .HugEn(r_HugEn), .DlyCrcEn(r_DlyCrcEn), 
        .RxData(RxData), .RxValid(RxValid), .RxStartFrm(RxStartFrm), 
        .RxEndFrm(RxEndFrm), .ByteCnt(RxByteCnt), .ByteCntEq0(RxByteCntEq0), 
        .ByteCntGreat2(RxByteCntGreat2), .ByteCntMaxFrame(RxByteCntMaxFrame), 
        .CrcError(RxCrcError), .StateIdle(RxStateIdle), .StatePreamble(
        RxStatePreamble), .StateSFD(RxStateSFD), .StateData(RxStateData), 
        .MAC(r_MAC), .r_Pro(r_Pro), .r_Bro(r_Bro), .r_HASH0(r_HASH0), 
        .r_HASH1(r_HASH1), .RxAbort(RxAbort), .AddressMiss(AddressMiss), 
        .PassAll(r_PassAll), .ControlFrmAddressOK(ControlFrmAddressOK), 
        .eth_top_test_point_11887_in(n218), .test_si(n145), .test_se(test_se)
         );
  eth_wishbone_test_1 wishbone ( .WB_CLK_I(n164), .WB_DAT_I(wb_dat_i), 
        .WB_DAT_O(BD_WB_DAT_O), .WB_ADR_I(wb_adr_i[9:2]), .WB_WE_I(wb_we_i), 
        .WB_ACK_O(BDAck), .BDCs(BDCs), .Reset(wb_rst_i), .m_wb_adr_o(
        m_wb_adr_o[31:2]), .m_wb_sel_o(m_wb_sel_o), .m_wb_we_o(m_wb_we_o), 
        .m_wb_dat_o(m_wb_dat_o), .m_wb_dat_i(m_wb_dat_i), .m_wb_cyc_o(
        m_wb_cyc_o), .m_wb_stb_o(m_wb_stb_o), .m_wb_ack_i(m_wb_ack_i), 
        .m_wb_err_i(m_wb_err_i), .MTxClk(n154), .TxStartFrm(TxStartFrm), 
        .TxEndFrm(TxEndFrm), .TxUsedData(TxUsedData), .TxData(TxData), 
        .TxRetry(TxRetry), .TxAbort(TxAbort), .TxUnderRun(TxUnderRun), 
        .TxDone(TxDone), .PerPacketCrcEn(PerPacketCrcEn), .PerPacketPad(
        PerPacketPad), .MRxClk(n152), .RxData(RxData), .RxValid(RxValid), 
        .RxStartFrm(RxStartFrm), .RxEndFrm(RxEndFrm), .RxAbort(RxAbort_wb), 
        .RxStatusWriteLatched_sync2(RxStatusWriteLatched_sync2), .r_TxEn(
        r_TxEn), .r_RxEn(r_RxEn), .r_TxBDNum(r_TxBDNum), .r_RxFlow(r_RxFlow), 
        .r_PassAll(r_PassAll), .TxB_IRQ(TxB_IRQ), .TxE_IRQ(TxE_IRQ), .RxB_IRQ(
        RxB_IRQ), .RxE_IRQ(RxE_IRQ), .Busy_IRQ(Busy_IRQ), .InvalidSymbol(
        InvalidSymbol), .LatchedCrcError(LatchedCrcError), .RxLateCollision(
        RxLateCollision), .ShortFrame(ShortFrame), .DribbleNibble(
        DribbleNibble), .ReceivedPacketTooBig(ReceivedPacketTooBig), 
        .RxLength(RxByteCnt), .LoadRxStatus(LoadRxStatus), 
        .ReceivedPacketGood(ReceivedPacketGood), .AddressMiss(AddressMiss), 
        .ReceivedPauseFrm(ReceivedPauseFrm), .RetryCntLatched(RetryCntLatched), 
        .RetryLimit(RetryLimit), .LateCollLatched(LateCollLatched), 
        .DeferLatched(DeferLatched), .RstDeferLatched(RstDeferLatched), 
        .CarrierSenseLost(CarrierSenseLost), .eth_top_test_point_11887_in(n150), .test_si8(test_si8), .test_si7(test_si7), .test_si6(test_si6), .test_si5(
        test_si5), .test_si4(test_si4), .test_si3(test_si3), .test_si2(
        test_si2), .test_si1(StatePreamble), .test_so7(test_so7), .test_so6(
        test_so6), .test_so5(test_so5), .test_so4(test_so4), .test_so3(
        test_so3), .test_so2(test_so2), .test_so1(n144), .test_se(test_se) );
  eth_macstatus_test_1 macstatus1 ( .MRxClk(n152), .Reset(wb_rst_i), 
        .ReceivedLengthOK(ReceivedLengthOK), .ReceiveEnd(ReceiveEnd), 
        .ReceivedPacketGood(ReceivedPacketGood), .RxCrcError(RxCrcError), 
        .MRxErr(MRxErr_Lb), .MRxDV(MRxDV_Lb), .RxStateSFD(RxStateSFD), 
        .RxStateData(RxStateData), .RxStatePreamble(RxStatePreamble), 
        .RxStateIdle(RxStateIdle), .Transmitting(Transmitting), .RxByteCnt(
        RxByteCnt), .RxByteCntEq0(RxByteCntEq0), .RxByteCntGreat2(
        RxByteCntGreat2), .RxByteCntMaxFrame(RxByteCntMaxFrame), 
        .InvalidSymbol(InvalidSymbol), .MRxD(MRxD_Lb), .LatchedCrcError(
        LatchedCrcError), .Collision(mcoll_pad_i), .CollValid(r_CollValid), 
        .RxLateCollision(RxLateCollision), .r_RecSmall(r_RecSmall), .r_MinFL(
        r_MinFL), .r_MaxFL(r_MaxFL), .ShortFrame(ShortFrame), .DribbleNibble(
        DribbleNibble), .ReceivedPacketTooBig(ReceivedPacketTooBig), .r_HugEn(
        r_HugEn), .LoadRxStatus(LoadRxStatus), .StartTxDone(StartTxDone), 
        .StartTxAbort(StartTxAbort), .RetryCnt(RetryCnt), .RetryCntLatched(
        RetryCntLatched), .MTxClk(n154), .MaxCollisionOccured(
        MaxCollisionOccured), .RetryLimit(RetryLimit), .LateCollision(
        LateCollision), .LateCollLatched(LateCollLatched), .DeferIndication(
        DeferIndication), .DeferLatched(DeferLatched), .RstDeferLatched(
        RstDeferLatched), .TxStartFrm(TxStartFrmOut), .StatePreamble(
        StatePreamble), .StateData(StateData), .CarrierSense(CarrierSense_Tx2), 
        .CarrierSenseLost(CarrierSenseLost), .TxUsedData(TxUsedDataIn), 
        .LatchedMRxErr(LatchedMRxErr), .Loopback(r_LoopBck), .r_FullD(r_FullD), 
        .eth_top_test_point_11887_in(n218), .test_si(WillSendControlFrame), 
        .test_se(test_se) );
  MUX21X1 U230 ( .IN1(wb_rst_i), .IN2(data_sourcea), .S(test_mode), .Q(n150)
         );
  INVX0 U231 ( .INP(n150), .ZN(n216) );
  INVX0 U232 ( .INP(n216), .ZN(n217) );
  INVX0 U233 ( .INP(n216), .ZN(n218) );
  NOR2X1 U234 ( .IN1(wb_we_i), .IN2(n220), .QN(n219) );
  INVX1 U235 ( .INP(n150), .ZN(n242) );
  MUX21X1 U236 ( .IN1(BD_WB_DAT_O[9]), .IN2(RegDataOut[9]), .S(n219), .Q(
        temp_wb_dat_o[9]) );
  MUX21X1 U237 ( .IN1(BD_WB_DAT_O[8]), .IN2(RegDataOut[8]), .S(n219), .Q(
        temp_wb_dat_o[8]) );
  MUX21X1 U238 ( .IN1(BD_WB_DAT_O[7]), .IN2(RegDataOut[7]), .S(n219), .Q(
        temp_wb_dat_o[7]) );
  MUX21X1 U239 ( .IN1(BD_WB_DAT_O[6]), .IN2(RegDataOut[6]), .S(n219), .Q(
        temp_wb_dat_o[6]) );
  MUX21X1 U240 ( .IN1(BD_WB_DAT_O[5]), .IN2(RegDataOut[5]), .S(n219), .Q(
        temp_wb_dat_o[5]) );
  MUX21X1 U241 ( .IN1(BD_WB_DAT_O[4]), .IN2(RegDataOut[4]), .S(n219), .Q(
        temp_wb_dat_o[4]) );
  MUX21X1 U242 ( .IN1(BD_WB_DAT_O[3]), .IN2(RegDataOut[3]), .S(n219), .Q(
        temp_wb_dat_o[3]) );
  MUX21X1 U243 ( .IN1(BD_WB_DAT_O[31]), .IN2(RegDataOut[31]), .S(n219), .Q(
        temp_wb_dat_o[31]) );
  MUX21X1 U244 ( .IN1(BD_WB_DAT_O[30]), .IN2(RegDataOut[30]), .S(n219), .Q(
        temp_wb_dat_o[30]) );
  MUX21X1 U245 ( .IN1(BD_WB_DAT_O[2]), .IN2(RegDataOut[2]), .S(n219), .Q(
        temp_wb_dat_o[2]) );
  MUX21X1 U246 ( .IN1(BD_WB_DAT_O[29]), .IN2(RegDataOut[29]), .S(n219), .Q(
        temp_wb_dat_o[29]) );
  MUX21X1 U247 ( .IN1(BD_WB_DAT_O[28]), .IN2(RegDataOut[28]), .S(n219), .Q(
        temp_wb_dat_o[28]) );
  MUX21X1 U248 ( .IN1(BD_WB_DAT_O[27]), .IN2(RegDataOut[27]), .S(n219), .Q(
        temp_wb_dat_o[27]) );
  MUX21X1 U249 ( .IN1(BD_WB_DAT_O[26]), .IN2(RegDataOut[26]), .S(n219), .Q(
        temp_wb_dat_o[26]) );
  MUX21X1 U250 ( .IN1(BD_WB_DAT_O[25]), .IN2(RegDataOut[25]), .S(n219), .Q(
        temp_wb_dat_o[25]) );
  MUX21X1 U251 ( .IN1(BD_WB_DAT_O[24]), .IN2(RegDataOut[24]), .S(n219), .Q(
        temp_wb_dat_o[24]) );
  MUX21X1 U252 ( .IN1(BD_WB_DAT_O[23]), .IN2(RegDataOut[23]), .S(n219), .Q(
        temp_wb_dat_o[23]) );
  MUX21X1 U253 ( .IN1(BD_WB_DAT_O[22]), .IN2(RegDataOut[22]), .S(n219), .Q(
        temp_wb_dat_o[22]) );
  MUX21X1 U254 ( .IN1(BD_WB_DAT_O[21]), .IN2(RegDataOut[21]), .S(n219), .Q(
        temp_wb_dat_o[21]) );
  MUX21X1 U255 ( .IN1(BD_WB_DAT_O[20]), .IN2(RegDataOut[20]), .S(n219), .Q(
        temp_wb_dat_o[20]) );
  MUX21X1 U256 ( .IN1(BD_WB_DAT_O[1]), .IN2(RegDataOut[1]), .S(n219), .Q(
        temp_wb_dat_o[1]) );
  MUX21X1 U257 ( .IN1(BD_WB_DAT_O[19]), .IN2(RegDataOut[19]), .S(n219), .Q(
        temp_wb_dat_o[19]) );
  MUX21X1 U258 ( .IN1(BD_WB_DAT_O[18]), .IN2(RegDataOut[18]), .S(n219), .Q(
        temp_wb_dat_o[18]) );
  MUX21X1 U259 ( .IN1(BD_WB_DAT_O[17]), .IN2(RegDataOut[17]), .S(n219), .Q(
        temp_wb_dat_o[17]) );
  MUX21X1 U260 ( .IN1(BD_WB_DAT_O[16]), .IN2(RegDataOut[16]), .S(n219), .Q(
        temp_wb_dat_o[16]) );
  MUX21X1 U261 ( .IN1(BD_WB_DAT_O[15]), .IN2(RegDataOut[15]), .S(n219), .Q(
        temp_wb_dat_o[15]) );
  MUX21X1 U262 ( .IN1(BD_WB_DAT_O[14]), .IN2(RegDataOut[14]), .S(n219), .Q(
        temp_wb_dat_o[14]) );
  MUX21X1 U263 ( .IN1(BD_WB_DAT_O[13]), .IN2(RegDataOut[13]), .S(n219), .Q(
        temp_wb_dat_o[13]) );
  MUX21X1 U264 ( .IN1(BD_WB_DAT_O[12]), .IN2(RegDataOut[12]), .S(n219), .Q(
        temp_wb_dat_o[12]) );
  MUX21X1 U265 ( .IN1(BD_WB_DAT_O[11]), .IN2(RegDataOut[11]), .S(n219), .Q(
        temp_wb_dat_o[11]) );
  MUX21X1 U266 ( .IN1(BD_WB_DAT_O[10]), .IN2(RegDataOut[10]), .S(n219), .Q(
        temp_wb_dat_o[10]) );
  MUX21X1 U267 ( .IN1(BD_WB_DAT_O[0]), .IN2(RegDataOut[0]), .S(n219), .Q(
        temp_wb_dat_o[0]) );
  NOR2X0 U268 ( .IN1(n220), .IN2(n221), .QN(n92) );
  NOR2X0 U269 ( .IN1(n220), .IN2(n222), .QN(n91) );
  NOR2X0 U270 ( .IN1(n220), .IN2(n223), .QN(n90) );
  NOR2X0 U271 ( .IN1(n220), .IN2(n224), .QN(n89) );
  INVX0 U272 ( .INP(n225), .ZN(n220) );
  AO221X1 U273 ( .IN1(ShortFrame), .IN2(n226), .IN3(n33), .IN4(RxAbort_latch), 
        .IN5(n227), .Q(n37) );
  AO221X1 U274 ( .IN1(LatchedMRxErr), .IN2(n228), .IN3(ReceivedPauseFrm), 
        .IN4(n229), .IN5(RxAbort), .Q(n227) );
  INVX0 U275 ( .INP(r_PassAll), .ZN(n229) );
  INVX0 U276 ( .INP(InvalidSymbol), .ZN(n228) );
  INVX0 U277 ( .INP(r_RecSmall), .ZN(n226) );
  MUX21X1 U278 ( .IN1(r_RxEn), .IN2(n122), .S(mrxdv_pad_i), .Q(n36) );
  NOR2X0 U279 ( .IN1(ResetCollision), .IN2(n230), .QN(n35) );
  NOR2X0 U280 ( .IN1(n123), .IN2(Collision_Tx1), .QN(n230) );
  AO21X1 U281 ( .IN1(wb_clk_i), .IN2(n231), .IN3(n232), .Q(n164) );
  AO21X1 U282 ( .IN1(mtx_clk_pad_i), .IN2(n231), .IN3(n232), .Q(n154) );
  AO21X1 U283 ( .IN1(mrx_clk_pad_i), .IN2(n231), .IN3(n232), .Q(n152) );
  AND2X1 U284 ( .IN1(data_source), .IN2(test_mode), .Q(n232) );
  INVX0 U285 ( .INP(test_mode), .ZN(n231) );
  OR2X1 U286 ( .IN1(PerPacketCrcEn), .IN2(r_CrcEn), .Q(_1_net_) );
  OR2X1 U287 ( .IN1(PerPacketPad), .IN2(r_Pad), .Q(_0_net_) );
  NOR2X0 U288 ( .IN1(r_FullD), .IN2(n27), .QN(TxCarrierSense) );
  NOR2X0 U289 ( .IN1(r_FullD), .IN2(n26), .QN(Transmitting) );
  OA21X1 U290 ( .IN1(n225), .IN2(BDAck), .IN3(n30), .Q(N9) );
  NOR2X0 U291 ( .IN1(n233), .IN2(wb_adr_i[10]), .QN(n225) );
  NOR2X0 U292 ( .IN1(n28), .IN2(TxPauseRq_sync3), .QN(N25) );
  AND2X1 U293 ( .IN1(r_TxPauseRq), .IN2(r_TxFlow), .Q(N24) );
  NOR2X0 U294 ( .IN1(n29), .IN2(WillSendControlFrame_sync3), .QN(N23) );
  NOR4X0 U295 ( .IN1(wb_err_o), .IN2(n234), .IN3(n235), .IN4(n236), .QN(N10)
         );
  INVX0 U296 ( .INP(wb_stb_i), .ZN(n236) );
  INVX0 U297 ( .INP(wb_cyc_i), .ZN(n235) );
  MUX21X1 U298 ( .IN1(n237), .IN2(mtxerr_pad_o), .S(r_LoopBck), .Q(MRxErr_Lb)
         );
  AND2X1 U299 ( .IN1(mrxerr_pad_i), .IN2(n122), .Q(n237) );
  MUX21X1 U300 ( .IN1(mrxd_pad_i[3]), .IN2(mtxd_pad_o[3]), .S(r_LoopBck), .Q(
        MRxD_Lb[3]) );
  MUX21X1 U301 ( .IN1(mrxd_pad_i[2]), .IN2(mtxd_pad_o[2]), .S(r_LoopBck), .Q(
        MRxD_Lb[2]) );
  MUX21X1 U302 ( .IN1(mrxd_pad_i[1]), .IN2(mtxd_pad_o[1]), .S(r_LoopBck), .Q(
        MRxD_Lb[1]) );
  MUX21X1 U303 ( .IN1(mrxd_pad_i[0]), .IN2(mtxd_pad_o[0]), .S(r_LoopBck), .Q(
        MRxD_Lb[0]) );
  MUX21X1 U304 ( .IN1(n238), .IN2(mtxen_pad_o), .S(r_LoopBck), .Q(MRxDV_Lb) );
  AND2X1 U305 ( .IN1(n122), .IN2(mrxdv_pad_i), .Q(n238) );
  NOR2X0 U306 ( .IN1(r_FullD), .IN2(n94), .QN(Collision) );
  NOR2X0 U307 ( .IN1(n221), .IN2(n239), .QN(BDCs[3]) );
  INVX0 U308 ( .INP(wb_sel_i[3]), .ZN(n221) );
  NOR2X0 U309 ( .IN1(n222), .IN2(n239), .QN(BDCs[2]) );
  INVX0 U310 ( .INP(wb_sel_i[2]), .ZN(n222) );
  NOR2X0 U311 ( .IN1(n223), .IN2(n239), .QN(BDCs[1]) );
  INVX0 U312 ( .INP(wb_sel_i[1]), .ZN(n223) );
  NOR2X0 U313 ( .IN1(n224), .IN2(n239), .QN(BDCs[0]) );
  NAND2X0 U314 ( .IN1(wb_adr_i[10]), .IN2(n240), .QN(n239) );
  INVX0 U315 ( .INP(n233), .ZN(n240) );
  NAND3X0 U316 ( .IN1(wb_cyc_i), .IN2(n234), .IN3(wb_stb_i), .QN(n233) );
  NOR2X0 U317 ( .IN1(n241), .IN2(wb_adr_i[11]), .QN(n234) );
  NOR4X0 U318 ( .IN1(wb_sel_i[3]), .IN2(wb_sel_i[2]), .IN3(wb_sel_i[1]), .IN4(
        wb_sel_i[0]), .QN(n241) );
  INVX0 U319 ( .INP(wb_sel_i[0]), .ZN(n224) );
endmodule

